module Hash(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [7:0]   io_pipe_phv_in_data_160,
  input  [7:0]   io_pipe_phv_in_data_161,
  input  [7:0]   io_pipe_phv_in_data_162,
  input  [7:0]   io_pipe_phv_in_data_163,
  input  [7:0]   io_pipe_phv_in_data_164,
  input  [7:0]   io_pipe_phv_in_data_165,
  input  [7:0]   io_pipe_phv_in_data_166,
  input  [7:0]   io_pipe_phv_in_data_167,
  input  [7:0]   io_pipe_phv_in_data_168,
  input  [7:0]   io_pipe_phv_in_data_169,
  input  [7:0]   io_pipe_phv_in_data_170,
  input  [7:0]   io_pipe_phv_in_data_171,
  input  [7:0]   io_pipe_phv_in_data_172,
  input  [7:0]   io_pipe_phv_in_data_173,
  input  [7:0]   io_pipe_phv_in_data_174,
  input  [7:0]   io_pipe_phv_in_data_175,
  input  [7:0]   io_pipe_phv_in_data_176,
  input  [7:0]   io_pipe_phv_in_data_177,
  input  [7:0]   io_pipe_phv_in_data_178,
  input  [7:0]   io_pipe_phv_in_data_179,
  input  [7:0]   io_pipe_phv_in_data_180,
  input  [7:0]   io_pipe_phv_in_data_181,
  input  [7:0]   io_pipe_phv_in_data_182,
  input  [7:0]   io_pipe_phv_in_data_183,
  input  [7:0]   io_pipe_phv_in_data_184,
  input  [7:0]   io_pipe_phv_in_data_185,
  input  [7:0]   io_pipe_phv_in_data_186,
  input  [7:0]   io_pipe_phv_in_data_187,
  input  [7:0]   io_pipe_phv_in_data_188,
  input  [7:0]   io_pipe_phv_in_data_189,
  input  [7:0]   io_pipe_phv_in_data_190,
  input  [7:0]   io_pipe_phv_in_data_191,
  input  [7:0]   io_pipe_phv_in_data_192,
  input  [7:0]   io_pipe_phv_in_data_193,
  input  [7:0]   io_pipe_phv_in_data_194,
  input  [7:0]   io_pipe_phv_in_data_195,
  input  [7:0]   io_pipe_phv_in_data_196,
  input  [7:0]   io_pipe_phv_in_data_197,
  input  [7:0]   io_pipe_phv_in_data_198,
  input  [7:0]   io_pipe_phv_in_data_199,
  input  [7:0]   io_pipe_phv_in_data_200,
  input  [7:0]   io_pipe_phv_in_data_201,
  input  [7:0]   io_pipe_phv_in_data_202,
  input  [7:0]   io_pipe_phv_in_data_203,
  input  [7:0]   io_pipe_phv_in_data_204,
  input  [7:0]   io_pipe_phv_in_data_205,
  input  [7:0]   io_pipe_phv_in_data_206,
  input  [7:0]   io_pipe_phv_in_data_207,
  input  [7:0]   io_pipe_phv_in_data_208,
  input  [7:0]   io_pipe_phv_in_data_209,
  input  [7:0]   io_pipe_phv_in_data_210,
  input  [7:0]   io_pipe_phv_in_data_211,
  input  [7:0]   io_pipe_phv_in_data_212,
  input  [7:0]   io_pipe_phv_in_data_213,
  input  [7:0]   io_pipe_phv_in_data_214,
  input  [7:0]   io_pipe_phv_in_data_215,
  input  [7:0]   io_pipe_phv_in_data_216,
  input  [7:0]   io_pipe_phv_in_data_217,
  input  [7:0]   io_pipe_phv_in_data_218,
  input  [7:0]   io_pipe_phv_in_data_219,
  input  [7:0]   io_pipe_phv_in_data_220,
  input  [7:0]   io_pipe_phv_in_data_221,
  input  [7:0]   io_pipe_phv_in_data_222,
  input  [7:0]   io_pipe_phv_in_data_223,
  input  [7:0]   io_pipe_phv_in_data_224,
  input  [7:0]   io_pipe_phv_in_data_225,
  input  [7:0]   io_pipe_phv_in_data_226,
  input  [7:0]   io_pipe_phv_in_data_227,
  input  [7:0]   io_pipe_phv_in_data_228,
  input  [7:0]   io_pipe_phv_in_data_229,
  input  [7:0]   io_pipe_phv_in_data_230,
  input  [7:0]   io_pipe_phv_in_data_231,
  input  [7:0]   io_pipe_phv_in_data_232,
  input  [7:0]   io_pipe_phv_in_data_233,
  input  [7:0]   io_pipe_phv_in_data_234,
  input  [7:0]   io_pipe_phv_in_data_235,
  input  [7:0]   io_pipe_phv_in_data_236,
  input  [7:0]   io_pipe_phv_in_data_237,
  input  [7:0]   io_pipe_phv_in_data_238,
  input  [7:0]   io_pipe_phv_in_data_239,
  input  [7:0]   io_pipe_phv_in_data_240,
  input  [7:0]   io_pipe_phv_in_data_241,
  input  [7:0]   io_pipe_phv_in_data_242,
  input  [7:0]   io_pipe_phv_in_data_243,
  input  [7:0]   io_pipe_phv_in_data_244,
  input  [7:0]   io_pipe_phv_in_data_245,
  input  [7:0]   io_pipe_phv_in_data_246,
  input  [7:0]   io_pipe_phv_in_data_247,
  input  [7:0]   io_pipe_phv_in_data_248,
  input  [7:0]   io_pipe_phv_in_data_249,
  input  [7:0]   io_pipe_phv_in_data_250,
  input  [7:0]   io_pipe_phv_in_data_251,
  input  [7:0]   io_pipe_phv_in_data_252,
  input  [7:0]   io_pipe_phv_in_data_253,
  input  [7:0]   io_pipe_phv_in_data_254,
  input  [7:0]   io_pipe_phv_in_data_255,
  input  [7:0]   io_pipe_phv_in_data_256,
  input  [7:0]   io_pipe_phv_in_data_257,
  input  [7:0]   io_pipe_phv_in_data_258,
  input  [7:0]   io_pipe_phv_in_data_259,
  input  [7:0]   io_pipe_phv_in_data_260,
  input  [7:0]   io_pipe_phv_in_data_261,
  input  [7:0]   io_pipe_phv_in_data_262,
  input  [7:0]   io_pipe_phv_in_data_263,
  input  [7:0]   io_pipe_phv_in_data_264,
  input  [7:0]   io_pipe_phv_in_data_265,
  input  [7:0]   io_pipe_phv_in_data_266,
  input  [7:0]   io_pipe_phv_in_data_267,
  input  [7:0]   io_pipe_phv_in_data_268,
  input  [7:0]   io_pipe_phv_in_data_269,
  input  [7:0]   io_pipe_phv_in_data_270,
  input  [7:0]   io_pipe_phv_in_data_271,
  input  [7:0]   io_pipe_phv_in_data_272,
  input  [7:0]   io_pipe_phv_in_data_273,
  input  [7:0]   io_pipe_phv_in_data_274,
  input  [7:0]   io_pipe_phv_in_data_275,
  input  [7:0]   io_pipe_phv_in_data_276,
  input  [7:0]   io_pipe_phv_in_data_277,
  input  [7:0]   io_pipe_phv_in_data_278,
  input  [7:0]   io_pipe_phv_in_data_279,
  input  [7:0]   io_pipe_phv_in_data_280,
  input  [7:0]   io_pipe_phv_in_data_281,
  input  [7:0]   io_pipe_phv_in_data_282,
  input  [7:0]   io_pipe_phv_in_data_283,
  input  [7:0]   io_pipe_phv_in_data_284,
  input  [7:0]   io_pipe_phv_in_data_285,
  input  [7:0]   io_pipe_phv_in_data_286,
  input  [7:0]   io_pipe_phv_in_data_287,
  input  [7:0]   io_pipe_phv_in_data_288,
  input  [7:0]   io_pipe_phv_in_data_289,
  input  [7:0]   io_pipe_phv_in_data_290,
  input  [7:0]   io_pipe_phv_in_data_291,
  input  [7:0]   io_pipe_phv_in_data_292,
  input  [7:0]   io_pipe_phv_in_data_293,
  input  [7:0]   io_pipe_phv_in_data_294,
  input  [7:0]   io_pipe_phv_in_data_295,
  input  [7:0]   io_pipe_phv_in_data_296,
  input  [7:0]   io_pipe_phv_in_data_297,
  input  [7:0]   io_pipe_phv_in_data_298,
  input  [7:0]   io_pipe_phv_in_data_299,
  input  [7:0]   io_pipe_phv_in_data_300,
  input  [7:0]   io_pipe_phv_in_data_301,
  input  [7:0]   io_pipe_phv_in_data_302,
  input  [7:0]   io_pipe_phv_in_data_303,
  input  [7:0]   io_pipe_phv_in_data_304,
  input  [7:0]   io_pipe_phv_in_data_305,
  input  [7:0]   io_pipe_phv_in_data_306,
  input  [7:0]   io_pipe_phv_in_data_307,
  input  [7:0]   io_pipe_phv_in_data_308,
  input  [7:0]   io_pipe_phv_in_data_309,
  input  [7:0]   io_pipe_phv_in_data_310,
  input  [7:0]   io_pipe_phv_in_data_311,
  input  [7:0]   io_pipe_phv_in_data_312,
  input  [7:0]   io_pipe_phv_in_data_313,
  input  [7:0]   io_pipe_phv_in_data_314,
  input  [7:0]   io_pipe_phv_in_data_315,
  input  [7:0]   io_pipe_phv_in_data_316,
  input  [7:0]   io_pipe_phv_in_data_317,
  input  [7:0]   io_pipe_phv_in_data_318,
  input  [7:0]   io_pipe_phv_in_data_319,
  input  [7:0]   io_pipe_phv_in_data_320,
  input  [7:0]   io_pipe_phv_in_data_321,
  input  [7:0]   io_pipe_phv_in_data_322,
  input  [7:0]   io_pipe_phv_in_data_323,
  input  [7:0]   io_pipe_phv_in_data_324,
  input  [7:0]   io_pipe_phv_in_data_325,
  input  [7:0]   io_pipe_phv_in_data_326,
  input  [7:0]   io_pipe_phv_in_data_327,
  input  [7:0]   io_pipe_phv_in_data_328,
  input  [7:0]   io_pipe_phv_in_data_329,
  input  [7:0]   io_pipe_phv_in_data_330,
  input  [7:0]   io_pipe_phv_in_data_331,
  input  [7:0]   io_pipe_phv_in_data_332,
  input  [7:0]   io_pipe_phv_in_data_333,
  input  [7:0]   io_pipe_phv_in_data_334,
  input  [7:0]   io_pipe_phv_in_data_335,
  input  [7:0]   io_pipe_phv_in_data_336,
  input  [7:0]   io_pipe_phv_in_data_337,
  input  [7:0]   io_pipe_phv_in_data_338,
  input  [7:0]   io_pipe_phv_in_data_339,
  input  [7:0]   io_pipe_phv_in_data_340,
  input  [7:0]   io_pipe_phv_in_data_341,
  input  [7:0]   io_pipe_phv_in_data_342,
  input  [7:0]   io_pipe_phv_in_data_343,
  input  [7:0]   io_pipe_phv_in_data_344,
  input  [7:0]   io_pipe_phv_in_data_345,
  input  [7:0]   io_pipe_phv_in_data_346,
  input  [7:0]   io_pipe_phv_in_data_347,
  input  [7:0]   io_pipe_phv_in_data_348,
  input  [7:0]   io_pipe_phv_in_data_349,
  input  [7:0]   io_pipe_phv_in_data_350,
  input  [7:0]   io_pipe_phv_in_data_351,
  input  [7:0]   io_pipe_phv_in_data_352,
  input  [7:0]   io_pipe_phv_in_data_353,
  input  [7:0]   io_pipe_phv_in_data_354,
  input  [7:0]   io_pipe_phv_in_data_355,
  input  [7:0]   io_pipe_phv_in_data_356,
  input  [7:0]   io_pipe_phv_in_data_357,
  input  [7:0]   io_pipe_phv_in_data_358,
  input  [7:0]   io_pipe_phv_in_data_359,
  input  [7:0]   io_pipe_phv_in_data_360,
  input  [7:0]   io_pipe_phv_in_data_361,
  input  [7:0]   io_pipe_phv_in_data_362,
  input  [7:0]   io_pipe_phv_in_data_363,
  input  [7:0]   io_pipe_phv_in_data_364,
  input  [7:0]   io_pipe_phv_in_data_365,
  input  [7:0]   io_pipe_phv_in_data_366,
  input  [7:0]   io_pipe_phv_in_data_367,
  input  [7:0]   io_pipe_phv_in_data_368,
  input  [7:0]   io_pipe_phv_in_data_369,
  input  [7:0]   io_pipe_phv_in_data_370,
  input  [7:0]   io_pipe_phv_in_data_371,
  input  [7:0]   io_pipe_phv_in_data_372,
  input  [7:0]   io_pipe_phv_in_data_373,
  input  [7:0]   io_pipe_phv_in_data_374,
  input  [7:0]   io_pipe_phv_in_data_375,
  input  [7:0]   io_pipe_phv_in_data_376,
  input  [7:0]   io_pipe_phv_in_data_377,
  input  [7:0]   io_pipe_phv_in_data_378,
  input  [7:0]   io_pipe_phv_in_data_379,
  input  [7:0]   io_pipe_phv_in_data_380,
  input  [7:0]   io_pipe_phv_in_data_381,
  input  [7:0]   io_pipe_phv_in_data_382,
  input  [7:0]   io_pipe_phv_in_data_383,
  input  [7:0]   io_pipe_phv_in_data_384,
  input  [7:0]   io_pipe_phv_in_data_385,
  input  [7:0]   io_pipe_phv_in_data_386,
  input  [7:0]   io_pipe_phv_in_data_387,
  input  [7:0]   io_pipe_phv_in_data_388,
  input  [7:0]   io_pipe_phv_in_data_389,
  input  [7:0]   io_pipe_phv_in_data_390,
  input  [7:0]   io_pipe_phv_in_data_391,
  input  [7:0]   io_pipe_phv_in_data_392,
  input  [7:0]   io_pipe_phv_in_data_393,
  input  [7:0]   io_pipe_phv_in_data_394,
  input  [7:0]   io_pipe_phv_in_data_395,
  input  [7:0]   io_pipe_phv_in_data_396,
  input  [7:0]   io_pipe_phv_in_data_397,
  input  [7:0]   io_pipe_phv_in_data_398,
  input  [7:0]   io_pipe_phv_in_data_399,
  input  [7:0]   io_pipe_phv_in_data_400,
  input  [7:0]   io_pipe_phv_in_data_401,
  input  [7:0]   io_pipe_phv_in_data_402,
  input  [7:0]   io_pipe_phv_in_data_403,
  input  [7:0]   io_pipe_phv_in_data_404,
  input  [7:0]   io_pipe_phv_in_data_405,
  input  [7:0]   io_pipe_phv_in_data_406,
  input  [7:0]   io_pipe_phv_in_data_407,
  input  [7:0]   io_pipe_phv_in_data_408,
  input  [7:0]   io_pipe_phv_in_data_409,
  input  [7:0]   io_pipe_phv_in_data_410,
  input  [7:0]   io_pipe_phv_in_data_411,
  input  [7:0]   io_pipe_phv_in_data_412,
  input  [7:0]   io_pipe_phv_in_data_413,
  input  [7:0]   io_pipe_phv_in_data_414,
  input  [7:0]   io_pipe_phv_in_data_415,
  input  [7:0]   io_pipe_phv_in_data_416,
  input  [7:0]   io_pipe_phv_in_data_417,
  input  [7:0]   io_pipe_phv_in_data_418,
  input  [7:0]   io_pipe_phv_in_data_419,
  input  [7:0]   io_pipe_phv_in_data_420,
  input  [7:0]   io_pipe_phv_in_data_421,
  input  [7:0]   io_pipe_phv_in_data_422,
  input  [7:0]   io_pipe_phv_in_data_423,
  input  [7:0]   io_pipe_phv_in_data_424,
  input  [7:0]   io_pipe_phv_in_data_425,
  input  [7:0]   io_pipe_phv_in_data_426,
  input  [7:0]   io_pipe_phv_in_data_427,
  input  [7:0]   io_pipe_phv_in_data_428,
  input  [7:0]   io_pipe_phv_in_data_429,
  input  [7:0]   io_pipe_phv_in_data_430,
  input  [7:0]   io_pipe_phv_in_data_431,
  input  [7:0]   io_pipe_phv_in_data_432,
  input  [7:0]   io_pipe_phv_in_data_433,
  input  [7:0]   io_pipe_phv_in_data_434,
  input  [7:0]   io_pipe_phv_in_data_435,
  input  [7:0]   io_pipe_phv_in_data_436,
  input  [7:0]   io_pipe_phv_in_data_437,
  input  [7:0]   io_pipe_phv_in_data_438,
  input  [7:0]   io_pipe_phv_in_data_439,
  input  [7:0]   io_pipe_phv_in_data_440,
  input  [7:0]   io_pipe_phv_in_data_441,
  input  [7:0]   io_pipe_phv_in_data_442,
  input  [7:0]   io_pipe_phv_in_data_443,
  input  [7:0]   io_pipe_phv_in_data_444,
  input  [7:0]   io_pipe_phv_in_data_445,
  input  [7:0]   io_pipe_phv_in_data_446,
  input  [7:0]   io_pipe_phv_in_data_447,
  input  [7:0]   io_pipe_phv_in_data_448,
  input  [7:0]   io_pipe_phv_in_data_449,
  input  [7:0]   io_pipe_phv_in_data_450,
  input  [7:0]   io_pipe_phv_in_data_451,
  input  [7:0]   io_pipe_phv_in_data_452,
  input  [7:0]   io_pipe_phv_in_data_453,
  input  [7:0]   io_pipe_phv_in_data_454,
  input  [7:0]   io_pipe_phv_in_data_455,
  input  [7:0]   io_pipe_phv_in_data_456,
  input  [7:0]   io_pipe_phv_in_data_457,
  input  [7:0]   io_pipe_phv_in_data_458,
  input  [7:0]   io_pipe_phv_in_data_459,
  input  [7:0]   io_pipe_phv_in_data_460,
  input  [7:0]   io_pipe_phv_in_data_461,
  input  [7:0]   io_pipe_phv_in_data_462,
  input  [7:0]   io_pipe_phv_in_data_463,
  input  [7:0]   io_pipe_phv_in_data_464,
  input  [7:0]   io_pipe_phv_in_data_465,
  input  [7:0]   io_pipe_phv_in_data_466,
  input  [7:0]   io_pipe_phv_in_data_467,
  input  [7:0]   io_pipe_phv_in_data_468,
  input  [7:0]   io_pipe_phv_in_data_469,
  input  [7:0]   io_pipe_phv_in_data_470,
  input  [7:0]   io_pipe_phv_in_data_471,
  input  [7:0]   io_pipe_phv_in_data_472,
  input  [7:0]   io_pipe_phv_in_data_473,
  input  [7:0]   io_pipe_phv_in_data_474,
  input  [7:0]   io_pipe_phv_in_data_475,
  input  [7:0]   io_pipe_phv_in_data_476,
  input  [7:0]   io_pipe_phv_in_data_477,
  input  [7:0]   io_pipe_phv_in_data_478,
  input  [7:0]   io_pipe_phv_in_data_479,
  input  [7:0]   io_pipe_phv_in_data_480,
  input  [7:0]   io_pipe_phv_in_data_481,
  input  [7:0]   io_pipe_phv_in_data_482,
  input  [7:0]   io_pipe_phv_in_data_483,
  input  [7:0]   io_pipe_phv_in_data_484,
  input  [7:0]   io_pipe_phv_in_data_485,
  input  [7:0]   io_pipe_phv_in_data_486,
  input  [7:0]   io_pipe_phv_in_data_487,
  input  [7:0]   io_pipe_phv_in_data_488,
  input  [7:0]   io_pipe_phv_in_data_489,
  input  [7:0]   io_pipe_phv_in_data_490,
  input  [7:0]   io_pipe_phv_in_data_491,
  input  [7:0]   io_pipe_phv_in_data_492,
  input  [7:0]   io_pipe_phv_in_data_493,
  input  [7:0]   io_pipe_phv_in_data_494,
  input  [7:0]   io_pipe_phv_in_data_495,
  input  [7:0]   io_pipe_phv_in_data_496,
  input  [7:0]   io_pipe_phv_in_data_497,
  input  [7:0]   io_pipe_phv_in_data_498,
  input  [7:0]   io_pipe_phv_in_data_499,
  input  [7:0]   io_pipe_phv_in_data_500,
  input  [7:0]   io_pipe_phv_in_data_501,
  input  [7:0]   io_pipe_phv_in_data_502,
  input  [7:0]   io_pipe_phv_in_data_503,
  input  [7:0]   io_pipe_phv_in_data_504,
  input  [7:0]   io_pipe_phv_in_data_505,
  input  [7:0]   io_pipe_phv_in_data_506,
  input  [7:0]   io_pipe_phv_in_data_507,
  input  [7:0]   io_pipe_phv_in_data_508,
  input  [7:0]   io_pipe_phv_in_data_509,
  input  [7:0]   io_pipe_phv_in_data_510,
  input  [7:0]   io_pipe_phv_in_data_511,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [7:0]   io_pipe_phv_out_data_160,
  output [7:0]   io_pipe_phv_out_data_161,
  output [7:0]   io_pipe_phv_out_data_162,
  output [7:0]   io_pipe_phv_out_data_163,
  output [7:0]   io_pipe_phv_out_data_164,
  output [7:0]   io_pipe_phv_out_data_165,
  output [7:0]   io_pipe_phv_out_data_166,
  output [7:0]   io_pipe_phv_out_data_167,
  output [7:0]   io_pipe_phv_out_data_168,
  output [7:0]   io_pipe_phv_out_data_169,
  output [7:0]   io_pipe_phv_out_data_170,
  output [7:0]   io_pipe_phv_out_data_171,
  output [7:0]   io_pipe_phv_out_data_172,
  output [7:0]   io_pipe_phv_out_data_173,
  output [7:0]   io_pipe_phv_out_data_174,
  output [7:0]   io_pipe_phv_out_data_175,
  output [7:0]   io_pipe_phv_out_data_176,
  output [7:0]   io_pipe_phv_out_data_177,
  output [7:0]   io_pipe_phv_out_data_178,
  output [7:0]   io_pipe_phv_out_data_179,
  output [7:0]   io_pipe_phv_out_data_180,
  output [7:0]   io_pipe_phv_out_data_181,
  output [7:0]   io_pipe_phv_out_data_182,
  output [7:0]   io_pipe_phv_out_data_183,
  output [7:0]   io_pipe_phv_out_data_184,
  output [7:0]   io_pipe_phv_out_data_185,
  output [7:0]   io_pipe_phv_out_data_186,
  output [7:0]   io_pipe_phv_out_data_187,
  output [7:0]   io_pipe_phv_out_data_188,
  output [7:0]   io_pipe_phv_out_data_189,
  output [7:0]   io_pipe_phv_out_data_190,
  output [7:0]   io_pipe_phv_out_data_191,
  output [7:0]   io_pipe_phv_out_data_192,
  output [7:0]   io_pipe_phv_out_data_193,
  output [7:0]   io_pipe_phv_out_data_194,
  output [7:0]   io_pipe_phv_out_data_195,
  output [7:0]   io_pipe_phv_out_data_196,
  output [7:0]   io_pipe_phv_out_data_197,
  output [7:0]   io_pipe_phv_out_data_198,
  output [7:0]   io_pipe_phv_out_data_199,
  output [7:0]   io_pipe_phv_out_data_200,
  output [7:0]   io_pipe_phv_out_data_201,
  output [7:0]   io_pipe_phv_out_data_202,
  output [7:0]   io_pipe_phv_out_data_203,
  output [7:0]   io_pipe_phv_out_data_204,
  output [7:0]   io_pipe_phv_out_data_205,
  output [7:0]   io_pipe_phv_out_data_206,
  output [7:0]   io_pipe_phv_out_data_207,
  output [7:0]   io_pipe_phv_out_data_208,
  output [7:0]   io_pipe_phv_out_data_209,
  output [7:0]   io_pipe_phv_out_data_210,
  output [7:0]   io_pipe_phv_out_data_211,
  output [7:0]   io_pipe_phv_out_data_212,
  output [7:0]   io_pipe_phv_out_data_213,
  output [7:0]   io_pipe_phv_out_data_214,
  output [7:0]   io_pipe_phv_out_data_215,
  output [7:0]   io_pipe_phv_out_data_216,
  output [7:0]   io_pipe_phv_out_data_217,
  output [7:0]   io_pipe_phv_out_data_218,
  output [7:0]   io_pipe_phv_out_data_219,
  output [7:0]   io_pipe_phv_out_data_220,
  output [7:0]   io_pipe_phv_out_data_221,
  output [7:0]   io_pipe_phv_out_data_222,
  output [7:0]   io_pipe_phv_out_data_223,
  output [7:0]   io_pipe_phv_out_data_224,
  output [7:0]   io_pipe_phv_out_data_225,
  output [7:0]   io_pipe_phv_out_data_226,
  output [7:0]   io_pipe_phv_out_data_227,
  output [7:0]   io_pipe_phv_out_data_228,
  output [7:0]   io_pipe_phv_out_data_229,
  output [7:0]   io_pipe_phv_out_data_230,
  output [7:0]   io_pipe_phv_out_data_231,
  output [7:0]   io_pipe_phv_out_data_232,
  output [7:0]   io_pipe_phv_out_data_233,
  output [7:0]   io_pipe_phv_out_data_234,
  output [7:0]   io_pipe_phv_out_data_235,
  output [7:0]   io_pipe_phv_out_data_236,
  output [7:0]   io_pipe_phv_out_data_237,
  output [7:0]   io_pipe_phv_out_data_238,
  output [7:0]   io_pipe_phv_out_data_239,
  output [7:0]   io_pipe_phv_out_data_240,
  output [7:0]   io_pipe_phv_out_data_241,
  output [7:0]   io_pipe_phv_out_data_242,
  output [7:0]   io_pipe_phv_out_data_243,
  output [7:0]   io_pipe_phv_out_data_244,
  output [7:0]   io_pipe_phv_out_data_245,
  output [7:0]   io_pipe_phv_out_data_246,
  output [7:0]   io_pipe_phv_out_data_247,
  output [7:0]   io_pipe_phv_out_data_248,
  output [7:0]   io_pipe_phv_out_data_249,
  output [7:0]   io_pipe_phv_out_data_250,
  output [7:0]   io_pipe_phv_out_data_251,
  output [7:0]   io_pipe_phv_out_data_252,
  output [7:0]   io_pipe_phv_out_data_253,
  output [7:0]   io_pipe_phv_out_data_254,
  output [7:0]   io_pipe_phv_out_data_255,
  output [7:0]   io_pipe_phv_out_data_256,
  output [7:0]   io_pipe_phv_out_data_257,
  output [7:0]   io_pipe_phv_out_data_258,
  output [7:0]   io_pipe_phv_out_data_259,
  output [7:0]   io_pipe_phv_out_data_260,
  output [7:0]   io_pipe_phv_out_data_261,
  output [7:0]   io_pipe_phv_out_data_262,
  output [7:0]   io_pipe_phv_out_data_263,
  output [7:0]   io_pipe_phv_out_data_264,
  output [7:0]   io_pipe_phv_out_data_265,
  output [7:0]   io_pipe_phv_out_data_266,
  output [7:0]   io_pipe_phv_out_data_267,
  output [7:0]   io_pipe_phv_out_data_268,
  output [7:0]   io_pipe_phv_out_data_269,
  output [7:0]   io_pipe_phv_out_data_270,
  output [7:0]   io_pipe_phv_out_data_271,
  output [7:0]   io_pipe_phv_out_data_272,
  output [7:0]   io_pipe_phv_out_data_273,
  output [7:0]   io_pipe_phv_out_data_274,
  output [7:0]   io_pipe_phv_out_data_275,
  output [7:0]   io_pipe_phv_out_data_276,
  output [7:0]   io_pipe_phv_out_data_277,
  output [7:0]   io_pipe_phv_out_data_278,
  output [7:0]   io_pipe_phv_out_data_279,
  output [7:0]   io_pipe_phv_out_data_280,
  output [7:0]   io_pipe_phv_out_data_281,
  output [7:0]   io_pipe_phv_out_data_282,
  output [7:0]   io_pipe_phv_out_data_283,
  output [7:0]   io_pipe_phv_out_data_284,
  output [7:0]   io_pipe_phv_out_data_285,
  output [7:0]   io_pipe_phv_out_data_286,
  output [7:0]   io_pipe_phv_out_data_287,
  output [7:0]   io_pipe_phv_out_data_288,
  output [7:0]   io_pipe_phv_out_data_289,
  output [7:0]   io_pipe_phv_out_data_290,
  output [7:0]   io_pipe_phv_out_data_291,
  output [7:0]   io_pipe_phv_out_data_292,
  output [7:0]   io_pipe_phv_out_data_293,
  output [7:0]   io_pipe_phv_out_data_294,
  output [7:0]   io_pipe_phv_out_data_295,
  output [7:0]   io_pipe_phv_out_data_296,
  output [7:0]   io_pipe_phv_out_data_297,
  output [7:0]   io_pipe_phv_out_data_298,
  output [7:0]   io_pipe_phv_out_data_299,
  output [7:0]   io_pipe_phv_out_data_300,
  output [7:0]   io_pipe_phv_out_data_301,
  output [7:0]   io_pipe_phv_out_data_302,
  output [7:0]   io_pipe_phv_out_data_303,
  output [7:0]   io_pipe_phv_out_data_304,
  output [7:0]   io_pipe_phv_out_data_305,
  output [7:0]   io_pipe_phv_out_data_306,
  output [7:0]   io_pipe_phv_out_data_307,
  output [7:0]   io_pipe_phv_out_data_308,
  output [7:0]   io_pipe_phv_out_data_309,
  output [7:0]   io_pipe_phv_out_data_310,
  output [7:0]   io_pipe_phv_out_data_311,
  output [7:0]   io_pipe_phv_out_data_312,
  output [7:0]   io_pipe_phv_out_data_313,
  output [7:0]   io_pipe_phv_out_data_314,
  output [7:0]   io_pipe_phv_out_data_315,
  output [7:0]   io_pipe_phv_out_data_316,
  output [7:0]   io_pipe_phv_out_data_317,
  output [7:0]   io_pipe_phv_out_data_318,
  output [7:0]   io_pipe_phv_out_data_319,
  output [7:0]   io_pipe_phv_out_data_320,
  output [7:0]   io_pipe_phv_out_data_321,
  output [7:0]   io_pipe_phv_out_data_322,
  output [7:0]   io_pipe_phv_out_data_323,
  output [7:0]   io_pipe_phv_out_data_324,
  output [7:0]   io_pipe_phv_out_data_325,
  output [7:0]   io_pipe_phv_out_data_326,
  output [7:0]   io_pipe_phv_out_data_327,
  output [7:0]   io_pipe_phv_out_data_328,
  output [7:0]   io_pipe_phv_out_data_329,
  output [7:0]   io_pipe_phv_out_data_330,
  output [7:0]   io_pipe_phv_out_data_331,
  output [7:0]   io_pipe_phv_out_data_332,
  output [7:0]   io_pipe_phv_out_data_333,
  output [7:0]   io_pipe_phv_out_data_334,
  output [7:0]   io_pipe_phv_out_data_335,
  output [7:0]   io_pipe_phv_out_data_336,
  output [7:0]   io_pipe_phv_out_data_337,
  output [7:0]   io_pipe_phv_out_data_338,
  output [7:0]   io_pipe_phv_out_data_339,
  output [7:0]   io_pipe_phv_out_data_340,
  output [7:0]   io_pipe_phv_out_data_341,
  output [7:0]   io_pipe_phv_out_data_342,
  output [7:0]   io_pipe_phv_out_data_343,
  output [7:0]   io_pipe_phv_out_data_344,
  output [7:0]   io_pipe_phv_out_data_345,
  output [7:0]   io_pipe_phv_out_data_346,
  output [7:0]   io_pipe_phv_out_data_347,
  output [7:0]   io_pipe_phv_out_data_348,
  output [7:0]   io_pipe_phv_out_data_349,
  output [7:0]   io_pipe_phv_out_data_350,
  output [7:0]   io_pipe_phv_out_data_351,
  output [7:0]   io_pipe_phv_out_data_352,
  output [7:0]   io_pipe_phv_out_data_353,
  output [7:0]   io_pipe_phv_out_data_354,
  output [7:0]   io_pipe_phv_out_data_355,
  output [7:0]   io_pipe_phv_out_data_356,
  output [7:0]   io_pipe_phv_out_data_357,
  output [7:0]   io_pipe_phv_out_data_358,
  output [7:0]   io_pipe_phv_out_data_359,
  output [7:0]   io_pipe_phv_out_data_360,
  output [7:0]   io_pipe_phv_out_data_361,
  output [7:0]   io_pipe_phv_out_data_362,
  output [7:0]   io_pipe_phv_out_data_363,
  output [7:0]   io_pipe_phv_out_data_364,
  output [7:0]   io_pipe_phv_out_data_365,
  output [7:0]   io_pipe_phv_out_data_366,
  output [7:0]   io_pipe_phv_out_data_367,
  output [7:0]   io_pipe_phv_out_data_368,
  output [7:0]   io_pipe_phv_out_data_369,
  output [7:0]   io_pipe_phv_out_data_370,
  output [7:0]   io_pipe_phv_out_data_371,
  output [7:0]   io_pipe_phv_out_data_372,
  output [7:0]   io_pipe_phv_out_data_373,
  output [7:0]   io_pipe_phv_out_data_374,
  output [7:0]   io_pipe_phv_out_data_375,
  output [7:0]   io_pipe_phv_out_data_376,
  output [7:0]   io_pipe_phv_out_data_377,
  output [7:0]   io_pipe_phv_out_data_378,
  output [7:0]   io_pipe_phv_out_data_379,
  output [7:0]   io_pipe_phv_out_data_380,
  output [7:0]   io_pipe_phv_out_data_381,
  output [7:0]   io_pipe_phv_out_data_382,
  output [7:0]   io_pipe_phv_out_data_383,
  output [7:0]   io_pipe_phv_out_data_384,
  output [7:0]   io_pipe_phv_out_data_385,
  output [7:0]   io_pipe_phv_out_data_386,
  output [7:0]   io_pipe_phv_out_data_387,
  output [7:0]   io_pipe_phv_out_data_388,
  output [7:0]   io_pipe_phv_out_data_389,
  output [7:0]   io_pipe_phv_out_data_390,
  output [7:0]   io_pipe_phv_out_data_391,
  output [7:0]   io_pipe_phv_out_data_392,
  output [7:0]   io_pipe_phv_out_data_393,
  output [7:0]   io_pipe_phv_out_data_394,
  output [7:0]   io_pipe_phv_out_data_395,
  output [7:0]   io_pipe_phv_out_data_396,
  output [7:0]   io_pipe_phv_out_data_397,
  output [7:0]   io_pipe_phv_out_data_398,
  output [7:0]   io_pipe_phv_out_data_399,
  output [7:0]   io_pipe_phv_out_data_400,
  output [7:0]   io_pipe_phv_out_data_401,
  output [7:0]   io_pipe_phv_out_data_402,
  output [7:0]   io_pipe_phv_out_data_403,
  output [7:0]   io_pipe_phv_out_data_404,
  output [7:0]   io_pipe_phv_out_data_405,
  output [7:0]   io_pipe_phv_out_data_406,
  output [7:0]   io_pipe_phv_out_data_407,
  output [7:0]   io_pipe_phv_out_data_408,
  output [7:0]   io_pipe_phv_out_data_409,
  output [7:0]   io_pipe_phv_out_data_410,
  output [7:0]   io_pipe_phv_out_data_411,
  output [7:0]   io_pipe_phv_out_data_412,
  output [7:0]   io_pipe_phv_out_data_413,
  output [7:0]   io_pipe_phv_out_data_414,
  output [7:0]   io_pipe_phv_out_data_415,
  output [7:0]   io_pipe_phv_out_data_416,
  output [7:0]   io_pipe_phv_out_data_417,
  output [7:0]   io_pipe_phv_out_data_418,
  output [7:0]   io_pipe_phv_out_data_419,
  output [7:0]   io_pipe_phv_out_data_420,
  output [7:0]   io_pipe_phv_out_data_421,
  output [7:0]   io_pipe_phv_out_data_422,
  output [7:0]   io_pipe_phv_out_data_423,
  output [7:0]   io_pipe_phv_out_data_424,
  output [7:0]   io_pipe_phv_out_data_425,
  output [7:0]   io_pipe_phv_out_data_426,
  output [7:0]   io_pipe_phv_out_data_427,
  output [7:0]   io_pipe_phv_out_data_428,
  output [7:0]   io_pipe_phv_out_data_429,
  output [7:0]   io_pipe_phv_out_data_430,
  output [7:0]   io_pipe_phv_out_data_431,
  output [7:0]   io_pipe_phv_out_data_432,
  output [7:0]   io_pipe_phv_out_data_433,
  output [7:0]   io_pipe_phv_out_data_434,
  output [7:0]   io_pipe_phv_out_data_435,
  output [7:0]   io_pipe_phv_out_data_436,
  output [7:0]   io_pipe_phv_out_data_437,
  output [7:0]   io_pipe_phv_out_data_438,
  output [7:0]   io_pipe_phv_out_data_439,
  output [7:0]   io_pipe_phv_out_data_440,
  output [7:0]   io_pipe_phv_out_data_441,
  output [7:0]   io_pipe_phv_out_data_442,
  output [7:0]   io_pipe_phv_out_data_443,
  output [7:0]   io_pipe_phv_out_data_444,
  output [7:0]   io_pipe_phv_out_data_445,
  output [7:0]   io_pipe_phv_out_data_446,
  output [7:0]   io_pipe_phv_out_data_447,
  output [7:0]   io_pipe_phv_out_data_448,
  output [7:0]   io_pipe_phv_out_data_449,
  output [7:0]   io_pipe_phv_out_data_450,
  output [7:0]   io_pipe_phv_out_data_451,
  output [7:0]   io_pipe_phv_out_data_452,
  output [7:0]   io_pipe_phv_out_data_453,
  output [7:0]   io_pipe_phv_out_data_454,
  output [7:0]   io_pipe_phv_out_data_455,
  output [7:0]   io_pipe_phv_out_data_456,
  output [7:0]   io_pipe_phv_out_data_457,
  output [7:0]   io_pipe_phv_out_data_458,
  output [7:0]   io_pipe_phv_out_data_459,
  output [7:0]   io_pipe_phv_out_data_460,
  output [7:0]   io_pipe_phv_out_data_461,
  output [7:0]   io_pipe_phv_out_data_462,
  output [7:0]   io_pipe_phv_out_data_463,
  output [7:0]   io_pipe_phv_out_data_464,
  output [7:0]   io_pipe_phv_out_data_465,
  output [7:0]   io_pipe_phv_out_data_466,
  output [7:0]   io_pipe_phv_out_data_467,
  output [7:0]   io_pipe_phv_out_data_468,
  output [7:0]   io_pipe_phv_out_data_469,
  output [7:0]   io_pipe_phv_out_data_470,
  output [7:0]   io_pipe_phv_out_data_471,
  output [7:0]   io_pipe_phv_out_data_472,
  output [7:0]   io_pipe_phv_out_data_473,
  output [7:0]   io_pipe_phv_out_data_474,
  output [7:0]   io_pipe_phv_out_data_475,
  output [7:0]   io_pipe_phv_out_data_476,
  output [7:0]   io_pipe_phv_out_data_477,
  output [7:0]   io_pipe_phv_out_data_478,
  output [7:0]   io_pipe_phv_out_data_479,
  output [7:0]   io_pipe_phv_out_data_480,
  output [7:0]   io_pipe_phv_out_data_481,
  output [7:0]   io_pipe_phv_out_data_482,
  output [7:0]   io_pipe_phv_out_data_483,
  output [7:0]   io_pipe_phv_out_data_484,
  output [7:0]   io_pipe_phv_out_data_485,
  output [7:0]   io_pipe_phv_out_data_486,
  output [7:0]   io_pipe_phv_out_data_487,
  output [7:0]   io_pipe_phv_out_data_488,
  output [7:0]   io_pipe_phv_out_data_489,
  output [7:0]   io_pipe_phv_out_data_490,
  output [7:0]   io_pipe_phv_out_data_491,
  output [7:0]   io_pipe_phv_out_data_492,
  output [7:0]   io_pipe_phv_out_data_493,
  output [7:0]   io_pipe_phv_out_data_494,
  output [7:0]   io_pipe_phv_out_data_495,
  output [7:0]   io_pipe_phv_out_data_496,
  output [7:0]   io_pipe_phv_out_data_497,
  output [7:0]   io_pipe_phv_out_data_498,
  output [7:0]   io_pipe_phv_out_data_499,
  output [7:0]   io_pipe_phv_out_data_500,
  output [7:0]   io_pipe_phv_out_data_501,
  output [7:0]   io_pipe_phv_out_data_502,
  output [7:0]   io_pipe_phv_out_data_503,
  output [7:0]   io_pipe_phv_out_data_504,
  output [7:0]   io_pipe_phv_out_data_505,
  output [7:0]   io_pipe_phv_out_data_506,
  output [7:0]   io_pipe_phv_out_data_507,
  output [7:0]   io_pipe_phv_out_data_508,
  output [7:0]   io_pipe_phv_out_data_509,
  output [7:0]   io_pipe_phv_out_data_510,
  output [7:0]   io_pipe_phv_out_data_511,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input          io_mod_hash_depth_mod,
  input          io_mod_config_id,
  input  [3:0]   io_mod_hash_depth,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  output [7:0]   io_hash_val,
  output [3:0]   io_hash_val_cs
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_256; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_257; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_258; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_259; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_260; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_261; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_262; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_263; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_264; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_265; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_266; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_267; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_268; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_269; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_270; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_271; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_272; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_273; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_274; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_275; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_276; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_277; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_278; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_279; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_280; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_281; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_282; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_283; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_284; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_285; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_286; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_287; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_288; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_289; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_290; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_291; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_292; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_293; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_294; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_295; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_296; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_297; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_298; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_299; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_300; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_301; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_302; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_303; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_304; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_305; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_306; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_307; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_308; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_309; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_310; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_311; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_312; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_313; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_314; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_315; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_316; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_317; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_318; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_319; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_320; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_321; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_322; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_323; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_324; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_325; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_326; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_327; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_328; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_329; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_330; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_331; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_332; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_333; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_334; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_335; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_336; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_337; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_338; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_339; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_340; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_341; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_342; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_343; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_344; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_345; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_346; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_347; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_348; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_349; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_350; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_351; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_352; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_353; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_354; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_355; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_356; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_357; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_358; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_359; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_360; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_361; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_362; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_363; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_364; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_365; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_366; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_367; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_368; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_369; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_370; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_371; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_372; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_373; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_374; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_375; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_376; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_377; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_378; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_379; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_380; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_381; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_382; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_383; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_384; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_385; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_386; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_387; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_388; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_389; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_390; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_391; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_392; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_393; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_394; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_395; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_396; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_397; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_398; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_399; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_400; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_401; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_402; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_403; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_404; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_405; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_406; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_407; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_408; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_409; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_410; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_411; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_412; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_413; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_414; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_415; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_416; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_417; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_418; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_419; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_420; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_421; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_422; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_423; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_424; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_425; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_426; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_427; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_428; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_429; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_430; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_431; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_432; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_433; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_434; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_435; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_436; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_437; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_438; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_439; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_440; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_441; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_442; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_443; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_444; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_445; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_446; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_447; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_448; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_449; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_450; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_451; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_452; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_453; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_454; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_455; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_456; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_457; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_458; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_459; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_460; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_461; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_462; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_463; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_464; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_465; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_466; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_467; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_468; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_469; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_470; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_471; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_472; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_473; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_474; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_475; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_476; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_477; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_478; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_479; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_480; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_481; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_482; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_483; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_484; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_485; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_486; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_487; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_488; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_489; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_490; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_491; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_492; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_493; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_494; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_495; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_496; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_497; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_498; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_499; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_500; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_501; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_502; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_503; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_504; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_505; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_506; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_507; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_508; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_509; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_510; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_511; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[hash.scala 127:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_256; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_257; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_258; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_259; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_260; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_261; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_262; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_263; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_264; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_265; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_266; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_267; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_268; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_269; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_270; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_271; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_272; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_273; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_274; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_275; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_276; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_277; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_278; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_279; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_280; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_281; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_282; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_283; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_284; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_285; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_286; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_287; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_288; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_289; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_290; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_291; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_292; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_293; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_294; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_295; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_296; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_297; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_298; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_299; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_300; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_301; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_302; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_303; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_304; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_305; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_306; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_307; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_308; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_309; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_310; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_311; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_312; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_313; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_314; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_315; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_316; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_317; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_318; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_319; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_320; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_321; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_322; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_323; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_324; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_325; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_326; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_327; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_328; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_329; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_330; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_331; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_332; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_333; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_334; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_335; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_336; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_337; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_338; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_339; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_340; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_341; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_342; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_343; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_344; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_345; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_346; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_347; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_348; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_349; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_350; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_351; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_352; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_353; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_354; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_355; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_356; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_357; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_358; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_359; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_360; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_361; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_362; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_363; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_364; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_365; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_366; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_367; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_368; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_369; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_370; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_371; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_372; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_373; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_374; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_375; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_376; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_377; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_378; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_379; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_380; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_381; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_382; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_383; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_384; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_385; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_386; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_387; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_388; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_389; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_390; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_391; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_392; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_393; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_394; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_395; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_396; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_397; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_398; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_399; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_400; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_401; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_402; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_403; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_404; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_405; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_406; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_407; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_408; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_409; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_410; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_411; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_412; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_413; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_414; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_415; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_416; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_417; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_418; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_419; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_420; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_421; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_422; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_423; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_424; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_425; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_426; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_427; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_428; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_429; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_430; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_431; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_432; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_433; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_434; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_435; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_436; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_437; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_438; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_439; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_440; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_441; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_442; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_443; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_444; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_445; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_446; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_447; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_448; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_449; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_450; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_451; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_452; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_453; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_454; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_455; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_456; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_457; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_458; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_459; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_460; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_461; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_462; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_463; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_464; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_465; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_466; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_467; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_468; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_469; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_470; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_471; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_472; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_473; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_474; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_475; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_476; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_477; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_478; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_479; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_480; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_481; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_482; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_483; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_484; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_485; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_486; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_487; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_488; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_489; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_490; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_491; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_492; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_493; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_494; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_495; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_496; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_497; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_498; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_499; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_500; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_501; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_502; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_503; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_504; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_505; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_506; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_507; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_508; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_509; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_510; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_511; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 127:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_key_in; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_key_out; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_sum_in; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_sum_out; // @[hash.scala 127:23]
  wire  pipe2_clock; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_256; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_257; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_258; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_259; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_260; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_261; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_262; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_263; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_264; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_265; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_266; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_267; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_268; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_269; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_270; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_271; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_272; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_273; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_274; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_275; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_276; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_277; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_278; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_279; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_280; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_281; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_282; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_283; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_284; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_285; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_286; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_287; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_288; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_289; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_290; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_291; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_292; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_293; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_294; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_295; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_296; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_297; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_298; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_299; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_300; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_301; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_302; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_303; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_304; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_305; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_306; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_307; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_308; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_309; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_310; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_311; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_312; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_313; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_314; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_315; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_316; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_317; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_318; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_319; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_320; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_321; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_322; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_323; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_324; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_325; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_326; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_327; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_328; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_329; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_330; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_331; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_332; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_333; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_334; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_335; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_336; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_337; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_338; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_339; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_340; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_341; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_342; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_343; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_344; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_345; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_346; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_347; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_348; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_349; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_350; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_351; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_352; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_353; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_354; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_355; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_356; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_357; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_358; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_359; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_360; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_361; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_362; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_363; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_364; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_365; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_366; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_367; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_368; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_369; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_370; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_371; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_372; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_373; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_374; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_375; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_376; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_377; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_378; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_379; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_380; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_381; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_382; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_383; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_384; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_385; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_386; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_387; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_388; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_389; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_390; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_391; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_392; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_393; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_394; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_395; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_396; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_397; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_398; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_399; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_400; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_401; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_402; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_403; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_404; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_405; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_406; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_407; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_408; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_409; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_410; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_411; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_412; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_413; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_414; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_415; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_416; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_417; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_418; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_419; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_420; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_421; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_422; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_423; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_424; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_425; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_426; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_427; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_428; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_429; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_430; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_431; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_432; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_433; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_434; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_435; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_436; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_437; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_438; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_439; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_440; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_441; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_442; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_443; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_444; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_445; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_446; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_447; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_448; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_449; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_450; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_451; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_452; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_453; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_454; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_455; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_456; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_457; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_458; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_459; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_460; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_461; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_462; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_463; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_464; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_465; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_466; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_467; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_468; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_469; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_470; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_471; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_472; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_473; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_474; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_475; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_476; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_477; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_478; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_479; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_480; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_481; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_482; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_483; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_484; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_485; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_486; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_487; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_488; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_489; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_490; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_491; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_492; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_493; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_494; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_495; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_496; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_497; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_498; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_499; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_500; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_501; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_502; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_503; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_504; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_505; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_506; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_507; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_508; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_509; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_510; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_511; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[hash.scala 128:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_256; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_257; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_258; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_259; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_260; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_261; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_262; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_263; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_264; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_265; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_266; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_267; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_268; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_269; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_270; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_271; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_272; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_273; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_274; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_275; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_276; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_277; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_278; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_279; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_280; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_281; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_282; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_283; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_284; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_285; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_286; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_287; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_288; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_289; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_290; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_291; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_292; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_293; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_294; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_295; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_296; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_297; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_298; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_299; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_300; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_301; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_302; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_303; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_304; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_305; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_306; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_307; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_308; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_309; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_310; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_311; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_312; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_313; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_314; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_315; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_316; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_317; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_318; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_319; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_320; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_321; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_322; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_323; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_324; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_325; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_326; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_327; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_328; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_329; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_330; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_331; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_332; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_333; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_334; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_335; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_336; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_337; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_338; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_339; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_340; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_341; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_342; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_343; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_344; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_345; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_346; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_347; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_348; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_349; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_350; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_351; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_352; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_353; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_354; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_355; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_356; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_357; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_358; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_359; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_360; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_361; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_362; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_363; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_364; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_365; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_366; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_367; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_368; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_369; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_370; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_371; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_372; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_373; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_374; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_375; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_376; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_377; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_378; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_379; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_380; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_381; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_382; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_383; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_384; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_385; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_386; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_387; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_388; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_389; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_390; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_391; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_392; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_393; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_394; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_395; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_396; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_397; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_398; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_399; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_400; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_401; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_402; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_403; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_404; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_405; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_406; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_407; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_408; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_409; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_410; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_411; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_412; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_413; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_414; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_415; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_416; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_417; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_418; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_419; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_420; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_421; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_422; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_423; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_424; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_425; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_426; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_427; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_428; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_429; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_430; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_431; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_432; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_433; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_434; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_435; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_436; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_437; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_438; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_439; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_440; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_441; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_442; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_443; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_444; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_445; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_446; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_447; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_448; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_449; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_450; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_451; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_452; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_453; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_454; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_455; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_456; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_457; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_458; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_459; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_460; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_461; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_462; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_463; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_464; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_465; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_466; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_467; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_468; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_469; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_470; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_471; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_472; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_473; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_474; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_475; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_476; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_477; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_478; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_479; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_480; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_481; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_482; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_483; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_484; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_485; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_486; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_487; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_488; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_489; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_490; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_491; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_492; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_493; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_494; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_495; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_496; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_497; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_498; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_499; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_500; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_501; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_502; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_503; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_504; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_505; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_506; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_507; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_508; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_509; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_510; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_511; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 128:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_key_in; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_key_out; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_sum_in; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_sum_out; // @[hash.scala 128:23]
  wire  pipe3_clock; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_160; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_161; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_162; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_163; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_164; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_165; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_166; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_167; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_168; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_169; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_170; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_171; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_172; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_173; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_174; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_175; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_176; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_177; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_178; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_179; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_180; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_181; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_182; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_183; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_184; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_185; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_186; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_187; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_188; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_189; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_190; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_191; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_192; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_193; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_194; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_195; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_196; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_197; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_198; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_199; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_200; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_201; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_202; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_203; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_204; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_205; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_206; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_207; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_208; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_209; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_210; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_211; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_212; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_213; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_214; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_215; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_216; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_217; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_218; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_219; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_220; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_221; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_222; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_223; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_224; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_225; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_226; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_227; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_228; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_229; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_230; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_231; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_232; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_233; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_234; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_235; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_236; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_237; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_238; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_239; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_240; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_241; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_242; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_243; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_244; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_245; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_246; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_247; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_248; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_249; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_250; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_251; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_252; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_253; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_254; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_255; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_256; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_257; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_258; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_259; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_260; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_261; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_262; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_263; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_264; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_265; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_266; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_267; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_268; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_269; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_270; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_271; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_272; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_273; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_274; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_275; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_276; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_277; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_278; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_279; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_280; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_281; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_282; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_283; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_284; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_285; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_286; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_287; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_288; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_289; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_290; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_291; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_292; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_293; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_294; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_295; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_296; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_297; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_298; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_299; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_300; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_301; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_302; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_303; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_304; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_305; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_306; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_307; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_308; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_309; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_310; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_311; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_312; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_313; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_314; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_315; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_316; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_317; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_318; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_319; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_320; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_321; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_322; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_323; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_324; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_325; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_326; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_327; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_328; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_329; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_330; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_331; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_332; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_333; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_334; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_335; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_336; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_337; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_338; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_339; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_340; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_341; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_342; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_343; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_344; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_345; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_346; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_347; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_348; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_349; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_350; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_351; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_352; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_353; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_354; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_355; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_356; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_357; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_358; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_359; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_360; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_361; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_362; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_363; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_364; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_365; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_366; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_367; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_368; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_369; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_370; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_371; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_372; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_373; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_374; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_375; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_376; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_377; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_378; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_379; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_380; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_381; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_382; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_383; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_384; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_385; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_386; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_387; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_388; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_389; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_390; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_391; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_392; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_393; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_394; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_395; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_396; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_397; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_398; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_399; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_400; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_401; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_402; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_403; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_404; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_405; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_406; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_407; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_408; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_409; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_410; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_411; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_412; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_413; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_414; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_415; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_416; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_417; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_418; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_419; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_420; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_421; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_422; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_423; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_424; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_425; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_426; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_427; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_428; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_429; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_430; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_431; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_432; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_433; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_434; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_435; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_436; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_437; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_438; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_439; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_440; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_441; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_442; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_443; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_444; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_445; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_446; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_447; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_448; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_449; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_450; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_451; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_452; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_453; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_454; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_455; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_456; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_457; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_458; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_459; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_460; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_461; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_462; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_463; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_464; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_465; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_466; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_467; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_468; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_469; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_470; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_471; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_472; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_473; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_474; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_475; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_476; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_477; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_478; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_479; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_480; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_481; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_482; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_483; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_484; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_485; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_486; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_487; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_488; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_489; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_490; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_491; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_492; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_493; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_494; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_495; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_496; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_497; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_498; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_499; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_500; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_501; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_502; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_503; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_504; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_505; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_506; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_507; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_508; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_509; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_510; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_511; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[hash.scala 129:23]
  wire [3:0] pipe3_io_pipe_phv_in_next_processor_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_160; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_161; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_162; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_163; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_164; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_165; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_166; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_167; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_168; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_169; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_170; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_171; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_172; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_173; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_174; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_175; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_176; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_177; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_178; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_179; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_180; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_181; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_182; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_183; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_184; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_185; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_186; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_187; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_188; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_189; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_190; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_191; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_192; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_193; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_194; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_195; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_196; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_197; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_198; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_199; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_200; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_201; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_202; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_203; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_204; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_205; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_206; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_207; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_208; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_209; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_210; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_211; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_212; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_213; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_214; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_215; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_216; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_217; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_218; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_219; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_220; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_221; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_222; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_223; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_224; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_225; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_226; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_227; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_228; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_229; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_230; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_231; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_232; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_233; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_234; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_235; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_236; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_237; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_238; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_239; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_240; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_241; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_242; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_243; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_244; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_245; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_246; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_247; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_248; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_249; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_250; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_251; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_252; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_253; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_254; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_255; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_256; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_257; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_258; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_259; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_260; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_261; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_262; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_263; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_264; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_265; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_266; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_267; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_268; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_269; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_270; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_271; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_272; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_273; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_274; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_275; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_276; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_277; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_278; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_279; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_280; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_281; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_282; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_283; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_284; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_285; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_286; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_287; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_288; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_289; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_290; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_291; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_292; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_293; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_294; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_295; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_296; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_297; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_298; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_299; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_300; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_301; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_302; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_303; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_304; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_305; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_306; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_307; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_308; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_309; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_310; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_311; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_312; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_313; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_314; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_315; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_316; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_317; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_318; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_319; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_320; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_321; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_322; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_323; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_324; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_325; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_326; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_327; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_328; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_329; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_330; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_331; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_332; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_333; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_334; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_335; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_336; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_337; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_338; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_339; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_340; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_341; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_342; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_343; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_344; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_345; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_346; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_347; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_348; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_349; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_350; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_351; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_352; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_353; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_354; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_355; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_356; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_357; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_358; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_359; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_360; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_361; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_362; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_363; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_364; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_365; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_366; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_367; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_368; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_369; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_370; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_371; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_372; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_373; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_374; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_375; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_376; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_377; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_378; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_379; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_380; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_381; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_382; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_383; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_384; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_385; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_386; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_387; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_388; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_389; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_390; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_391; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_392; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_393; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_394; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_395; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_396; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_397; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_398; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_399; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_400; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_401; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_402; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_403; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_404; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_405; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_406; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_407; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_408; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_409; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_410; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_411; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_412; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_413; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_414; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_415; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_416; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_417; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_418; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_419; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_420; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_421; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_422; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_423; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_424; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_425; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_426; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_427; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_428; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_429; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_430; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_431; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_432; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_433; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_434; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_435; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_436; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_437; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_438; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_439; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_440; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_441; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_442; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_443; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_444; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_445; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_446; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_447; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_448; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_449; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_450; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_451; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_452; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_453; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_454; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_455; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_456; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_457; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_458; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_459; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_460; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_461; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_462; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_463; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_464; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_465; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_466; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_467; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_468; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_469; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_470; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_471; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_472; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_473; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_474; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_475; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_476; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_477; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_478; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_479; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_480; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_481; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_482; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_483; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_484; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_485; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_486; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_487; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_488; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_489; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_490; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_491; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_492; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_493; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_494; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_495; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_496; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_497; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_498; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_499; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_500; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_501; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_502; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_503; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_504; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_505; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_506; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_507; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_508; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_509; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_510; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_511; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 129:23]
  wire [3:0] pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_key_in; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_key_out; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_sum_in; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_sum_out; // @[hash.scala 129:23]
  wire  pipe4_clock; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_160; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_161; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_162; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_163; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_164; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_165; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_166; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_167; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_168; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_169; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_170; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_171; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_172; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_173; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_174; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_175; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_176; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_177; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_178; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_179; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_180; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_181; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_182; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_183; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_184; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_185; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_186; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_187; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_188; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_189; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_190; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_191; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_192; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_193; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_194; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_195; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_196; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_197; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_198; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_199; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_200; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_201; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_202; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_203; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_204; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_205; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_206; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_207; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_208; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_209; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_210; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_211; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_212; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_213; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_214; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_215; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_216; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_217; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_218; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_219; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_220; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_221; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_222; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_223; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_224; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_225; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_226; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_227; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_228; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_229; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_230; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_231; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_232; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_233; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_234; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_235; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_236; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_237; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_238; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_239; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_240; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_241; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_242; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_243; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_244; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_245; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_246; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_247; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_248; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_249; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_250; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_251; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_252; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_253; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_254; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_255; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_256; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_257; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_258; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_259; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_260; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_261; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_262; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_263; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_264; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_265; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_266; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_267; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_268; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_269; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_270; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_271; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_272; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_273; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_274; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_275; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_276; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_277; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_278; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_279; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_280; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_281; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_282; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_283; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_284; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_285; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_286; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_287; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_288; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_289; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_290; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_291; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_292; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_293; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_294; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_295; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_296; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_297; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_298; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_299; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_300; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_301; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_302; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_303; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_304; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_305; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_306; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_307; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_308; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_309; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_310; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_311; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_312; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_313; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_314; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_315; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_316; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_317; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_318; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_319; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_320; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_321; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_322; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_323; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_324; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_325; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_326; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_327; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_328; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_329; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_330; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_331; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_332; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_333; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_334; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_335; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_336; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_337; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_338; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_339; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_340; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_341; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_342; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_343; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_344; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_345; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_346; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_347; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_348; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_349; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_350; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_351; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_352; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_353; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_354; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_355; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_356; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_357; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_358; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_359; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_360; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_361; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_362; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_363; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_364; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_365; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_366; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_367; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_368; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_369; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_370; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_371; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_372; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_373; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_374; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_375; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_376; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_377; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_378; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_379; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_380; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_381; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_382; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_383; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_384; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_385; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_386; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_387; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_388; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_389; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_390; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_391; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_392; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_393; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_394; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_395; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_396; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_397; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_398; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_399; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_400; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_401; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_402; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_403; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_404; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_405; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_406; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_407; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_408; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_409; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_410; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_411; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_412; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_413; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_414; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_415; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_416; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_417; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_418; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_419; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_420; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_421; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_422; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_423; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_424; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_425; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_426; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_427; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_428; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_429; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_430; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_431; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_432; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_433; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_434; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_435; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_436; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_437; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_438; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_439; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_440; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_441; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_442; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_443; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_444; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_445; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_446; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_447; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_448; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_449; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_450; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_451; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_452; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_453; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_454; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_455; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_456; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_457; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_458; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_459; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_460; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_461; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_462; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_463; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_464; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_465; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_466; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_467; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_468; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_469; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_470; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_471; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_472; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_473; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_474; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_475; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_476; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_477; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_478; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_479; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_480; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_481; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_482; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_483; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_484; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_485; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_486; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_487; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_488; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_489; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_490; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_491; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_492; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_493; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_494; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_495; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_496; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_497; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_498; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_499; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_500; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_501; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_502; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_503; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_504; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_505; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_506; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_507; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_508; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_509; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_510; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_511; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[hash.scala 130:23]
  wire [3:0] pipe4_io_pipe_phv_in_next_processor_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_160; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_161; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_162; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_163; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_164; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_165; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_166; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_167; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_168; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_169; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_170; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_171; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_172; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_173; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_174; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_175; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_176; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_177; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_178; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_179; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_180; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_181; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_182; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_183; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_184; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_185; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_186; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_187; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_188; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_189; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_190; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_191; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_192; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_193; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_194; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_195; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_196; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_197; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_198; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_199; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_200; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_201; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_202; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_203; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_204; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_205; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_206; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_207; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_208; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_209; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_210; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_211; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_212; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_213; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_214; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_215; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_216; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_217; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_218; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_219; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_220; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_221; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_222; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_223; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_224; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_225; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_226; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_227; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_228; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_229; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_230; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_231; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_232; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_233; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_234; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_235; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_236; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_237; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_238; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_239; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_240; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_241; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_242; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_243; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_244; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_245; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_246; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_247; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_248; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_249; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_250; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_251; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_252; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_253; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_254; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_255; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_256; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_257; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_258; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_259; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_260; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_261; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_262; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_263; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_264; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_265; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_266; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_267; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_268; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_269; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_270; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_271; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_272; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_273; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_274; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_275; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_276; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_277; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_278; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_279; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_280; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_281; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_282; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_283; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_284; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_285; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_286; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_287; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_288; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_289; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_290; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_291; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_292; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_293; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_294; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_295; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_296; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_297; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_298; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_299; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_300; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_301; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_302; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_303; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_304; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_305; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_306; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_307; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_308; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_309; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_310; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_311; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_312; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_313; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_314; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_315; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_316; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_317; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_318; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_319; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_320; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_321; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_322; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_323; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_324; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_325; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_326; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_327; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_328; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_329; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_330; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_331; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_332; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_333; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_334; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_335; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_336; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_337; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_338; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_339; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_340; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_341; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_342; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_343; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_344; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_345; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_346; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_347; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_348; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_349; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_350; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_351; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_352; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_353; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_354; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_355; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_356; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_357; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_358; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_359; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_360; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_361; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_362; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_363; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_364; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_365; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_366; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_367; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_368; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_369; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_370; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_371; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_372; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_373; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_374; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_375; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_376; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_377; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_378; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_379; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_380; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_381; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_382; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_383; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_384; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_385; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_386; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_387; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_388; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_389; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_390; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_391; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_392; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_393; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_394; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_395; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_396; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_397; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_398; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_399; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_400; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_401; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_402; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_403; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_404; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_405; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_406; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_407; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_408; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_409; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_410; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_411; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_412; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_413; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_414; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_415; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_416; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_417; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_418; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_419; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_420; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_421; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_422; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_423; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_424; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_425; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_426; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_427; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_428; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_429; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_430; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_431; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_432; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_433; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_434; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_435; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_436; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_437; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_438; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_439; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_440; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_441; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_442; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_443; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_444; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_445; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_446; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_447; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_448; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_449; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_450; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_451; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_452; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_453; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_454; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_455; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_456; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_457; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_458; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_459; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_460; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_461; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_462; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_463; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_464; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_465; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_466; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_467; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_468; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_469; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_470; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_471; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_472; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_473; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_474; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_475; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_476; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_477; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_478; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_479; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_480; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_481; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_482; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_483; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_484; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_485; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_486; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_487; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_488; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_489; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_490; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_491; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_492; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_493; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_494; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_495; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_496; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_497; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_498; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_499; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_500; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_501; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_502; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_503; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_504; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_505; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_506; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_507; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_508; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_509; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_510; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_511; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 130:23]
  wire [3:0] pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_key_in; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_key_out; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_sum_in; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_sum_out; // @[hash.scala 130:23]
  wire  pipe5_clock; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_96; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_97; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_98; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_99; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_100; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_101; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_102; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_103; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_104; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_105; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_106; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_107; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_108; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_109; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_110; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_111; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_112; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_113; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_114; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_115; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_116; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_117; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_118; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_119; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_120; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_121; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_122; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_123; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_124; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_125; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_126; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_127; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_128; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_129; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_130; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_131; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_132; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_133; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_134; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_135; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_136; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_137; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_138; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_139; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_140; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_141; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_142; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_143; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_144; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_145; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_146; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_147; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_148; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_149; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_150; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_151; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_152; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_153; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_154; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_155; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_156; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_157; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_158; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_159; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_160; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_161; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_162; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_163; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_164; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_165; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_166; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_167; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_168; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_169; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_170; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_171; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_172; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_173; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_174; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_175; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_176; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_177; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_178; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_179; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_180; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_181; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_182; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_183; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_184; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_185; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_186; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_187; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_188; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_189; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_190; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_191; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_192; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_193; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_194; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_195; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_196; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_197; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_198; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_199; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_200; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_201; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_202; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_203; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_204; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_205; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_206; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_207; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_208; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_209; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_210; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_211; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_212; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_213; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_214; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_215; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_216; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_217; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_218; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_219; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_220; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_221; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_222; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_223; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_224; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_225; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_226; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_227; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_228; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_229; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_230; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_231; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_232; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_233; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_234; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_235; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_236; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_237; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_238; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_239; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_240; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_241; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_242; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_243; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_244; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_245; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_246; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_247; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_248; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_249; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_250; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_251; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_252; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_253; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_254; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_255; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_256; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_257; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_258; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_259; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_260; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_261; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_262; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_263; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_264; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_265; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_266; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_267; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_268; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_269; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_270; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_271; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_272; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_273; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_274; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_275; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_276; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_277; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_278; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_279; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_280; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_281; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_282; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_283; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_284; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_285; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_286; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_287; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_288; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_289; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_290; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_291; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_292; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_293; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_294; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_295; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_296; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_297; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_298; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_299; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_300; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_301; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_302; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_303; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_304; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_305; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_306; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_307; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_308; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_309; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_310; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_311; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_312; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_313; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_314; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_315; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_316; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_317; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_318; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_319; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_320; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_321; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_322; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_323; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_324; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_325; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_326; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_327; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_328; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_329; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_330; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_331; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_332; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_333; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_334; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_335; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_336; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_337; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_338; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_339; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_340; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_341; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_342; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_343; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_344; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_345; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_346; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_347; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_348; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_349; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_350; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_351; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_352; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_353; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_354; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_355; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_356; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_357; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_358; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_359; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_360; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_361; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_362; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_363; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_364; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_365; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_366; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_367; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_368; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_369; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_370; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_371; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_372; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_373; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_374; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_375; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_376; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_377; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_378; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_379; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_380; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_381; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_382; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_383; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_384; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_385; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_386; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_387; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_388; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_389; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_390; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_391; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_392; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_393; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_394; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_395; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_396; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_397; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_398; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_399; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_400; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_401; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_402; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_403; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_404; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_405; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_406; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_407; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_408; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_409; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_410; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_411; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_412; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_413; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_414; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_415; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_416; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_417; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_418; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_419; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_420; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_421; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_422; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_423; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_424; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_425; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_426; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_427; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_428; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_429; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_430; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_431; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_432; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_433; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_434; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_435; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_436; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_437; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_438; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_439; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_440; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_441; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_442; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_443; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_444; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_445; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_446; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_447; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_448; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_449; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_450; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_451; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_452; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_453; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_454; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_455; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_456; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_457; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_458; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_459; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_460; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_461; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_462; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_463; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_464; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_465; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_466; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_467; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_468; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_469; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_470; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_471; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_472; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_473; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_474; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_475; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_476; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_477; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_478; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_479; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_480; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_481; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_482; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_483; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_484; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_485; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_486; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_487; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_488; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_489; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_490; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_491; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_492; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_493; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_494; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_495; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_496; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_497; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_498; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_499; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_500; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_501; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_502; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_503; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_504; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_505; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_506; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_507; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_508; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_509; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_510; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_511; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_pipe_phv_in_next_processor_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_96; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_97; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_98; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_99; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_100; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_101; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_102; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_103; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_104; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_105; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_106; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_107; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_108; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_109; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_110; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_111; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_112; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_113; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_114; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_115; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_116; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_117; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_118; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_119; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_120; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_121; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_122; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_123; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_124; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_125; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_126; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_127; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_128; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_129; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_130; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_131; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_132; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_133; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_134; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_135; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_136; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_137; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_138; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_139; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_140; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_141; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_142; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_143; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_144; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_145; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_146; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_147; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_148; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_149; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_150; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_151; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_152; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_153; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_154; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_155; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_156; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_157; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_158; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_159; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_160; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_161; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_162; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_163; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_164; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_165; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_166; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_167; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_168; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_169; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_170; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_171; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_172; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_173; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_174; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_175; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_176; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_177; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_178; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_179; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_180; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_181; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_182; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_183; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_184; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_185; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_186; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_187; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_188; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_189; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_190; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_191; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_192; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_193; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_194; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_195; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_196; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_197; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_198; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_199; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_200; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_201; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_202; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_203; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_204; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_205; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_206; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_207; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_208; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_209; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_210; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_211; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_212; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_213; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_214; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_215; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_216; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_217; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_218; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_219; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_220; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_221; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_222; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_223; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_224; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_225; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_226; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_227; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_228; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_229; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_230; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_231; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_232; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_233; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_234; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_235; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_236; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_237; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_238; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_239; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_240; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_241; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_242; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_243; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_244; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_245; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_246; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_247; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_248; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_249; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_250; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_251; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_252; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_253; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_254; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_255; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_256; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_257; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_258; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_259; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_260; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_261; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_262; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_263; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_264; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_265; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_266; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_267; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_268; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_269; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_270; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_271; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_272; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_273; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_274; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_275; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_276; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_277; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_278; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_279; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_280; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_281; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_282; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_283; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_284; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_285; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_286; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_287; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_288; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_289; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_290; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_291; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_292; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_293; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_294; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_295; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_296; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_297; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_298; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_299; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_300; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_301; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_302; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_303; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_304; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_305; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_306; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_307; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_308; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_309; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_310; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_311; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_312; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_313; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_314; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_315; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_316; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_317; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_318; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_319; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_320; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_321; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_322; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_323; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_324; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_325; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_326; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_327; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_328; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_329; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_330; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_331; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_332; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_333; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_334; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_335; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_336; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_337; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_338; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_339; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_340; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_341; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_342; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_343; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_344; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_345; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_346; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_347; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_348; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_349; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_350; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_351; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_352; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_353; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_354; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_355; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_356; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_357; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_358; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_359; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_360; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_361; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_362; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_363; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_364; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_365; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_366; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_367; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_368; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_369; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_370; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_371; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_372; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_373; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_374; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_375; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_376; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_377; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_378; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_379; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_380; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_381; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_382; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_383; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_384; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_385; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_386; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_387; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_388; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_389; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_390; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_391; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_392; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_393; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_394; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_395; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_396; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_397; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_398; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_399; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_400; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_401; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_402; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_403; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_404; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_405; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_406; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_407; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_408; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_409; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_410; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_411; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_412; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_413; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_414; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_415; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_416; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_417; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_418; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_419; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_420; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_421; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_422; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_423; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_424; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_425; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_426; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_427; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_428; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_429; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_430; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_431; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_432; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_433; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_434; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_435; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_436; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_437; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_438; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_439; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_440; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_441; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_442; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_443; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_444; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_445; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_446; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_447; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_448; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_449; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_450; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_451; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_452; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_453; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_454; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_455; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_456; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_457; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_458; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_459; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_460; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_461; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_462; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_463; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_464; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_465; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_466; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_467; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_468; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_469; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_470; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_471; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_472; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_473; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_474; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_475; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_476; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_477; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_478; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_479; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_480; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_481; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_482; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_483; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_484; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_485; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_486; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_487; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_488; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_489; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_490; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_491; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_492; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_493; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_494; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_495; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_496; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_497; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_498; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_499; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_500; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_501; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_502; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_503; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_504; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_505; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_506; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_507; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_508; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_509; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_510; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_511; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_hash_depth_0; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_hash_depth_1; // @[hash.scala 131:23]
  wire [191:0] pipe5_io_key_in; // @[hash.scala 131:23]
  wire [191:0] pipe5_io_key_out; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_sum_in; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_sum_out; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_val_out; // @[hash.scala 131:23]
  wire  pipe6_clock; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_96; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_97; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_98; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_99; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_100; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_101; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_102; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_103; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_104; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_105; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_106; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_107; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_108; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_109; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_110; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_111; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_112; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_113; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_114; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_115; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_116; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_117; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_118; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_119; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_120; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_121; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_122; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_123; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_124; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_125; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_126; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_127; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_128; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_129; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_130; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_131; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_132; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_133; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_134; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_135; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_136; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_137; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_138; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_139; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_140; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_141; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_142; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_143; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_144; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_145; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_146; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_147; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_148; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_149; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_150; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_151; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_152; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_153; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_154; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_155; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_156; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_157; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_158; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_159; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_160; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_161; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_162; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_163; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_164; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_165; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_166; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_167; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_168; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_169; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_170; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_171; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_172; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_173; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_174; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_175; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_176; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_177; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_178; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_179; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_180; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_181; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_182; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_183; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_184; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_185; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_186; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_187; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_188; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_189; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_190; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_191; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_192; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_193; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_194; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_195; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_196; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_197; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_198; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_199; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_200; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_201; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_202; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_203; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_204; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_205; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_206; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_207; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_208; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_209; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_210; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_211; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_212; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_213; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_214; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_215; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_216; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_217; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_218; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_219; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_220; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_221; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_222; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_223; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_224; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_225; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_226; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_227; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_228; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_229; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_230; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_231; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_232; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_233; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_234; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_235; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_236; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_237; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_238; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_239; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_240; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_241; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_242; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_243; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_244; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_245; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_246; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_247; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_248; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_249; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_250; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_251; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_252; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_253; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_254; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_255; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_256; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_257; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_258; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_259; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_260; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_261; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_262; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_263; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_264; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_265; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_266; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_267; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_268; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_269; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_270; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_271; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_272; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_273; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_274; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_275; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_276; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_277; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_278; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_279; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_280; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_281; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_282; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_283; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_284; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_285; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_286; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_287; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_288; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_289; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_290; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_291; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_292; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_293; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_294; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_295; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_296; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_297; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_298; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_299; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_300; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_301; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_302; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_303; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_304; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_305; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_306; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_307; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_308; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_309; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_310; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_311; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_312; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_313; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_314; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_315; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_316; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_317; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_318; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_319; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_320; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_321; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_322; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_323; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_324; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_325; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_326; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_327; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_328; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_329; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_330; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_331; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_332; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_333; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_334; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_335; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_336; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_337; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_338; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_339; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_340; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_341; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_342; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_343; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_344; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_345; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_346; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_347; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_348; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_349; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_350; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_351; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_352; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_353; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_354; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_355; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_356; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_357; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_358; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_359; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_360; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_361; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_362; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_363; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_364; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_365; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_366; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_367; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_368; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_369; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_370; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_371; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_372; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_373; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_374; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_375; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_376; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_377; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_378; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_379; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_380; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_381; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_382; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_383; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_384; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_385; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_386; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_387; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_388; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_389; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_390; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_391; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_392; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_393; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_394; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_395; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_396; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_397; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_398; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_399; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_400; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_401; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_402; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_403; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_404; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_405; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_406; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_407; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_408; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_409; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_410; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_411; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_412; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_413; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_414; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_415; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_416; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_417; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_418; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_419; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_420; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_421; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_422; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_423; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_424; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_425; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_426; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_427; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_428; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_429; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_430; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_431; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_432; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_433; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_434; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_435; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_436; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_437; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_438; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_439; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_440; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_441; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_442; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_443; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_444; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_445; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_446; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_447; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_448; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_449; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_450; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_451; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_452; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_453; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_454; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_455; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_456; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_457; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_458; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_459; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_460; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_461; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_462; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_463; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_464; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_465; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_466; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_467; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_468; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_469; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_470; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_471; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_472; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_473; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_474; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_475; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_476; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_477; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_478; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_479; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_480; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_481; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_482; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_483; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_484; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_485; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_486; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_487; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_488; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_489; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_490; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_491; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_492; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_493; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_494; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_495; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_496; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_497; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_498; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_499; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_500; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_501; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_502; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_503; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_504; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_505; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_506; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_507; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_508; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_509; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_510; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_511; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_pipe_phv_in_next_processor_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_96; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_97; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_98; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_99; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_100; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_101; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_102; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_103; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_104; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_105; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_106; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_107; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_108; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_109; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_110; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_111; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_112; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_113; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_114; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_115; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_116; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_117; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_118; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_119; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_120; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_121; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_122; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_123; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_124; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_125; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_126; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_127; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_128; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_129; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_130; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_131; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_132; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_133; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_134; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_135; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_136; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_137; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_138; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_139; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_140; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_141; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_142; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_143; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_144; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_145; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_146; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_147; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_148; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_149; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_150; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_151; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_152; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_153; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_154; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_155; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_156; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_157; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_158; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_159; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_160; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_161; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_162; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_163; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_164; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_165; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_166; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_167; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_168; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_169; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_170; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_171; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_172; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_173; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_174; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_175; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_176; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_177; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_178; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_179; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_180; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_181; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_182; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_183; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_184; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_185; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_186; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_187; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_188; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_189; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_190; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_191; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_192; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_193; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_194; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_195; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_196; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_197; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_198; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_199; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_200; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_201; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_202; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_203; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_204; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_205; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_206; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_207; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_208; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_209; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_210; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_211; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_212; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_213; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_214; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_215; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_216; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_217; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_218; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_219; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_220; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_221; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_222; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_223; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_224; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_225; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_226; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_227; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_228; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_229; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_230; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_231; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_232; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_233; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_234; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_235; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_236; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_237; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_238; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_239; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_240; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_241; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_242; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_243; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_244; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_245; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_246; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_247; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_248; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_249; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_250; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_251; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_252; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_253; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_254; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_255; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_256; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_257; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_258; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_259; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_260; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_261; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_262; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_263; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_264; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_265; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_266; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_267; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_268; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_269; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_270; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_271; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_272; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_273; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_274; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_275; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_276; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_277; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_278; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_279; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_280; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_281; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_282; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_283; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_284; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_285; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_286; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_287; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_288; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_289; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_290; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_291; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_292; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_293; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_294; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_295; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_296; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_297; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_298; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_299; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_300; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_301; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_302; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_303; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_304; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_305; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_306; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_307; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_308; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_309; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_310; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_311; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_312; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_313; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_314; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_315; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_316; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_317; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_318; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_319; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_320; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_321; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_322; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_323; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_324; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_325; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_326; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_327; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_328; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_329; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_330; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_331; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_332; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_333; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_334; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_335; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_336; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_337; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_338; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_339; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_340; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_341; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_342; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_343; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_344; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_345; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_346; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_347; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_348; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_349; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_350; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_351; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_352; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_353; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_354; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_355; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_356; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_357; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_358; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_359; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_360; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_361; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_362; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_363; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_364; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_365; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_366; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_367; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_368; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_369; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_370; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_371; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_372; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_373; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_374; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_375; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_376; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_377; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_378; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_379; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_380; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_381; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_382; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_383; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_384; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_385; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_386; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_387; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_388; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_389; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_390; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_391; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_392; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_393; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_394; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_395; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_396; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_397; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_398; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_399; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_400; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_401; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_402; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_403; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_404; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_405; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_406; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_407; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_408; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_409; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_410; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_411; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_412; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_413; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_414; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_415; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_416; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_417; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_418; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_419; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_420; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_421; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_422; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_423; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_424; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_425; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_426; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_427; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_428; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_429; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_430; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_431; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_432; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_433; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_434; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_435; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_436; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_437; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_438; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_439; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_440; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_441; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_442; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_443; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_444; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_445; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_446; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_447; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_448; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_449; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_450; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_451; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_452; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_453; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_454; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_455; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_456; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_457; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_458; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_459; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_460; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_461; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_462; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_463; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_464; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_465; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_466; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_467; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_468; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_469; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_470; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_471; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_472; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_473; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_474; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_475; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_476; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_477; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_478; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_479; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_480; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_481; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_482; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_483; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_484; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_485; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_486; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_487; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_488; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_489; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_490; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_491; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_492; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_493; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_494; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_495; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_496; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_497; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_498; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_499; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_500; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_501; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_502; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_503; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_504; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_505; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_506; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_507; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_508; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_509; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_510; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_511; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_hash_depth_0; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_hash_depth_1; // @[hash.scala 132:23]
  wire [191:0] pipe6_io_key_in; // @[hash.scala 132:23]
  wire [191:0] pipe6_io_key_out; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_sum_in; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_sum_out; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_val_in; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_val_out; // @[hash.scala 132:23]
  wire  pipe7_clock; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_0; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_1; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_2; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_3; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_4; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_5; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_6; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_7; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_8; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_9; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_10; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_11; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_12; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_13; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_14; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_16; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_17; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_18; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_19; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_20; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_21; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_22; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_23; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_24; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_25; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_26; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_27; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_28; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_29; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_30; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_31; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_32; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_33; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_34; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_35; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_36; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_37; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_38; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_39; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_40; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_41; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_42; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_43; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_44; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_45; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_46; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_47; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_48; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_49; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_50; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_51; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_52; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_53; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_54; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_55; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_56; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_57; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_58; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_59; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_60; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_61; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_62; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_63; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_64; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_65; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_66; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_67; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_68; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_69; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_70; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_71; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_72; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_73; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_74; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_75; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_76; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_77; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_78; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_79; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_80; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_81; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_82; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_83; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_84; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_85; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_86; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_87; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_88; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_89; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_90; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_91; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_92; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_93; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_94; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_95; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_96; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_97; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_98; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_99; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_100; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_101; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_102; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_103; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_104; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_105; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_106; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_107; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_108; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_109; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_110; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_111; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_112; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_113; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_114; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_115; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_116; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_117; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_118; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_119; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_120; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_121; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_122; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_123; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_124; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_125; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_126; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_127; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_128; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_129; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_130; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_131; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_132; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_133; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_134; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_135; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_136; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_137; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_138; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_139; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_140; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_141; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_142; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_143; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_144; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_145; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_146; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_147; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_148; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_149; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_150; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_151; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_152; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_153; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_154; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_155; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_156; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_157; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_158; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_159; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_160; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_161; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_162; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_163; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_164; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_165; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_166; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_167; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_168; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_169; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_170; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_171; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_172; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_173; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_174; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_175; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_176; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_177; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_178; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_179; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_180; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_181; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_182; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_183; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_184; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_185; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_186; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_187; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_188; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_189; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_190; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_191; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_192; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_193; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_194; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_195; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_196; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_197; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_198; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_199; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_200; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_201; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_202; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_203; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_204; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_205; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_206; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_207; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_208; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_209; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_210; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_211; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_212; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_213; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_214; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_215; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_216; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_217; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_218; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_219; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_220; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_221; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_222; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_223; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_224; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_225; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_226; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_227; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_228; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_229; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_230; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_231; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_232; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_233; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_234; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_235; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_236; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_237; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_238; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_239; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_240; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_241; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_242; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_243; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_244; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_245; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_246; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_247; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_248; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_249; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_250; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_251; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_252; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_253; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_254; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_255; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_256; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_257; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_258; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_259; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_260; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_261; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_262; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_263; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_264; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_265; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_266; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_267; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_268; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_269; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_270; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_271; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_272; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_273; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_274; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_275; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_276; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_277; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_278; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_279; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_280; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_281; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_282; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_283; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_284; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_285; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_286; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_287; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_288; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_289; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_290; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_291; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_292; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_293; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_294; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_295; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_296; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_297; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_298; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_299; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_300; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_301; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_302; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_303; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_304; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_305; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_306; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_307; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_308; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_309; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_310; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_311; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_312; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_313; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_314; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_315; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_316; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_317; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_318; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_319; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_320; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_321; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_322; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_323; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_324; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_325; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_326; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_327; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_328; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_329; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_330; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_331; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_332; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_333; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_334; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_335; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_336; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_337; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_338; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_339; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_340; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_341; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_342; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_343; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_344; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_345; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_346; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_347; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_348; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_349; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_350; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_351; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_352; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_353; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_354; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_355; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_356; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_357; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_358; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_359; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_360; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_361; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_362; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_363; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_364; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_365; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_366; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_367; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_368; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_369; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_370; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_371; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_372; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_373; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_374; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_375; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_376; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_377; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_378; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_379; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_380; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_381; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_382; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_383; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_384; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_385; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_386; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_387; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_388; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_389; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_390; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_391; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_392; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_393; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_394; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_395; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_396; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_397; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_398; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_399; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_400; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_401; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_402; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_403; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_404; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_405; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_406; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_407; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_408; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_409; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_410; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_411; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_412; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_413; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_414; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_415; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_416; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_417; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_418; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_419; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_420; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_421; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_422; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_423; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_424; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_425; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_426; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_427; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_428; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_429; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_430; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_431; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_432; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_433; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_434; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_435; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_436; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_437; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_438; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_439; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_440; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_441; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_442; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_443; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_444; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_445; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_446; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_447; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_448; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_449; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_450; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_451; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_452; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_453; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_454; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_455; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_456; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_457; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_458; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_459; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_460; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_461; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_462; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_463; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_464; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_465; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_466; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_467; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_468; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_469; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_470; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_471; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_472; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_473; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_474; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_475; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_476; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_477; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_478; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_479; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_480; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_481; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_482; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_483; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_484; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_485; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_486; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_487; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_488; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_489; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_490; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_491; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_492; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_493; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_494; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_495; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_496; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_497; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_498; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_499; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_500; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_501; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_502; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_503; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_504; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_505; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_506; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_507; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_508; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_509; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_510; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_511; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_0; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_1; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_2; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_3; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_4; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_5; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_6; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_7; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_8; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_9; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_10; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_11; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_12; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_13; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_14; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_parse_current_state; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_parse_current_offset; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_parse_transition_field; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_pipe_phv_in_next_processor_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_in_next_config_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_in_is_valid_processor; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_0; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_1; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_2; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_3; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_4; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_5; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_6; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_7; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_8; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_9; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_10; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_11; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_12; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_13; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_14; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_16; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_17; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_18; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_19; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_20; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_21; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_22; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_23; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_24; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_25; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_26; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_27; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_28; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_29; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_30; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_31; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_32; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_33; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_34; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_35; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_36; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_37; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_38; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_39; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_40; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_41; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_42; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_43; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_44; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_45; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_46; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_47; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_48; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_49; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_50; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_51; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_52; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_53; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_54; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_55; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_56; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_57; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_58; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_59; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_60; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_61; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_62; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_63; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_64; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_65; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_66; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_67; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_68; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_69; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_70; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_71; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_72; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_73; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_74; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_75; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_76; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_77; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_78; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_79; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_80; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_81; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_82; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_83; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_84; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_85; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_86; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_87; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_88; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_89; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_90; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_91; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_92; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_93; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_94; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_95; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_96; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_97; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_98; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_99; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_100; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_101; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_102; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_103; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_104; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_105; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_106; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_107; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_108; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_109; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_110; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_111; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_112; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_113; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_114; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_115; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_116; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_117; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_118; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_119; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_120; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_121; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_122; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_123; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_124; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_125; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_126; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_127; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_128; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_129; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_130; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_131; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_132; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_133; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_134; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_135; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_136; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_137; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_138; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_139; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_140; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_141; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_142; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_143; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_144; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_145; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_146; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_147; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_148; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_149; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_150; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_151; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_152; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_153; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_154; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_155; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_156; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_157; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_158; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_159; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_160; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_161; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_162; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_163; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_164; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_165; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_166; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_167; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_168; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_169; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_170; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_171; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_172; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_173; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_174; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_175; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_176; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_177; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_178; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_179; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_180; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_181; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_182; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_183; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_184; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_185; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_186; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_187; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_188; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_189; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_190; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_191; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_192; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_193; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_194; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_195; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_196; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_197; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_198; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_199; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_200; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_201; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_202; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_203; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_204; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_205; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_206; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_207; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_208; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_209; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_210; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_211; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_212; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_213; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_214; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_215; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_216; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_217; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_218; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_219; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_220; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_221; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_222; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_223; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_224; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_225; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_226; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_227; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_228; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_229; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_230; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_231; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_232; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_233; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_234; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_235; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_236; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_237; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_238; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_239; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_240; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_241; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_242; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_243; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_244; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_245; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_246; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_247; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_248; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_249; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_250; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_251; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_252; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_253; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_254; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_255; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_256; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_257; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_258; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_259; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_260; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_261; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_262; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_263; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_264; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_265; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_266; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_267; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_268; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_269; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_270; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_271; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_272; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_273; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_274; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_275; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_276; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_277; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_278; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_279; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_280; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_281; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_282; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_283; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_284; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_285; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_286; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_287; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_288; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_289; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_290; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_291; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_292; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_293; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_294; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_295; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_296; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_297; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_298; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_299; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_300; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_301; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_302; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_303; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_304; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_305; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_306; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_307; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_308; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_309; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_310; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_311; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_312; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_313; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_314; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_315; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_316; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_317; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_318; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_319; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_320; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_321; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_322; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_323; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_324; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_325; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_326; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_327; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_328; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_329; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_330; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_331; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_332; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_333; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_334; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_335; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_336; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_337; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_338; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_339; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_340; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_341; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_342; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_343; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_344; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_345; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_346; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_347; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_348; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_349; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_350; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_351; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_352; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_353; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_354; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_355; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_356; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_357; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_358; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_359; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_360; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_361; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_362; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_363; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_364; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_365; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_366; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_367; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_368; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_369; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_370; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_371; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_372; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_373; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_374; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_375; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_376; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_377; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_378; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_379; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_380; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_381; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_382; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_383; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_384; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_385; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_386; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_387; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_388; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_389; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_390; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_391; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_392; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_393; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_394; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_395; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_396; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_397; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_398; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_399; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_400; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_401; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_402; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_403; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_404; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_405; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_406; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_407; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_408; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_409; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_410; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_411; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_412; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_413; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_414; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_415; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_416; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_417; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_418; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_419; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_420; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_421; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_422; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_423; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_424; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_425; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_426; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_427; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_428; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_429; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_430; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_431; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_432; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_433; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_434; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_435; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_436; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_437; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_438; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_439; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_440; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_441; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_442; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_443; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_444; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_445; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_446; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_447; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_448; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_449; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_450; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_451; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_452; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_453; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_454; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_455; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_456; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_457; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_458; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_459; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_460; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_461; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_462; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_463; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_464; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_465; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_466; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_467; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_468; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_469; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_470; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_471; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_472; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_473; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_474; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_475; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_476; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_477; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_478; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_479; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_480; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_481; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_482; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_483; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_484; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_485; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_486; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_487; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_488; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_489; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_490; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_491; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_492; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_493; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_494; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_495; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_496; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_497; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_498; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_499; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_500; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_501; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_502; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_503; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_504; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_505; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_506; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_507; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_508; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_509; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_510; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_511; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_0; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_1; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_2; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_3; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_4; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_5; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_6; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_7; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_8; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_9; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_10; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_11; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_12; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_13; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_14; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_parse_current_state; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_parse_current_offset; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_parse_transition_field; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_pipe_phv_out_next_processor_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_out_next_config_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_out_is_valid_processor; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_hash_depth_0; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_hash_depth_1; // @[hash.scala 133:23]
  wire [191:0] pipe7_io_key_in; // @[hash.scala 133:23]
  wire [191:0] pipe7_io_key_out; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_sum_in; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_sum_out; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_val_in; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_val_out; // @[hash.scala 133:23]
  wire  pipe8_clock; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_0; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_1; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_2; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_3; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_4; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_5; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_6; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_7; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_8; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_9; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_10; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_11; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_12; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_13; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_14; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_16; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_17; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_18; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_19; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_20; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_21; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_22; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_23; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_24; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_25; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_26; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_27; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_28; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_29; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_30; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_31; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_32; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_33; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_34; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_35; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_36; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_37; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_38; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_39; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_40; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_41; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_42; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_43; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_44; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_45; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_46; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_47; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_48; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_49; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_50; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_51; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_52; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_53; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_54; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_55; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_56; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_57; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_58; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_59; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_60; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_61; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_62; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_63; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_64; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_65; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_66; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_67; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_68; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_69; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_70; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_71; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_72; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_73; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_74; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_75; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_76; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_77; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_78; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_79; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_80; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_81; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_82; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_83; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_84; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_85; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_86; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_87; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_88; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_89; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_90; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_91; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_92; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_93; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_94; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_95; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_96; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_97; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_98; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_99; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_100; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_101; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_102; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_103; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_104; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_105; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_106; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_107; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_108; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_109; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_110; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_111; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_112; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_113; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_114; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_115; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_116; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_117; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_118; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_119; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_120; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_121; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_122; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_123; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_124; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_125; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_126; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_127; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_128; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_129; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_130; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_131; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_132; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_133; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_134; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_135; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_136; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_137; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_138; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_139; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_140; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_141; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_142; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_143; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_144; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_145; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_146; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_147; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_148; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_149; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_150; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_151; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_152; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_153; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_154; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_155; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_156; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_157; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_158; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_159; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_160; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_161; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_162; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_163; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_164; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_165; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_166; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_167; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_168; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_169; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_170; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_171; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_172; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_173; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_174; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_175; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_176; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_177; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_178; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_179; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_180; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_181; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_182; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_183; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_184; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_185; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_186; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_187; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_188; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_189; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_190; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_191; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_192; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_193; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_194; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_195; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_196; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_197; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_198; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_199; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_200; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_201; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_202; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_203; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_204; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_205; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_206; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_207; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_208; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_209; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_210; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_211; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_212; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_213; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_214; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_215; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_216; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_217; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_218; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_219; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_220; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_221; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_222; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_223; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_224; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_225; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_226; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_227; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_228; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_229; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_230; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_231; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_232; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_233; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_234; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_235; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_236; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_237; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_238; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_239; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_240; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_241; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_242; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_243; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_244; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_245; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_246; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_247; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_248; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_249; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_250; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_251; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_252; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_253; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_254; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_255; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_256; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_257; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_258; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_259; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_260; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_261; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_262; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_263; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_264; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_265; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_266; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_267; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_268; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_269; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_270; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_271; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_272; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_273; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_274; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_275; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_276; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_277; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_278; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_279; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_280; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_281; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_282; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_283; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_284; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_285; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_286; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_287; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_288; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_289; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_290; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_291; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_292; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_293; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_294; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_295; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_296; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_297; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_298; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_299; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_300; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_301; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_302; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_303; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_304; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_305; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_306; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_307; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_308; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_309; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_310; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_311; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_312; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_313; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_314; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_315; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_316; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_317; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_318; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_319; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_320; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_321; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_322; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_323; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_324; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_325; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_326; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_327; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_328; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_329; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_330; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_331; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_332; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_333; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_334; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_335; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_336; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_337; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_338; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_339; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_340; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_341; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_342; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_343; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_344; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_345; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_346; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_347; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_348; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_349; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_350; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_351; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_352; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_353; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_354; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_355; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_356; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_357; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_358; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_359; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_360; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_361; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_362; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_363; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_364; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_365; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_366; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_367; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_368; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_369; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_370; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_371; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_372; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_373; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_374; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_375; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_376; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_377; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_378; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_379; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_380; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_381; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_382; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_383; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_384; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_385; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_386; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_387; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_388; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_389; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_390; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_391; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_392; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_393; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_394; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_395; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_396; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_397; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_398; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_399; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_400; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_401; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_402; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_403; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_404; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_405; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_406; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_407; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_408; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_409; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_410; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_411; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_412; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_413; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_414; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_415; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_416; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_417; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_418; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_419; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_420; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_421; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_422; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_423; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_424; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_425; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_426; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_427; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_428; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_429; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_430; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_431; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_432; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_433; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_434; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_435; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_436; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_437; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_438; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_439; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_440; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_441; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_442; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_443; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_444; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_445; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_446; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_447; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_448; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_449; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_450; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_451; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_452; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_453; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_454; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_455; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_456; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_457; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_458; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_459; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_460; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_461; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_462; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_463; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_464; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_465; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_466; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_467; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_468; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_469; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_470; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_471; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_472; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_473; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_474; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_475; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_476; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_477; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_478; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_479; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_480; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_481; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_482; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_483; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_484; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_485; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_486; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_487; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_488; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_489; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_490; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_491; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_492; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_493; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_494; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_495; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_496; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_497; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_498; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_499; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_500; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_501; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_502; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_503; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_504; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_505; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_506; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_507; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_508; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_509; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_510; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_511; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_0; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_1; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_2; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_3; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_4; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_5; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_6; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_7; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_8; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_9; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_10; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_11; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_12; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_13; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_14; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_parse_current_state; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_parse_current_offset; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_parse_transition_field; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_pipe_phv_in_next_processor_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_in_next_config_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_in_is_valid_processor; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_0; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_1; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_2; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_3; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_4; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_5; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_6; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_7; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_8; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_9; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_10; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_11; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_12; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_13; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_14; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_16; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_17; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_18; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_19; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_20; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_21; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_22; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_23; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_24; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_25; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_26; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_27; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_28; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_29; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_30; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_31; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_32; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_33; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_34; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_35; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_36; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_37; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_38; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_39; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_40; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_41; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_42; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_43; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_44; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_45; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_46; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_47; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_48; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_49; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_50; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_51; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_52; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_53; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_54; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_55; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_56; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_57; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_58; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_59; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_60; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_61; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_62; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_63; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_64; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_65; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_66; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_67; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_68; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_69; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_70; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_71; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_72; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_73; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_74; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_75; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_76; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_77; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_78; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_79; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_80; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_81; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_82; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_83; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_84; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_85; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_86; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_87; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_88; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_89; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_90; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_91; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_92; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_93; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_94; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_95; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_96; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_97; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_98; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_99; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_100; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_101; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_102; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_103; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_104; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_105; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_106; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_107; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_108; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_109; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_110; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_111; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_112; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_113; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_114; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_115; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_116; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_117; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_118; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_119; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_120; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_121; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_122; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_123; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_124; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_125; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_126; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_127; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_128; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_129; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_130; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_131; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_132; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_133; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_134; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_135; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_136; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_137; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_138; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_139; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_140; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_141; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_142; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_143; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_144; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_145; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_146; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_147; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_148; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_149; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_150; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_151; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_152; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_153; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_154; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_155; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_156; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_157; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_158; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_159; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_160; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_161; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_162; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_163; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_164; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_165; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_166; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_167; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_168; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_169; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_170; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_171; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_172; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_173; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_174; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_175; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_176; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_177; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_178; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_179; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_180; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_181; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_182; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_183; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_184; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_185; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_186; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_187; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_188; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_189; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_190; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_191; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_192; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_193; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_194; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_195; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_196; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_197; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_198; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_199; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_200; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_201; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_202; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_203; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_204; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_205; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_206; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_207; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_208; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_209; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_210; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_211; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_212; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_213; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_214; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_215; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_216; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_217; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_218; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_219; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_220; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_221; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_222; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_223; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_224; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_225; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_226; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_227; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_228; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_229; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_230; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_231; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_232; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_233; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_234; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_235; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_236; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_237; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_238; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_239; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_240; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_241; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_242; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_243; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_244; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_245; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_246; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_247; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_248; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_249; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_250; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_251; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_252; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_253; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_254; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_255; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_256; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_257; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_258; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_259; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_260; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_261; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_262; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_263; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_264; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_265; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_266; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_267; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_268; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_269; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_270; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_271; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_272; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_273; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_274; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_275; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_276; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_277; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_278; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_279; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_280; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_281; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_282; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_283; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_284; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_285; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_286; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_287; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_288; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_289; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_290; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_291; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_292; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_293; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_294; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_295; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_296; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_297; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_298; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_299; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_300; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_301; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_302; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_303; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_304; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_305; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_306; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_307; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_308; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_309; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_310; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_311; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_312; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_313; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_314; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_315; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_316; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_317; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_318; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_319; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_320; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_321; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_322; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_323; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_324; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_325; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_326; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_327; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_328; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_329; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_330; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_331; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_332; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_333; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_334; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_335; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_336; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_337; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_338; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_339; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_340; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_341; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_342; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_343; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_344; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_345; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_346; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_347; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_348; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_349; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_350; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_351; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_352; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_353; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_354; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_355; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_356; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_357; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_358; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_359; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_360; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_361; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_362; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_363; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_364; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_365; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_366; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_367; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_368; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_369; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_370; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_371; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_372; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_373; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_374; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_375; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_376; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_377; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_378; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_379; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_380; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_381; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_382; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_383; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_384; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_385; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_386; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_387; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_388; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_389; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_390; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_391; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_392; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_393; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_394; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_395; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_396; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_397; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_398; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_399; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_400; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_401; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_402; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_403; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_404; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_405; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_406; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_407; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_408; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_409; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_410; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_411; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_412; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_413; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_414; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_415; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_416; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_417; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_418; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_419; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_420; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_421; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_422; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_423; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_424; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_425; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_426; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_427; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_428; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_429; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_430; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_431; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_432; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_433; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_434; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_435; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_436; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_437; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_438; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_439; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_440; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_441; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_442; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_443; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_444; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_445; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_446; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_447; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_448; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_449; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_450; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_451; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_452; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_453; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_454; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_455; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_456; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_457; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_458; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_459; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_460; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_461; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_462; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_463; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_464; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_465; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_466; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_467; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_468; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_469; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_470; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_471; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_472; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_473; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_474; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_475; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_476; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_477; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_478; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_479; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_480; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_481; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_482; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_483; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_484; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_485; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_486; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_487; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_488; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_489; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_490; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_491; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_492; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_493; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_494; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_495; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_496; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_497; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_498; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_499; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_500; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_501; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_502; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_503; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_504; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_505; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_506; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_507; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_508; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_509; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_510; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_511; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_0; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_1; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_2; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_3; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_4; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_5; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_6; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_7; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_8; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_9; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_10; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_11; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_12; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_13; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_14; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_parse_current_state; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_parse_current_offset; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_parse_transition_field; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_pipe_phv_out_next_processor_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_out_next_config_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_out_is_valid_processor; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_hash_depth_0; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_hash_depth_1; // @[hash.scala 134:23]
  wire [191:0] pipe8_io_key_in; // @[hash.scala 134:23]
  wire [191:0] pipe8_io_key_out; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_sum_in; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_sum_out; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_val_in; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_val_out; // @[hash.scala 134:23]
  reg [3:0] hash_depth_0; // @[hash.scala 18:26]
  reg [3:0] hash_depth_1; // @[hash.scala 18:26]
  HashSumLevel pipe1 ( // @[hash.scala 127:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe1_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe1_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe1_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe1_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe1_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe1_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe1_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe1_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe1_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe1_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe1_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe1_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe1_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe1_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe1_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe1_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe1_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe1_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe1_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe1_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe1_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe1_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe1_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe1_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe1_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe1_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe1_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe1_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe1_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe1_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe1_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe1_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe1_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe1_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe1_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe1_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe1_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe1_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe1_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe1_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe1_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe1_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe1_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe1_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe1_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe1_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe1_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe1_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe1_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe1_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe1_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe1_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe1_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe1_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe1_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe1_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe1_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe1_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe1_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe1_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe1_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe1_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe1_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe1_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe1_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe1_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe1_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe1_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe1_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe1_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe1_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe1_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe1_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe1_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe1_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe1_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe1_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe1_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe1_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe1_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe1_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe1_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe1_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe1_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe1_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe1_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe1_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe1_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe1_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe1_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe1_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe1_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe1_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe1_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe1_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe1_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe1_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe1_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe1_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe1_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe1_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe1_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe1_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe1_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe1_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe1_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe1_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe1_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe1_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe1_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe1_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe1_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe1_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe1_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe1_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe1_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe1_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe1_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe1_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe1_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe1_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe1_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe1_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe1_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe1_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe1_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe1_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe1_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe1_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe1_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe1_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe1_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe1_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe1_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe1_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe1_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe1_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe1_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe1_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe1_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe1_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe1_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe1_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe1_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe1_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe1_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe1_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe1_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe1_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe1_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe1_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe1_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe1_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe1_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe1_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe1_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe1_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe1_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe1_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe1_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe1_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe1_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe1_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe1_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe1_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe1_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe1_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe1_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe1_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe1_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe1_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe1_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe1_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe1_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe1_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe1_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe1_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe1_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe1_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe1_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe1_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe1_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe1_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe1_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe1_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe1_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe1_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe1_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe1_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe1_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe1_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe1_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe1_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe1_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe1_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe1_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe1_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe1_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe1_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe1_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe1_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe1_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe1_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe1_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe1_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe1_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe1_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe1_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe1_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe1_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe1_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe1_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe1_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe1_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe1_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe1_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe1_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe1_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe1_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe1_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe1_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe1_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe1_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe1_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe1_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe1_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe1_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe1_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe1_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe1_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe1_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe1_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe1_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe1_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe1_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe1_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe1_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe1_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe1_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe1_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe1_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe1_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe1_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe1_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe1_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe1_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe1_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe1_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe1_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe1_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe1_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe1_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe1_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe1_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe1_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe1_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe1_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe1_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe1_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe1_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe1_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe1_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe1_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe1_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe1_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe1_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe1_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe1_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe1_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe1_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe1_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe1_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe1_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe1_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe1_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe1_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe1_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe1_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe1_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe1_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe1_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe1_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe1_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe1_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe1_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe1_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe1_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe1_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe1_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe1_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe1_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe1_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe1_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe1_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe1_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe1_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe1_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe1_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe1_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe1_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe1_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe1_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe1_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe1_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe1_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe1_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe1_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe1_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe1_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe1_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe1_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe1_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe1_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe1_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe1_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe1_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe1_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe1_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe1_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe1_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe1_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe1_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe1_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe1_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe1_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe1_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe1_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe1_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe1_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe1_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe1_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe1_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe1_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe1_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe1_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe1_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe1_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe1_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe1_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe1_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe1_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe1_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe1_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe1_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe1_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe1_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe1_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe1_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe1_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe1_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe1_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe1_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe1_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe1_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe1_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe1_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe1_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe1_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe1_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe1_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe1_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe1_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe1_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe1_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe1_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe1_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe1_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe1_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe1_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe1_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe1_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe1_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe1_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe1_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe1_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe1_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe1_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe1_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe1_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe1_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe1_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe1_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe1_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe1_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe1_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe1_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe1_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe1_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe1_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe1_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe1_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe1_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe1_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe1_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe1_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe1_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe1_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe1_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe1_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe1_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe1_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe1_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe1_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe1_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe1_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe1_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe1_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe1_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe1_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe1_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe1_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe1_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe1_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe1_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe1_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe1_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe1_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe1_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe1_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe1_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe1_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe1_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe1_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe1_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe1_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe1_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe1_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe1_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe1_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe1_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe1_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe1_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe1_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe1_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe1_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe1_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe1_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe1_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe1_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe1_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe1_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe1_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe1_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe1_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe1_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe1_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe1_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe1_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe1_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe1_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe1_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe1_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe1_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe1_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe1_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe1_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe1_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe1_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe1_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe1_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe1_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe1_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe1_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe1_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe1_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe1_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe1_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe1_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe1_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe1_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe1_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe1_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe1_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe1_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe1_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe1_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe1_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe1_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe1_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe1_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe1_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe1_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe1_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe1_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe1_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe1_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe1_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe1_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe1_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe1_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe1_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe1_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe1_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe1_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe1_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe1_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe1_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe1_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe1_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe1_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe1_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe1_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe1_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe1_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe1_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe1_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe1_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe1_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe1_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe1_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe1_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe1_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe1_io_key_in),
    .io_key_out(pipe1_io_key_out),
    .io_sum_in(pipe1_io_sum_in),
    .io_sum_out(pipe1_io_sum_out)
  );
  HashSumLevel_1 pipe2 ( // @[hash.scala 128:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe2_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe2_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe2_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe2_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe2_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe2_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe2_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe2_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe2_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe2_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe2_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe2_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe2_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe2_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe2_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe2_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe2_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe2_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe2_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe2_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe2_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe2_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe2_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe2_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe2_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe2_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe2_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe2_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe2_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe2_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe2_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe2_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe2_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe2_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe2_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe2_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe2_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe2_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe2_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe2_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe2_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe2_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe2_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe2_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe2_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe2_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe2_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe2_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe2_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe2_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe2_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe2_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe2_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe2_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe2_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe2_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe2_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe2_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe2_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe2_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe2_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe2_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe2_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe2_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe2_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe2_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe2_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe2_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe2_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe2_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe2_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe2_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe2_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe2_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe2_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe2_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe2_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe2_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe2_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe2_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe2_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe2_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe2_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe2_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe2_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe2_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe2_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe2_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe2_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe2_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe2_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe2_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe2_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe2_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe2_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe2_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe2_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe2_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe2_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe2_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe2_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe2_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe2_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe2_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe2_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe2_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe2_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe2_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe2_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe2_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe2_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe2_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe2_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe2_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe2_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe2_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe2_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe2_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe2_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe2_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe2_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe2_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe2_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe2_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe2_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe2_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe2_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe2_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe2_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe2_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe2_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe2_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe2_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe2_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe2_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe2_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe2_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe2_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe2_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe2_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe2_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe2_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe2_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe2_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe2_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe2_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe2_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe2_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe2_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe2_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe2_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe2_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe2_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe2_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe2_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe2_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe2_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe2_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe2_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe2_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe2_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe2_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe2_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe2_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe2_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe2_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe2_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe2_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe2_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe2_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe2_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe2_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe2_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe2_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe2_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe2_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe2_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe2_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe2_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe2_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe2_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe2_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe2_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe2_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe2_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe2_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe2_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe2_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe2_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe2_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe2_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe2_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe2_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe2_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe2_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe2_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe2_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe2_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe2_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe2_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe2_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe2_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe2_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe2_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe2_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe2_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe2_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe2_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe2_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe2_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe2_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe2_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe2_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe2_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe2_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe2_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe2_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe2_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe2_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe2_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe2_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe2_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe2_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe2_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe2_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe2_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe2_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe2_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe2_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe2_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe2_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe2_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe2_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe2_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe2_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe2_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe2_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe2_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe2_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe2_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe2_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe2_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe2_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe2_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe2_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe2_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe2_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe2_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe2_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe2_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe2_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe2_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe2_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe2_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe2_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe2_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe2_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe2_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe2_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe2_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe2_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe2_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe2_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe2_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe2_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe2_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe2_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe2_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe2_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe2_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe2_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe2_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe2_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe2_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe2_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe2_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe2_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe2_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe2_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe2_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe2_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe2_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe2_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe2_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe2_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe2_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe2_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe2_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe2_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe2_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe2_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe2_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe2_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe2_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe2_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe2_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe2_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe2_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe2_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe2_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe2_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe2_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe2_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe2_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe2_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe2_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe2_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe2_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe2_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe2_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe2_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe2_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe2_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe2_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe2_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe2_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe2_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe2_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe2_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe2_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe2_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe2_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe2_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe2_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe2_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe2_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe2_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe2_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe2_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe2_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe2_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe2_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe2_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe2_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe2_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe2_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe2_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe2_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe2_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe2_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe2_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe2_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe2_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe2_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe2_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe2_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe2_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe2_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe2_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe2_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe2_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe2_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe2_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe2_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe2_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe2_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe2_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe2_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe2_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe2_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe2_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe2_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe2_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe2_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe2_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe2_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe2_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe2_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe2_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe2_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe2_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe2_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe2_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe2_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe2_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe2_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe2_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe2_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe2_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe2_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe2_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe2_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe2_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe2_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe2_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe2_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe2_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe2_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe2_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe2_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe2_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe2_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe2_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe2_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe2_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe2_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe2_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe2_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe2_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe2_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe2_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe2_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe2_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe2_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe2_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe2_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe2_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe2_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe2_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe2_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe2_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe2_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe2_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe2_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe2_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe2_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe2_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe2_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe2_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe2_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe2_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe2_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe2_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe2_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe2_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe2_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe2_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe2_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe2_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe2_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe2_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe2_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe2_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe2_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe2_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe2_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe2_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe2_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe2_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe2_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe2_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe2_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe2_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe2_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe2_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe2_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe2_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe2_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe2_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe2_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe2_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe2_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe2_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe2_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe2_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe2_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe2_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe2_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe2_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe2_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe2_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe2_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe2_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe2_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe2_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe2_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe2_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe2_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe2_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe2_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe2_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe2_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe2_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe2_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe2_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe2_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe2_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe2_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe2_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe2_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe2_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe2_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe2_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe2_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe2_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe2_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe2_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe2_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe2_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe2_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe2_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe2_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe2_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe2_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe2_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe2_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe2_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe2_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe2_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe2_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe2_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe2_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe2_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe2_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe2_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe2_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe2_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe2_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe2_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe2_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe2_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe2_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe2_io_key_in),
    .io_key_out(pipe2_io_key_out),
    .io_sum_in(pipe2_io_sum_in),
    .io_sum_out(pipe2_io_sum_out)
  );
  HashSumLevel_2 pipe3 ( // @[hash.scala 129:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe3_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe3_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe3_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe3_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe3_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe3_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe3_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe3_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe3_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe3_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe3_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe3_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe3_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe3_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe3_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe3_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe3_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe3_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe3_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe3_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe3_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe3_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe3_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe3_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe3_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe3_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe3_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe3_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe3_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe3_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe3_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe3_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe3_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe3_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe3_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe3_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe3_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe3_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe3_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe3_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe3_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe3_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe3_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe3_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe3_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe3_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe3_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe3_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe3_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe3_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe3_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe3_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe3_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe3_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe3_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe3_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe3_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe3_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe3_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe3_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe3_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe3_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe3_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe3_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe3_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe3_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe3_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe3_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe3_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe3_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe3_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe3_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe3_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe3_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe3_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe3_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe3_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe3_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe3_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe3_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe3_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe3_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe3_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe3_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe3_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe3_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe3_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe3_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe3_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe3_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe3_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe3_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe3_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe3_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe3_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe3_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe3_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe3_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe3_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe3_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe3_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe3_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe3_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe3_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe3_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe3_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe3_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe3_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe3_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe3_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe3_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe3_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe3_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe3_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe3_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe3_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe3_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe3_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe3_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe3_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe3_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe3_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe3_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe3_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe3_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe3_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe3_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe3_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe3_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe3_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe3_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe3_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe3_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe3_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe3_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe3_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe3_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe3_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe3_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe3_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe3_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe3_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe3_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe3_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe3_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe3_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe3_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe3_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe3_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe3_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe3_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe3_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe3_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe3_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe3_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe3_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe3_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe3_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe3_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe3_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe3_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe3_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe3_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe3_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe3_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe3_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe3_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe3_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe3_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe3_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe3_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe3_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe3_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe3_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe3_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe3_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe3_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe3_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe3_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe3_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe3_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe3_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe3_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe3_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe3_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe3_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe3_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe3_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe3_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe3_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe3_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe3_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe3_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe3_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe3_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe3_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe3_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe3_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe3_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe3_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe3_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe3_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe3_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe3_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe3_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe3_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe3_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe3_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe3_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe3_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe3_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe3_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe3_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe3_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe3_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe3_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe3_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe3_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe3_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe3_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe3_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe3_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe3_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe3_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe3_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe3_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe3_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe3_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe3_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe3_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe3_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe3_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe3_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe3_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe3_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe3_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe3_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe3_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe3_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe3_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe3_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe3_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe3_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe3_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe3_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe3_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe3_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe3_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe3_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe3_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe3_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe3_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe3_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe3_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe3_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe3_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe3_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe3_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe3_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe3_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe3_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe3_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe3_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe3_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe3_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe3_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe3_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe3_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe3_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe3_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe3_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe3_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe3_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe3_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe3_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe3_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe3_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe3_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe3_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe3_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe3_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe3_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe3_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe3_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe3_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe3_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe3_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe3_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe3_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe3_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe3_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe3_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe3_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe3_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe3_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe3_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe3_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe3_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe3_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe3_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe3_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe3_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe3_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe3_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe3_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe3_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe3_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe3_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe3_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe3_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe3_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe3_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe3_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe3_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe3_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe3_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe3_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe3_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe3_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe3_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe3_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe3_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe3_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe3_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe3_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe3_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe3_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe3_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe3_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe3_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe3_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe3_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe3_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe3_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe3_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe3_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe3_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe3_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe3_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe3_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe3_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe3_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe3_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe3_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe3_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe3_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe3_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe3_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe3_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe3_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe3_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe3_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe3_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe3_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe3_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe3_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe3_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe3_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe3_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe3_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe3_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe3_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe3_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe3_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe3_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe3_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe3_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe3_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe3_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe3_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe3_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe3_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe3_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe3_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe3_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe3_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe3_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe3_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe3_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe3_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe3_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe3_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe3_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe3_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe3_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe3_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe3_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe3_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe3_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe3_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe3_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe3_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe3_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe3_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe3_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe3_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe3_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe3_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe3_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe3_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe3_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe3_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe3_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe3_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe3_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe3_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe3_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe3_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe3_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe3_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe3_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe3_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe3_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe3_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe3_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe3_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe3_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe3_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe3_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe3_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe3_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe3_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe3_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe3_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe3_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe3_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe3_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe3_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe3_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe3_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe3_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe3_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe3_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe3_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe3_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe3_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe3_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe3_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe3_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe3_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe3_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe3_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe3_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe3_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe3_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe3_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe3_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe3_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe3_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe3_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe3_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe3_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe3_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe3_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe3_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe3_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe3_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe3_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe3_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe3_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe3_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe3_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe3_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe3_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe3_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe3_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe3_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe3_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe3_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe3_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe3_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe3_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe3_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe3_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe3_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe3_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe3_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe3_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe3_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe3_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe3_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe3_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe3_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe3_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe3_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe3_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe3_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe3_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe3_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe3_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe3_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe3_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe3_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe3_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe3_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe3_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe3_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe3_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe3_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe3_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe3_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe3_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe3_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe3_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe3_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe3_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe3_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe3_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe3_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe3_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe3_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe3_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe3_io_key_in),
    .io_key_out(pipe3_io_key_out),
    .io_sum_in(pipe3_io_sum_in),
    .io_sum_out(pipe3_io_sum_out)
  );
  HashSumLevel_3 pipe4 ( // @[hash.scala 130:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe4_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe4_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe4_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe4_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe4_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe4_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe4_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe4_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe4_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe4_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe4_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe4_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe4_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe4_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe4_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe4_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe4_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe4_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe4_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe4_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe4_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe4_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe4_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe4_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe4_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe4_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe4_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe4_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe4_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe4_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe4_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe4_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe4_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe4_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe4_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe4_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe4_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe4_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe4_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe4_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe4_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe4_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe4_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe4_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe4_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe4_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe4_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe4_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe4_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe4_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe4_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe4_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe4_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe4_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe4_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe4_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe4_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe4_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe4_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe4_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe4_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe4_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe4_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe4_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe4_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe4_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe4_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe4_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe4_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe4_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe4_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe4_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe4_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe4_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe4_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe4_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe4_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe4_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe4_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe4_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe4_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe4_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe4_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe4_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe4_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe4_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe4_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe4_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe4_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe4_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe4_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe4_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe4_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe4_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe4_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe4_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe4_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe4_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe4_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe4_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe4_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe4_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe4_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe4_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe4_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe4_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe4_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe4_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe4_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe4_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe4_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe4_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe4_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe4_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe4_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe4_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe4_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe4_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe4_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe4_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe4_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe4_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe4_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe4_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe4_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe4_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe4_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe4_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe4_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe4_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe4_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe4_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe4_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe4_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe4_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe4_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe4_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe4_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe4_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe4_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe4_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe4_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe4_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe4_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe4_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe4_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe4_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe4_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe4_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe4_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe4_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe4_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe4_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe4_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe4_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe4_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe4_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe4_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe4_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe4_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe4_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe4_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe4_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe4_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe4_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe4_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe4_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe4_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe4_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe4_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe4_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe4_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe4_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe4_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe4_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe4_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe4_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe4_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe4_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe4_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe4_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe4_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe4_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe4_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe4_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe4_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe4_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe4_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe4_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe4_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe4_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe4_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe4_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe4_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe4_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe4_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe4_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe4_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe4_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe4_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe4_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe4_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe4_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe4_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe4_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe4_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe4_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe4_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe4_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe4_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe4_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe4_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe4_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe4_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe4_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe4_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe4_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe4_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe4_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe4_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe4_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe4_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe4_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe4_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe4_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe4_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe4_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe4_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe4_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe4_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe4_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe4_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe4_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe4_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe4_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe4_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe4_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe4_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe4_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe4_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe4_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe4_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe4_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe4_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe4_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe4_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe4_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe4_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe4_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe4_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe4_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe4_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe4_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe4_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe4_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe4_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe4_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe4_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe4_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe4_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe4_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe4_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe4_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe4_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe4_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe4_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe4_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe4_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe4_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe4_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe4_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe4_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe4_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe4_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe4_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe4_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe4_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe4_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe4_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe4_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe4_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe4_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe4_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe4_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe4_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe4_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe4_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe4_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe4_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe4_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe4_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe4_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe4_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe4_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe4_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe4_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe4_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe4_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe4_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe4_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe4_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe4_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe4_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe4_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe4_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe4_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe4_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe4_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe4_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe4_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe4_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe4_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe4_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe4_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe4_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe4_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe4_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe4_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe4_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe4_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe4_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe4_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe4_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe4_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe4_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe4_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe4_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe4_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe4_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe4_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe4_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe4_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe4_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe4_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe4_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe4_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe4_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe4_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe4_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe4_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe4_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe4_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe4_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe4_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe4_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe4_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe4_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe4_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe4_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe4_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe4_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe4_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe4_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe4_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe4_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe4_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe4_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe4_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe4_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe4_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe4_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe4_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe4_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe4_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe4_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe4_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe4_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe4_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe4_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe4_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe4_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe4_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe4_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe4_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe4_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe4_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe4_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe4_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe4_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe4_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe4_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe4_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe4_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe4_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe4_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe4_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe4_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe4_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe4_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe4_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe4_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe4_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe4_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe4_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe4_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe4_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe4_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe4_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe4_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe4_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe4_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe4_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe4_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe4_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe4_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe4_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe4_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe4_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe4_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe4_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe4_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe4_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe4_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe4_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe4_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe4_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe4_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe4_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe4_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe4_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe4_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe4_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe4_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe4_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe4_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe4_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe4_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe4_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe4_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe4_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe4_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe4_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe4_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe4_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe4_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe4_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe4_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe4_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe4_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe4_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe4_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe4_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe4_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe4_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe4_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe4_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe4_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe4_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe4_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe4_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe4_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe4_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe4_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe4_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe4_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe4_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe4_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe4_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe4_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe4_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe4_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe4_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe4_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe4_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe4_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe4_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe4_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe4_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe4_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe4_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe4_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe4_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe4_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe4_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe4_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe4_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe4_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe4_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe4_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe4_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe4_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe4_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe4_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe4_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe4_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe4_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe4_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe4_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe4_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe4_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe4_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe4_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe4_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe4_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe4_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe4_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe4_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe4_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe4_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe4_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe4_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe4_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe4_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe4_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe4_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe4_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe4_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe4_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe4_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe4_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe4_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe4_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe4_io_key_in),
    .io_key_out(pipe4_io_key_out),
    .io_sum_in(pipe4_io_sum_in),
    .io_sum_out(pipe4_io_sum_out)
  );
  HashReshapeLevel pipe5 ( // @[hash.scala 131:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe5_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe5_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe5_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe5_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe5_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe5_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe5_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe5_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe5_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe5_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe5_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe5_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe5_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe5_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe5_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe5_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe5_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe5_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe5_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe5_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe5_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe5_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe5_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe5_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe5_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe5_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe5_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe5_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe5_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe5_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe5_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe5_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe5_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe5_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe5_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe5_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe5_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe5_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe5_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe5_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe5_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe5_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe5_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe5_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe5_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe5_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe5_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe5_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe5_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe5_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe5_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe5_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe5_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe5_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe5_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe5_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe5_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe5_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe5_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe5_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe5_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe5_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe5_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe5_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe5_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe5_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe5_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe5_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe5_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe5_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe5_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe5_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe5_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe5_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe5_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe5_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe5_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe5_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe5_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe5_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe5_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe5_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe5_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe5_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe5_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe5_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe5_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe5_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe5_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe5_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe5_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe5_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe5_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe5_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe5_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe5_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe5_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe5_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe5_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe5_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe5_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe5_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe5_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe5_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe5_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe5_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe5_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe5_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe5_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe5_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe5_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe5_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe5_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe5_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe5_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe5_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe5_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe5_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe5_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe5_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe5_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe5_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe5_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe5_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe5_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe5_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe5_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe5_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe5_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe5_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe5_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe5_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe5_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe5_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe5_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe5_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe5_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe5_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe5_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe5_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe5_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe5_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe5_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe5_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe5_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe5_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe5_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe5_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe5_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe5_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe5_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe5_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe5_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe5_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe5_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe5_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe5_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe5_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe5_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe5_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe5_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe5_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe5_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe5_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe5_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe5_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe5_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe5_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe5_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe5_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe5_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe5_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe5_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe5_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe5_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe5_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe5_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe5_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe5_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe5_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe5_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe5_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe5_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe5_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe5_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe5_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe5_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe5_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe5_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe5_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe5_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe5_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe5_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe5_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe5_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe5_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe5_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe5_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe5_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe5_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe5_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe5_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe5_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe5_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe5_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe5_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe5_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe5_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe5_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe5_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe5_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe5_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe5_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe5_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe5_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe5_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe5_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe5_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe5_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe5_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe5_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe5_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe5_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe5_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe5_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe5_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe5_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe5_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe5_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe5_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe5_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe5_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe5_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe5_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe5_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe5_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe5_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe5_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe5_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe5_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe5_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe5_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe5_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe5_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe5_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe5_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe5_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe5_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe5_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe5_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe5_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe5_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe5_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe5_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe5_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe5_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe5_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe5_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe5_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe5_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe5_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe5_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe5_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe5_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe5_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe5_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe5_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe5_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe5_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe5_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe5_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe5_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe5_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe5_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe5_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe5_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe5_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe5_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe5_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe5_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe5_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe5_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe5_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe5_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe5_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe5_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe5_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe5_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe5_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe5_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe5_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe5_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe5_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe5_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe5_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe5_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe5_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe5_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe5_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe5_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe5_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe5_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe5_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe5_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe5_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe5_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe5_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe5_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe5_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe5_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe5_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe5_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe5_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe5_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe5_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe5_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe5_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe5_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe5_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe5_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe5_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe5_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe5_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe5_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe5_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe5_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe5_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe5_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe5_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe5_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe5_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe5_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe5_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe5_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe5_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe5_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe5_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe5_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe5_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe5_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe5_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe5_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe5_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe5_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe5_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe5_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe5_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe5_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe5_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe5_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe5_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe5_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe5_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe5_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe5_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe5_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe5_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe5_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe5_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe5_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe5_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe5_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe5_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe5_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe5_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe5_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe5_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe5_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe5_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe5_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe5_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe5_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe5_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe5_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe5_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe5_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe5_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe5_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe5_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe5_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe5_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe5_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe5_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe5_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe5_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe5_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe5_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe5_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe5_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe5_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe5_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe5_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe5_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe5_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe5_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe5_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe5_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe5_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe5_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe5_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe5_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe5_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe5_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe5_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe5_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe5_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe5_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe5_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe5_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe5_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe5_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe5_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe5_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe5_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe5_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe5_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe5_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe5_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe5_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe5_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe5_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe5_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe5_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe5_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe5_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe5_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe5_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe5_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe5_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe5_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe5_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe5_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe5_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe5_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe5_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe5_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe5_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe5_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe5_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe5_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe5_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe5_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe5_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe5_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe5_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe5_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe5_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe5_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe5_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe5_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe5_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe5_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe5_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe5_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe5_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe5_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe5_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe5_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe5_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe5_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe5_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe5_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe5_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe5_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe5_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe5_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe5_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe5_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe5_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe5_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe5_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe5_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe5_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe5_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe5_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe5_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe5_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe5_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe5_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe5_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe5_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe5_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe5_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe5_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe5_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe5_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe5_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe5_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe5_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe5_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe5_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe5_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe5_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe5_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe5_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe5_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe5_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe5_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe5_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe5_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe5_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe5_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe5_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe5_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe5_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe5_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe5_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe5_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe5_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe5_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe5_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe5_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe5_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe5_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe5_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe5_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe5_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe5_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe5_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe5_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe5_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe5_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe5_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe5_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe5_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe5_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe5_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe5_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe5_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe5_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe5_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe5_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe5_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe5_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe5_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe5_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe5_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe5_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe5_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe5_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe5_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe5_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe5_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe5_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe5_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe5_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe5_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe5_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe5_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe5_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe5_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe5_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe5_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe5_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe5_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe5_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe5_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe5_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe5_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe5_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe5_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe5_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe5_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe5_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe5_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe5_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe5_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe5_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe5_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe5_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe5_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe5_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe5_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe5_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe5_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe5_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe5_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe5_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe5_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe5_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe5_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe5_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe5_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe5_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe5_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe5_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe5_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe5_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe5_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe5_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe5_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe5_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe5_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe5_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe5_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe5_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe5_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe5_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe5_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe5_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe5_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe5_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe5_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe5_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe5_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe5_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe5_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe5_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe5_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe5_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe5_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe5_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe5_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe5_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe5_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe5_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe5_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe5_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe5_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe5_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe5_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe5_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe5_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe5_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe5_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe5_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe5_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe5_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe5_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe5_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe5_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe5_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe5_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe5_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe5_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe5_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe5_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe5_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe5_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe5_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe5_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe5_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe5_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe5_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe5_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe5_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe5_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe5_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe5_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe5_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe5_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe5_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe5_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe5_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe5_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe5_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe5_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe5_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe5_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe5_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe5_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe5_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe5_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe5_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe5_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe5_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe5_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe5_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe5_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe5_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe5_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe5_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe5_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe5_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe5_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe5_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe5_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe5_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe5_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe5_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe5_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe5_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe5_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe5_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe5_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe5_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe5_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe5_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe5_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe5_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe5_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe5_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe5_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe5_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe5_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe5_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe5_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe5_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe5_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe5_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe5_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe5_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe5_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe5_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe5_io_hash_depth_0),
    .io_hash_depth_1(pipe5_io_hash_depth_1),
    .io_key_in(pipe5_io_key_in),
    .io_key_out(pipe5_io_key_out),
    .io_sum_in(pipe5_io_sum_in),
    .io_sum_out(pipe5_io_sum_out),
    .io_val_out(pipe5_io_val_out)
  );
  HashReshapeLevel_1 pipe6 ( // @[hash.scala 132:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe6_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe6_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe6_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe6_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe6_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe6_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe6_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe6_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe6_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe6_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe6_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe6_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe6_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe6_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe6_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe6_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe6_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe6_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe6_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe6_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe6_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe6_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe6_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe6_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe6_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe6_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe6_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe6_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe6_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe6_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe6_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe6_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe6_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe6_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe6_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe6_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe6_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe6_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe6_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe6_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe6_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe6_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe6_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe6_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe6_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe6_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe6_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe6_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe6_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe6_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe6_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe6_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe6_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe6_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe6_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe6_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe6_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe6_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe6_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe6_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe6_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe6_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe6_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe6_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe6_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe6_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe6_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe6_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe6_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe6_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe6_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe6_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe6_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe6_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe6_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe6_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe6_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe6_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe6_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe6_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe6_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe6_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe6_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe6_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe6_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe6_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe6_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe6_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe6_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe6_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe6_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe6_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe6_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe6_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe6_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe6_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe6_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe6_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe6_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe6_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe6_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe6_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe6_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe6_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe6_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe6_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe6_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe6_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe6_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe6_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe6_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe6_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe6_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe6_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe6_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe6_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe6_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe6_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe6_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe6_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe6_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe6_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe6_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe6_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe6_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe6_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe6_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe6_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe6_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe6_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe6_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe6_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe6_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe6_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe6_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe6_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe6_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe6_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe6_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe6_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe6_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe6_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe6_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe6_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe6_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe6_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe6_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe6_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe6_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe6_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe6_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe6_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe6_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe6_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe6_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe6_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe6_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe6_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe6_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe6_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe6_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe6_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe6_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe6_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe6_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe6_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe6_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe6_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe6_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe6_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe6_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe6_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe6_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe6_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe6_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe6_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe6_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe6_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe6_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe6_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe6_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe6_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe6_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe6_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe6_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe6_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe6_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe6_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe6_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe6_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe6_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe6_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe6_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe6_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe6_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe6_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe6_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe6_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe6_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe6_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe6_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe6_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe6_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe6_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe6_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe6_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe6_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe6_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe6_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe6_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe6_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe6_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe6_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe6_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe6_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe6_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe6_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe6_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe6_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe6_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe6_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe6_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe6_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe6_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe6_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe6_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe6_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe6_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe6_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe6_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe6_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe6_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe6_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe6_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe6_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe6_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe6_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe6_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe6_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe6_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe6_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe6_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe6_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe6_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe6_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe6_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe6_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe6_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe6_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe6_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe6_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe6_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe6_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe6_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe6_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe6_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe6_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe6_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe6_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe6_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe6_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe6_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe6_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe6_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe6_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe6_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe6_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe6_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe6_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe6_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe6_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe6_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe6_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe6_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe6_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe6_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe6_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe6_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe6_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe6_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe6_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe6_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe6_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe6_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe6_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe6_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe6_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe6_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe6_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe6_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe6_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe6_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe6_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe6_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe6_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe6_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe6_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe6_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe6_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe6_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe6_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe6_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe6_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe6_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe6_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe6_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe6_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe6_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe6_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe6_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe6_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe6_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe6_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe6_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe6_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe6_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe6_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe6_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe6_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe6_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe6_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe6_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe6_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe6_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe6_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe6_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe6_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe6_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe6_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe6_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe6_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe6_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe6_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe6_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe6_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe6_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe6_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe6_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe6_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe6_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe6_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe6_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe6_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe6_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe6_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe6_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe6_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe6_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe6_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe6_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe6_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe6_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe6_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe6_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe6_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe6_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe6_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe6_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe6_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe6_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe6_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe6_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe6_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe6_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe6_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe6_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe6_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe6_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe6_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe6_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe6_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe6_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe6_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe6_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe6_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe6_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe6_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe6_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe6_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe6_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe6_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe6_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe6_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe6_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe6_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe6_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe6_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe6_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe6_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe6_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe6_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe6_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe6_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe6_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe6_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe6_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe6_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe6_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe6_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe6_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe6_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe6_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe6_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe6_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe6_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe6_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe6_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe6_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe6_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe6_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe6_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe6_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe6_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe6_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe6_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe6_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe6_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe6_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe6_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe6_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe6_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe6_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe6_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe6_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe6_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe6_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe6_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe6_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe6_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe6_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe6_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe6_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe6_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe6_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe6_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe6_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe6_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe6_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe6_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe6_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe6_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe6_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe6_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe6_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe6_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe6_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe6_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe6_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe6_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe6_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe6_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe6_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe6_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe6_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe6_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe6_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe6_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe6_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe6_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe6_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe6_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe6_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe6_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe6_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe6_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe6_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe6_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe6_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe6_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe6_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe6_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe6_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe6_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe6_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe6_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe6_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe6_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe6_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe6_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe6_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe6_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe6_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe6_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe6_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe6_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe6_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe6_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe6_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe6_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe6_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe6_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe6_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe6_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe6_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe6_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe6_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe6_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe6_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe6_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe6_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe6_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe6_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe6_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe6_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe6_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe6_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe6_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe6_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe6_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe6_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe6_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe6_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe6_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe6_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe6_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe6_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe6_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe6_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe6_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe6_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe6_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe6_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe6_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe6_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe6_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe6_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe6_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe6_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe6_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe6_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe6_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe6_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe6_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe6_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe6_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe6_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe6_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe6_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe6_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe6_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe6_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe6_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe6_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe6_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe6_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe6_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe6_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe6_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe6_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe6_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe6_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe6_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe6_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe6_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe6_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe6_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe6_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe6_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe6_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe6_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe6_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe6_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe6_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe6_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe6_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe6_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe6_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe6_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe6_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe6_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe6_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe6_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe6_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe6_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe6_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe6_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe6_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe6_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe6_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe6_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe6_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe6_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe6_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe6_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe6_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe6_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe6_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe6_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe6_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe6_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe6_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe6_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe6_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe6_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe6_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe6_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe6_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe6_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe6_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe6_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe6_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe6_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe6_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe6_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe6_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe6_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe6_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe6_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe6_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe6_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe6_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe6_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe6_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe6_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe6_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe6_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe6_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe6_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe6_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe6_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe6_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe6_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe6_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe6_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe6_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe6_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe6_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe6_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe6_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe6_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe6_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe6_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe6_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe6_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe6_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe6_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe6_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe6_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe6_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe6_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe6_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe6_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe6_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe6_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe6_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe6_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe6_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe6_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe6_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe6_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe6_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe6_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe6_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe6_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe6_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe6_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe6_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe6_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe6_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe6_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe6_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe6_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe6_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe6_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe6_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe6_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe6_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe6_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe6_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe6_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe6_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe6_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe6_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe6_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe6_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe6_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe6_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe6_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe6_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe6_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe6_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe6_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe6_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe6_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe6_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe6_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe6_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe6_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe6_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe6_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe6_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe6_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe6_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe6_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe6_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe6_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe6_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe6_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe6_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe6_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe6_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe6_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe6_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe6_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe6_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe6_io_hash_depth_0),
    .io_hash_depth_1(pipe6_io_hash_depth_1),
    .io_key_in(pipe6_io_key_in),
    .io_key_out(pipe6_io_key_out),
    .io_sum_in(pipe6_io_sum_in),
    .io_sum_out(pipe6_io_sum_out),
    .io_val_in(pipe6_io_val_in),
    .io_val_out(pipe6_io_val_out)
  );
  HashReshapeLevel_2 pipe7 ( // @[hash.scala 133:23]
    .clock(pipe7_clock),
    .io_pipe_phv_in_data_0(pipe7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe7_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe7_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe7_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe7_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe7_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe7_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe7_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe7_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe7_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe7_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe7_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe7_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe7_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe7_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe7_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe7_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe7_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe7_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe7_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe7_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe7_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe7_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe7_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe7_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe7_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe7_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe7_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe7_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe7_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe7_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe7_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe7_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe7_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe7_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe7_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe7_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe7_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe7_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe7_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe7_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe7_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe7_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe7_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe7_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe7_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe7_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe7_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe7_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe7_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe7_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe7_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe7_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe7_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe7_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe7_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe7_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe7_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe7_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe7_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe7_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe7_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe7_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe7_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe7_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe7_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe7_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe7_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe7_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe7_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe7_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe7_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe7_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe7_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe7_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe7_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe7_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe7_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe7_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe7_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe7_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe7_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe7_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe7_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe7_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe7_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe7_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe7_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe7_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe7_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe7_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe7_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe7_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe7_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe7_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe7_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe7_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe7_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe7_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe7_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe7_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe7_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe7_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe7_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe7_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe7_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe7_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe7_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe7_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe7_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe7_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe7_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe7_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe7_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe7_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe7_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe7_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe7_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe7_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe7_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe7_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe7_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe7_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe7_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe7_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe7_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe7_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe7_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe7_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe7_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe7_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe7_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe7_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe7_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe7_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe7_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe7_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe7_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe7_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe7_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe7_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe7_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe7_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe7_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe7_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe7_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe7_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe7_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe7_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe7_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe7_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe7_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe7_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe7_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe7_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe7_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe7_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe7_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe7_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe7_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe7_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe7_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe7_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe7_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe7_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe7_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe7_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe7_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe7_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe7_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe7_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe7_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe7_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe7_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe7_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe7_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe7_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe7_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe7_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe7_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe7_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe7_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe7_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe7_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe7_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe7_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe7_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe7_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe7_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe7_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe7_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe7_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe7_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe7_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe7_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe7_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe7_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe7_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe7_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe7_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe7_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe7_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe7_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe7_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe7_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe7_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe7_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe7_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe7_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe7_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe7_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe7_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe7_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe7_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe7_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe7_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe7_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe7_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe7_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe7_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe7_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe7_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe7_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe7_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe7_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe7_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe7_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe7_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe7_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe7_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe7_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe7_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe7_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe7_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe7_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe7_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe7_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe7_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe7_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe7_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe7_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe7_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe7_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe7_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe7_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe7_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe7_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe7_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe7_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe7_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe7_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe7_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe7_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe7_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe7_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe7_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe7_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe7_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe7_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe7_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe7_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe7_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe7_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe7_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe7_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe7_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe7_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe7_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe7_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe7_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe7_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe7_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe7_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe7_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe7_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe7_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe7_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe7_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe7_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe7_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe7_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe7_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe7_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe7_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe7_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe7_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe7_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe7_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe7_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe7_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe7_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe7_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe7_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe7_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe7_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe7_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe7_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe7_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe7_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe7_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe7_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe7_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe7_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe7_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe7_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe7_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe7_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe7_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe7_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe7_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe7_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe7_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe7_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe7_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe7_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe7_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe7_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe7_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe7_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe7_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe7_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe7_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe7_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe7_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe7_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe7_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe7_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe7_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe7_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe7_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe7_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe7_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe7_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe7_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe7_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe7_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe7_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe7_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe7_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe7_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe7_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe7_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe7_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe7_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe7_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe7_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe7_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe7_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe7_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe7_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe7_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe7_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe7_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe7_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe7_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe7_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe7_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe7_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe7_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe7_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe7_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe7_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe7_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe7_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe7_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe7_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe7_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe7_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe7_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe7_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe7_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe7_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe7_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe7_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe7_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe7_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe7_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe7_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe7_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe7_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe7_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe7_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe7_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe7_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe7_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe7_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe7_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe7_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe7_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe7_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe7_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe7_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe7_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe7_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe7_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe7_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe7_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe7_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe7_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe7_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe7_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe7_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe7_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe7_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe7_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe7_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe7_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe7_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe7_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe7_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe7_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe7_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe7_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe7_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe7_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe7_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe7_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe7_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe7_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe7_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe7_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe7_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe7_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe7_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe7_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe7_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe7_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe7_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe7_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe7_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe7_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe7_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe7_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe7_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe7_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe7_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe7_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe7_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe7_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe7_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe7_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe7_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe7_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe7_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe7_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe7_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe7_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe7_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe7_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe7_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe7_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe7_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe7_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe7_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe7_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe7_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe7_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe7_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe7_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe7_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe7_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe7_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe7_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe7_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe7_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe7_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe7_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe7_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe7_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe7_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe7_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe7_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe7_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe7_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe7_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe7_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe7_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe7_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe7_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe7_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe7_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe7_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe7_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe7_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe7_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe7_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe7_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe7_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe7_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe7_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe7_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe7_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe7_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe7_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe7_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe7_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe7_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe7_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe7_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe7_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe7_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe7_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe7_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe7_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe7_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe7_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe7_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe7_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe7_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe7_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe7_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe7_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe7_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe7_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe7_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe7_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe7_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe7_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe7_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe7_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe7_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe7_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe7_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe7_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe7_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe7_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe7_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe7_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe7_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe7_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe7_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe7_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe7_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe7_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe7_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe7_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe7_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe7_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe7_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe7_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe7_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe7_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe7_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe7_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe7_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe7_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe7_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe7_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe7_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe7_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe7_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe7_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe7_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe7_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe7_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe7_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe7_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe7_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe7_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe7_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe7_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe7_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe7_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe7_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe7_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe7_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe7_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe7_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe7_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe7_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe7_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe7_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe7_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe7_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe7_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe7_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe7_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe7_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe7_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe7_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe7_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe7_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe7_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe7_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe7_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe7_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe7_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe7_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe7_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe7_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe7_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe7_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe7_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe7_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe7_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe7_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe7_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe7_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe7_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe7_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe7_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe7_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe7_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe7_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe7_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe7_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe7_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe7_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe7_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe7_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe7_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe7_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe7_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe7_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe7_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe7_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe7_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe7_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe7_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe7_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe7_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe7_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe7_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe7_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe7_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe7_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe7_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe7_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe7_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe7_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe7_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe7_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe7_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe7_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe7_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe7_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe7_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe7_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe7_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe7_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe7_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe7_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe7_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe7_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe7_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe7_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe7_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe7_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe7_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe7_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe7_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe7_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe7_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe7_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe7_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe7_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe7_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe7_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe7_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe7_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe7_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe7_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe7_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe7_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe7_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe7_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe7_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe7_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe7_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe7_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe7_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe7_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe7_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe7_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe7_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe7_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe7_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe7_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe7_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe7_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe7_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe7_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe7_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe7_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe7_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe7_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe7_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe7_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe7_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe7_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe7_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe7_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe7_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe7_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe7_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe7_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe7_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe7_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe7_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe7_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe7_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe7_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe7_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe7_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe7_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe7_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe7_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe7_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe7_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe7_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe7_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe7_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe7_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe7_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe7_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe7_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe7_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe7_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe7_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe7_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe7_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe7_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe7_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe7_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe7_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe7_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe7_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe7_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe7_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe7_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe7_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe7_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe7_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe7_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe7_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe7_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe7_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe7_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe7_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe7_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe7_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe7_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe7_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe7_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe7_io_hash_depth_0),
    .io_hash_depth_1(pipe7_io_hash_depth_1),
    .io_key_in(pipe7_io_key_in),
    .io_key_out(pipe7_io_key_out),
    .io_sum_in(pipe7_io_sum_in),
    .io_sum_out(pipe7_io_sum_out),
    .io_val_in(pipe7_io_val_in),
    .io_val_out(pipe7_io_val_out)
  );
  HashReshapeLevel_3 pipe8 ( // @[hash.scala 134:23]
    .clock(pipe8_clock),
    .io_pipe_phv_in_data_0(pipe8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe8_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe8_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe8_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe8_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe8_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe8_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe8_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe8_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe8_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe8_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe8_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe8_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe8_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe8_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe8_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe8_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe8_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe8_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe8_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe8_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe8_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe8_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe8_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe8_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe8_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe8_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe8_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe8_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe8_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe8_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe8_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe8_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe8_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe8_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe8_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe8_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe8_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe8_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe8_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe8_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe8_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe8_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe8_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe8_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe8_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe8_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe8_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe8_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe8_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe8_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe8_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe8_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe8_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe8_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe8_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe8_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe8_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe8_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe8_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe8_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe8_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe8_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe8_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe8_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe8_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe8_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe8_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe8_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe8_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe8_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe8_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe8_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe8_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe8_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe8_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe8_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe8_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe8_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe8_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe8_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe8_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe8_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe8_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe8_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe8_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe8_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe8_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe8_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe8_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe8_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe8_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe8_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe8_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe8_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe8_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe8_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe8_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe8_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe8_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe8_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe8_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe8_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe8_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe8_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe8_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe8_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe8_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe8_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe8_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe8_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe8_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe8_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe8_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe8_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe8_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe8_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe8_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe8_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe8_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe8_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe8_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe8_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe8_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe8_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe8_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe8_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe8_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe8_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe8_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe8_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe8_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe8_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe8_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe8_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe8_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe8_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe8_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe8_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe8_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe8_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe8_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe8_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe8_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe8_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe8_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe8_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe8_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe8_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe8_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe8_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe8_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe8_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe8_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe8_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe8_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe8_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe8_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe8_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe8_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe8_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe8_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe8_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe8_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe8_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe8_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe8_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe8_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe8_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe8_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe8_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe8_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe8_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe8_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe8_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe8_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe8_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe8_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe8_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe8_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe8_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe8_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe8_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe8_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe8_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe8_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe8_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe8_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe8_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe8_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe8_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe8_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe8_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe8_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe8_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe8_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe8_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe8_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe8_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe8_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe8_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe8_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe8_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe8_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe8_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe8_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe8_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe8_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe8_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe8_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe8_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe8_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe8_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe8_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe8_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe8_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe8_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe8_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe8_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe8_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe8_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe8_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe8_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe8_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe8_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe8_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe8_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe8_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe8_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe8_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe8_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe8_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe8_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe8_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe8_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe8_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe8_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe8_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe8_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe8_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe8_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe8_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe8_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe8_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe8_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe8_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe8_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe8_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe8_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe8_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe8_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe8_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe8_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe8_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe8_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe8_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe8_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe8_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe8_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe8_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe8_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe8_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe8_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe8_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe8_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe8_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe8_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe8_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe8_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe8_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe8_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe8_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe8_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe8_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe8_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe8_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe8_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe8_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe8_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe8_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe8_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe8_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe8_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe8_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe8_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe8_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe8_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe8_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe8_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe8_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe8_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe8_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe8_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe8_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe8_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe8_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe8_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe8_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe8_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe8_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe8_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe8_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe8_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe8_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe8_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe8_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe8_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe8_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe8_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe8_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe8_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe8_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe8_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe8_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe8_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe8_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe8_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe8_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe8_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe8_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe8_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe8_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe8_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe8_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe8_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe8_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe8_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe8_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe8_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe8_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe8_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe8_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe8_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe8_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe8_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe8_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe8_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe8_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe8_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe8_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe8_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe8_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe8_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe8_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe8_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe8_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe8_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe8_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe8_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe8_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe8_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe8_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe8_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe8_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe8_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe8_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe8_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe8_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe8_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe8_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe8_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe8_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe8_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe8_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe8_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe8_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe8_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe8_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe8_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe8_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe8_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe8_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe8_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe8_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe8_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe8_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe8_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe8_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe8_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe8_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe8_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe8_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe8_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe8_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe8_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe8_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe8_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe8_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe8_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe8_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe8_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe8_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe8_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe8_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe8_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe8_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe8_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe8_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe8_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe8_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe8_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe8_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe8_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe8_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe8_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe8_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe8_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe8_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe8_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe8_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe8_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe8_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe8_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe8_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe8_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe8_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe8_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe8_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe8_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe8_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe8_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe8_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe8_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe8_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe8_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe8_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe8_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe8_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe8_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe8_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe8_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe8_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe8_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe8_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe8_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe8_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe8_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe8_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe8_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe8_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe8_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe8_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe8_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe8_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe8_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe8_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe8_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe8_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe8_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe8_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe8_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe8_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe8_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe8_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe8_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe8_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe8_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe8_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe8_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe8_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe8_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe8_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe8_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe8_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe8_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe8_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe8_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe8_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe8_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe8_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe8_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe8_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe8_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe8_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe8_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe8_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe8_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe8_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe8_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe8_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe8_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe8_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe8_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe8_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe8_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe8_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe8_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe8_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe8_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe8_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe8_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe8_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe8_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe8_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe8_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe8_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe8_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe8_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe8_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe8_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe8_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe8_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe8_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe8_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe8_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe8_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe8_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe8_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe8_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe8_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe8_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe8_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe8_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe8_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe8_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe8_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe8_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe8_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe8_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe8_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe8_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe8_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe8_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe8_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe8_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe8_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe8_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe8_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe8_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe8_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe8_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe8_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe8_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe8_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe8_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe8_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe8_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe8_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe8_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe8_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe8_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe8_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe8_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe8_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe8_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe8_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe8_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe8_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe8_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe8_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe8_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe8_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe8_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe8_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe8_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe8_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe8_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe8_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe8_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe8_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe8_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe8_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe8_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe8_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe8_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe8_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe8_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe8_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe8_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe8_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe8_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe8_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe8_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe8_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe8_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe8_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe8_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe8_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe8_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe8_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe8_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe8_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe8_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe8_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe8_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe8_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe8_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe8_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe8_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe8_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe8_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe8_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe8_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe8_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe8_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe8_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe8_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe8_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe8_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe8_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe8_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe8_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe8_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe8_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe8_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe8_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe8_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe8_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe8_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe8_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe8_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe8_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe8_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe8_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe8_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe8_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe8_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe8_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe8_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe8_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe8_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe8_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe8_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe8_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe8_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe8_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe8_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe8_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe8_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe8_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe8_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe8_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe8_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe8_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe8_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe8_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe8_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe8_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe8_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe8_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe8_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe8_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe8_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe8_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe8_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe8_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe8_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe8_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe8_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe8_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe8_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe8_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe8_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe8_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe8_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe8_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe8_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe8_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe8_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe8_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe8_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe8_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe8_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe8_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe8_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe8_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe8_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe8_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe8_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe8_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe8_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe8_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe8_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe8_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe8_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe8_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe8_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe8_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe8_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe8_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe8_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe8_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe8_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe8_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe8_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe8_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe8_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe8_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe8_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe8_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe8_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe8_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe8_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe8_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe8_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe8_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe8_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe8_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe8_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe8_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe8_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe8_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe8_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe8_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe8_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe8_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe8_io_hash_depth_0),
    .io_hash_depth_1(pipe8_io_hash_depth_1),
    .io_key_in(pipe8_io_key_in),
    .io_key_out(pipe8_io_key_out),
    .io_sum_in(pipe8_io_sum_in),
    .io_sum_out(pipe8_io_sum_out),
    .io_val_in(pipe8_io_val_in),
    .io_val_out(pipe8_io_val_out)
  );
  assign io_pipe_phv_out_data_0 = pipe8_io_pipe_phv_out_data_0; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_1 = pipe8_io_pipe_phv_out_data_1; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_2 = pipe8_io_pipe_phv_out_data_2; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_3 = pipe8_io_pipe_phv_out_data_3; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_4 = pipe8_io_pipe_phv_out_data_4; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_5 = pipe8_io_pipe_phv_out_data_5; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_6 = pipe8_io_pipe_phv_out_data_6; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_7 = pipe8_io_pipe_phv_out_data_7; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_8 = pipe8_io_pipe_phv_out_data_8; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_9 = pipe8_io_pipe_phv_out_data_9; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_10 = pipe8_io_pipe_phv_out_data_10; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_11 = pipe8_io_pipe_phv_out_data_11; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_12 = pipe8_io_pipe_phv_out_data_12; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_13 = pipe8_io_pipe_phv_out_data_13; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_14 = pipe8_io_pipe_phv_out_data_14; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_15 = pipe8_io_pipe_phv_out_data_15; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_16 = pipe8_io_pipe_phv_out_data_16; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_17 = pipe8_io_pipe_phv_out_data_17; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_18 = pipe8_io_pipe_phv_out_data_18; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_19 = pipe8_io_pipe_phv_out_data_19; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_20 = pipe8_io_pipe_phv_out_data_20; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_21 = pipe8_io_pipe_phv_out_data_21; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_22 = pipe8_io_pipe_phv_out_data_22; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_23 = pipe8_io_pipe_phv_out_data_23; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_24 = pipe8_io_pipe_phv_out_data_24; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_25 = pipe8_io_pipe_phv_out_data_25; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_26 = pipe8_io_pipe_phv_out_data_26; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_27 = pipe8_io_pipe_phv_out_data_27; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_28 = pipe8_io_pipe_phv_out_data_28; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_29 = pipe8_io_pipe_phv_out_data_29; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_30 = pipe8_io_pipe_phv_out_data_30; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_31 = pipe8_io_pipe_phv_out_data_31; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_32 = pipe8_io_pipe_phv_out_data_32; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_33 = pipe8_io_pipe_phv_out_data_33; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_34 = pipe8_io_pipe_phv_out_data_34; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_35 = pipe8_io_pipe_phv_out_data_35; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_36 = pipe8_io_pipe_phv_out_data_36; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_37 = pipe8_io_pipe_phv_out_data_37; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_38 = pipe8_io_pipe_phv_out_data_38; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_39 = pipe8_io_pipe_phv_out_data_39; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_40 = pipe8_io_pipe_phv_out_data_40; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_41 = pipe8_io_pipe_phv_out_data_41; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_42 = pipe8_io_pipe_phv_out_data_42; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_43 = pipe8_io_pipe_phv_out_data_43; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_44 = pipe8_io_pipe_phv_out_data_44; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_45 = pipe8_io_pipe_phv_out_data_45; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_46 = pipe8_io_pipe_phv_out_data_46; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_47 = pipe8_io_pipe_phv_out_data_47; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_48 = pipe8_io_pipe_phv_out_data_48; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_49 = pipe8_io_pipe_phv_out_data_49; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_50 = pipe8_io_pipe_phv_out_data_50; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_51 = pipe8_io_pipe_phv_out_data_51; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_52 = pipe8_io_pipe_phv_out_data_52; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_53 = pipe8_io_pipe_phv_out_data_53; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_54 = pipe8_io_pipe_phv_out_data_54; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_55 = pipe8_io_pipe_phv_out_data_55; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_56 = pipe8_io_pipe_phv_out_data_56; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_57 = pipe8_io_pipe_phv_out_data_57; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_58 = pipe8_io_pipe_phv_out_data_58; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_59 = pipe8_io_pipe_phv_out_data_59; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_60 = pipe8_io_pipe_phv_out_data_60; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_61 = pipe8_io_pipe_phv_out_data_61; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_62 = pipe8_io_pipe_phv_out_data_62; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_63 = pipe8_io_pipe_phv_out_data_63; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_64 = pipe8_io_pipe_phv_out_data_64; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_65 = pipe8_io_pipe_phv_out_data_65; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_66 = pipe8_io_pipe_phv_out_data_66; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_67 = pipe8_io_pipe_phv_out_data_67; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_68 = pipe8_io_pipe_phv_out_data_68; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_69 = pipe8_io_pipe_phv_out_data_69; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_70 = pipe8_io_pipe_phv_out_data_70; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_71 = pipe8_io_pipe_phv_out_data_71; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_72 = pipe8_io_pipe_phv_out_data_72; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_73 = pipe8_io_pipe_phv_out_data_73; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_74 = pipe8_io_pipe_phv_out_data_74; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_75 = pipe8_io_pipe_phv_out_data_75; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_76 = pipe8_io_pipe_phv_out_data_76; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_77 = pipe8_io_pipe_phv_out_data_77; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_78 = pipe8_io_pipe_phv_out_data_78; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_79 = pipe8_io_pipe_phv_out_data_79; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_80 = pipe8_io_pipe_phv_out_data_80; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_81 = pipe8_io_pipe_phv_out_data_81; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_82 = pipe8_io_pipe_phv_out_data_82; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_83 = pipe8_io_pipe_phv_out_data_83; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_84 = pipe8_io_pipe_phv_out_data_84; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_85 = pipe8_io_pipe_phv_out_data_85; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_86 = pipe8_io_pipe_phv_out_data_86; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_87 = pipe8_io_pipe_phv_out_data_87; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_88 = pipe8_io_pipe_phv_out_data_88; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_89 = pipe8_io_pipe_phv_out_data_89; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_90 = pipe8_io_pipe_phv_out_data_90; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_91 = pipe8_io_pipe_phv_out_data_91; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_92 = pipe8_io_pipe_phv_out_data_92; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_93 = pipe8_io_pipe_phv_out_data_93; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_94 = pipe8_io_pipe_phv_out_data_94; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_95 = pipe8_io_pipe_phv_out_data_95; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_96 = pipe8_io_pipe_phv_out_data_96; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_97 = pipe8_io_pipe_phv_out_data_97; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_98 = pipe8_io_pipe_phv_out_data_98; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_99 = pipe8_io_pipe_phv_out_data_99; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_100 = pipe8_io_pipe_phv_out_data_100; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_101 = pipe8_io_pipe_phv_out_data_101; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_102 = pipe8_io_pipe_phv_out_data_102; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_103 = pipe8_io_pipe_phv_out_data_103; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_104 = pipe8_io_pipe_phv_out_data_104; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_105 = pipe8_io_pipe_phv_out_data_105; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_106 = pipe8_io_pipe_phv_out_data_106; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_107 = pipe8_io_pipe_phv_out_data_107; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_108 = pipe8_io_pipe_phv_out_data_108; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_109 = pipe8_io_pipe_phv_out_data_109; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_110 = pipe8_io_pipe_phv_out_data_110; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_111 = pipe8_io_pipe_phv_out_data_111; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_112 = pipe8_io_pipe_phv_out_data_112; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_113 = pipe8_io_pipe_phv_out_data_113; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_114 = pipe8_io_pipe_phv_out_data_114; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_115 = pipe8_io_pipe_phv_out_data_115; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_116 = pipe8_io_pipe_phv_out_data_116; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_117 = pipe8_io_pipe_phv_out_data_117; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_118 = pipe8_io_pipe_phv_out_data_118; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_119 = pipe8_io_pipe_phv_out_data_119; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_120 = pipe8_io_pipe_phv_out_data_120; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_121 = pipe8_io_pipe_phv_out_data_121; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_122 = pipe8_io_pipe_phv_out_data_122; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_123 = pipe8_io_pipe_phv_out_data_123; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_124 = pipe8_io_pipe_phv_out_data_124; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_125 = pipe8_io_pipe_phv_out_data_125; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_126 = pipe8_io_pipe_phv_out_data_126; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_127 = pipe8_io_pipe_phv_out_data_127; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_128 = pipe8_io_pipe_phv_out_data_128; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_129 = pipe8_io_pipe_phv_out_data_129; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_130 = pipe8_io_pipe_phv_out_data_130; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_131 = pipe8_io_pipe_phv_out_data_131; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_132 = pipe8_io_pipe_phv_out_data_132; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_133 = pipe8_io_pipe_phv_out_data_133; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_134 = pipe8_io_pipe_phv_out_data_134; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_135 = pipe8_io_pipe_phv_out_data_135; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_136 = pipe8_io_pipe_phv_out_data_136; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_137 = pipe8_io_pipe_phv_out_data_137; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_138 = pipe8_io_pipe_phv_out_data_138; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_139 = pipe8_io_pipe_phv_out_data_139; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_140 = pipe8_io_pipe_phv_out_data_140; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_141 = pipe8_io_pipe_phv_out_data_141; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_142 = pipe8_io_pipe_phv_out_data_142; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_143 = pipe8_io_pipe_phv_out_data_143; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_144 = pipe8_io_pipe_phv_out_data_144; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_145 = pipe8_io_pipe_phv_out_data_145; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_146 = pipe8_io_pipe_phv_out_data_146; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_147 = pipe8_io_pipe_phv_out_data_147; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_148 = pipe8_io_pipe_phv_out_data_148; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_149 = pipe8_io_pipe_phv_out_data_149; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_150 = pipe8_io_pipe_phv_out_data_150; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_151 = pipe8_io_pipe_phv_out_data_151; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_152 = pipe8_io_pipe_phv_out_data_152; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_153 = pipe8_io_pipe_phv_out_data_153; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_154 = pipe8_io_pipe_phv_out_data_154; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_155 = pipe8_io_pipe_phv_out_data_155; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_156 = pipe8_io_pipe_phv_out_data_156; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_157 = pipe8_io_pipe_phv_out_data_157; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_158 = pipe8_io_pipe_phv_out_data_158; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_159 = pipe8_io_pipe_phv_out_data_159; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_160 = pipe8_io_pipe_phv_out_data_160; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_161 = pipe8_io_pipe_phv_out_data_161; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_162 = pipe8_io_pipe_phv_out_data_162; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_163 = pipe8_io_pipe_phv_out_data_163; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_164 = pipe8_io_pipe_phv_out_data_164; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_165 = pipe8_io_pipe_phv_out_data_165; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_166 = pipe8_io_pipe_phv_out_data_166; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_167 = pipe8_io_pipe_phv_out_data_167; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_168 = pipe8_io_pipe_phv_out_data_168; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_169 = pipe8_io_pipe_phv_out_data_169; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_170 = pipe8_io_pipe_phv_out_data_170; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_171 = pipe8_io_pipe_phv_out_data_171; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_172 = pipe8_io_pipe_phv_out_data_172; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_173 = pipe8_io_pipe_phv_out_data_173; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_174 = pipe8_io_pipe_phv_out_data_174; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_175 = pipe8_io_pipe_phv_out_data_175; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_176 = pipe8_io_pipe_phv_out_data_176; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_177 = pipe8_io_pipe_phv_out_data_177; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_178 = pipe8_io_pipe_phv_out_data_178; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_179 = pipe8_io_pipe_phv_out_data_179; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_180 = pipe8_io_pipe_phv_out_data_180; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_181 = pipe8_io_pipe_phv_out_data_181; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_182 = pipe8_io_pipe_phv_out_data_182; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_183 = pipe8_io_pipe_phv_out_data_183; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_184 = pipe8_io_pipe_phv_out_data_184; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_185 = pipe8_io_pipe_phv_out_data_185; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_186 = pipe8_io_pipe_phv_out_data_186; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_187 = pipe8_io_pipe_phv_out_data_187; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_188 = pipe8_io_pipe_phv_out_data_188; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_189 = pipe8_io_pipe_phv_out_data_189; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_190 = pipe8_io_pipe_phv_out_data_190; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_191 = pipe8_io_pipe_phv_out_data_191; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_192 = pipe8_io_pipe_phv_out_data_192; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_193 = pipe8_io_pipe_phv_out_data_193; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_194 = pipe8_io_pipe_phv_out_data_194; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_195 = pipe8_io_pipe_phv_out_data_195; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_196 = pipe8_io_pipe_phv_out_data_196; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_197 = pipe8_io_pipe_phv_out_data_197; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_198 = pipe8_io_pipe_phv_out_data_198; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_199 = pipe8_io_pipe_phv_out_data_199; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_200 = pipe8_io_pipe_phv_out_data_200; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_201 = pipe8_io_pipe_phv_out_data_201; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_202 = pipe8_io_pipe_phv_out_data_202; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_203 = pipe8_io_pipe_phv_out_data_203; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_204 = pipe8_io_pipe_phv_out_data_204; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_205 = pipe8_io_pipe_phv_out_data_205; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_206 = pipe8_io_pipe_phv_out_data_206; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_207 = pipe8_io_pipe_phv_out_data_207; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_208 = pipe8_io_pipe_phv_out_data_208; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_209 = pipe8_io_pipe_phv_out_data_209; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_210 = pipe8_io_pipe_phv_out_data_210; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_211 = pipe8_io_pipe_phv_out_data_211; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_212 = pipe8_io_pipe_phv_out_data_212; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_213 = pipe8_io_pipe_phv_out_data_213; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_214 = pipe8_io_pipe_phv_out_data_214; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_215 = pipe8_io_pipe_phv_out_data_215; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_216 = pipe8_io_pipe_phv_out_data_216; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_217 = pipe8_io_pipe_phv_out_data_217; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_218 = pipe8_io_pipe_phv_out_data_218; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_219 = pipe8_io_pipe_phv_out_data_219; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_220 = pipe8_io_pipe_phv_out_data_220; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_221 = pipe8_io_pipe_phv_out_data_221; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_222 = pipe8_io_pipe_phv_out_data_222; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_223 = pipe8_io_pipe_phv_out_data_223; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_224 = pipe8_io_pipe_phv_out_data_224; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_225 = pipe8_io_pipe_phv_out_data_225; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_226 = pipe8_io_pipe_phv_out_data_226; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_227 = pipe8_io_pipe_phv_out_data_227; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_228 = pipe8_io_pipe_phv_out_data_228; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_229 = pipe8_io_pipe_phv_out_data_229; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_230 = pipe8_io_pipe_phv_out_data_230; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_231 = pipe8_io_pipe_phv_out_data_231; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_232 = pipe8_io_pipe_phv_out_data_232; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_233 = pipe8_io_pipe_phv_out_data_233; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_234 = pipe8_io_pipe_phv_out_data_234; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_235 = pipe8_io_pipe_phv_out_data_235; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_236 = pipe8_io_pipe_phv_out_data_236; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_237 = pipe8_io_pipe_phv_out_data_237; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_238 = pipe8_io_pipe_phv_out_data_238; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_239 = pipe8_io_pipe_phv_out_data_239; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_240 = pipe8_io_pipe_phv_out_data_240; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_241 = pipe8_io_pipe_phv_out_data_241; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_242 = pipe8_io_pipe_phv_out_data_242; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_243 = pipe8_io_pipe_phv_out_data_243; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_244 = pipe8_io_pipe_phv_out_data_244; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_245 = pipe8_io_pipe_phv_out_data_245; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_246 = pipe8_io_pipe_phv_out_data_246; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_247 = pipe8_io_pipe_phv_out_data_247; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_248 = pipe8_io_pipe_phv_out_data_248; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_249 = pipe8_io_pipe_phv_out_data_249; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_250 = pipe8_io_pipe_phv_out_data_250; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_251 = pipe8_io_pipe_phv_out_data_251; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_252 = pipe8_io_pipe_phv_out_data_252; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_253 = pipe8_io_pipe_phv_out_data_253; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_254 = pipe8_io_pipe_phv_out_data_254; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_255 = pipe8_io_pipe_phv_out_data_255; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_256 = pipe8_io_pipe_phv_out_data_256; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_257 = pipe8_io_pipe_phv_out_data_257; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_258 = pipe8_io_pipe_phv_out_data_258; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_259 = pipe8_io_pipe_phv_out_data_259; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_260 = pipe8_io_pipe_phv_out_data_260; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_261 = pipe8_io_pipe_phv_out_data_261; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_262 = pipe8_io_pipe_phv_out_data_262; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_263 = pipe8_io_pipe_phv_out_data_263; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_264 = pipe8_io_pipe_phv_out_data_264; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_265 = pipe8_io_pipe_phv_out_data_265; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_266 = pipe8_io_pipe_phv_out_data_266; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_267 = pipe8_io_pipe_phv_out_data_267; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_268 = pipe8_io_pipe_phv_out_data_268; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_269 = pipe8_io_pipe_phv_out_data_269; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_270 = pipe8_io_pipe_phv_out_data_270; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_271 = pipe8_io_pipe_phv_out_data_271; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_272 = pipe8_io_pipe_phv_out_data_272; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_273 = pipe8_io_pipe_phv_out_data_273; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_274 = pipe8_io_pipe_phv_out_data_274; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_275 = pipe8_io_pipe_phv_out_data_275; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_276 = pipe8_io_pipe_phv_out_data_276; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_277 = pipe8_io_pipe_phv_out_data_277; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_278 = pipe8_io_pipe_phv_out_data_278; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_279 = pipe8_io_pipe_phv_out_data_279; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_280 = pipe8_io_pipe_phv_out_data_280; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_281 = pipe8_io_pipe_phv_out_data_281; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_282 = pipe8_io_pipe_phv_out_data_282; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_283 = pipe8_io_pipe_phv_out_data_283; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_284 = pipe8_io_pipe_phv_out_data_284; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_285 = pipe8_io_pipe_phv_out_data_285; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_286 = pipe8_io_pipe_phv_out_data_286; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_287 = pipe8_io_pipe_phv_out_data_287; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_288 = pipe8_io_pipe_phv_out_data_288; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_289 = pipe8_io_pipe_phv_out_data_289; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_290 = pipe8_io_pipe_phv_out_data_290; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_291 = pipe8_io_pipe_phv_out_data_291; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_292 = pipe8_io_pipe_phv_out_data_292; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_293 = pipe8_io_pipe_phv_out_data_293; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_294 = pipe8_io_pipe_phv_out_data_294; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_295 = pipe8_io_pipe_phv_out_data_295; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_296 = pipe8_io_pipe_phv_out_data_296; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_297 = pipe8_io_pipe_phv_out_data_297; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_298 = pipe8_io_pipe_phv_out_data_298; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_299 = pipe8_io_pipe_phv_out_data_299; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_300 = pipe8_io_pipe_phv_out_data_300; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_301 = pipe8_io_pipe_phv_out_data_301; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_302 = pipe8_io_pipe_phv_out_data_302; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_303 = pipe8_io_pipe_phv_out_data_303; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_304 = pipe8_io_pipe_phv_out_data_304; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_305 = pipe8_io_pipe_phv_out_data_305; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_306 = pipe8_io_pipe_phv_out_data_306; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_307 = pipe8_io_pipe_phv_out_data_307; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_308 = pipe8_io_pipe_phv_out_data_308; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_309 = pipe8_io_pipe_phv_out_data_309; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_310 = pipe8_io_pipe_phv_out_data_310; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_311 = pipe8_io_pipe_phv_out_data_311; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_312 = pipe8_io_pipe_phv_out_data_312; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_313 = pipe8_io_pipe_phv_out_data_313; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_314 = pipe8_io_pipe_phv_out_data_314; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_315 = pipe8_io_pipe_phv_out_data_315; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_316 = pipe8_io_pipe_phv_out_data_316; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_317 = pipe8_io_pipe_phv_out_data_317; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_318 = pipe8_io_pipe_phv_out_data_318; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_319 = pipe8_io_pipe_phv_out_data_319; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_320 = pipe8_io_pipe_phv_out_data_320; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_321 = pipe8_io_pipe_phv_out_data_321; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_322 = pipe8_io_pipe_phv_out_data_322; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_323 = pipe8_io_pipe_phv_out_data_323; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_324 = pipe8_io_pipe_phv_out_data_324; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_325 = pipe8_io_pipe_phv_out_data_325; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_326 = pipe8_io_pipe_phv_out_data_326; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_327 = pipe8_io_pipe_phv_out_data_327; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_328 = pipe8_io_pipe_phv_out_data_328; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_329 = pipe8_io_pipe_phv_out_data_329; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_330 = pipe8_io_pipe_phv_out_data_330; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_331 = pipe8_io_pipe_phv_out_data_331; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_332 = pipe8_io_pipe_phv_out_data_332; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_333 = pipe8_io_pipe_phv_out_data_333; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_334 = pipe8_io_pipe_phv_out_data_334; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_335 = pipe8_io_pipe_phv_out_data_335; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_336 = pipe8_io_pipe_phv_out_data_336; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_337 = pipe8_io_pipe_phv_out_data_337; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_338 = pipe8_io_pipe_phv_out_data_338; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_339 = pipe8_io_pipe_phv_out_data_339; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_340 = pipe8_io_pipe_phv_out_data_340; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_341 = pipe8_io_pipe_phv_out_data_341; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_342 = pipe8_io_pipe_phv_out_data_342; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_343 = pipe8_io_pipe_phv_out_data_343; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_344 = pipe8_io_pipe_phv_out_data_344; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_345 = pipe8_io_pipe_phv_out_data_345; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_346 = pipe8_io_pipe_phv_out_data_346; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_347 = pipe8_io_pipe_phv_out_data_347; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_348 = pipe8_io_pipe_phv_out_data_348; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_349 = pipe8_io_pipe_phv_out_data_349; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_350 = pipe8_io_pipe_phv_out_data_350; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_351 = pipe8_io_pipe_phv_out_data_351; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_352 = pipe8_io_pipe_phv_out_data_352; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_353 = pipe8_io_pipe_phv_out_data_353; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_354 = pipe8_io_pipe_phv_out_data_354; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_355 = pipe8_io_pipe_phv_out_data_355; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_356 = pipe8_io_pipe_phv_out_data_356; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_357 = pipe8_io_pipe_phv_out_data_357; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_358 = pipe8_io_pipe_phv_out_data_358; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_359 = pipe8_io_pipe_phv_out_data_359; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_360 = pipe8_io_pipe_phv_out_data_360; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_361 = pipe8_io_pipe_phv_out_data_361; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_362 = pipe8_io_pipe_phv_out_data_362; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_363 = pipe8_io_pipe_phv_out_data_363; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_364 = pipe8_io_pipe_phv_out_data_364; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_365 = pipe8_io_pipe_phv_out_data_365; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_366 = pipe8_io_pipe_phv_out_data_366; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_367 = pipe8_io_pipe_phv_out_data_367; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_368 = pipe8_io_pipe_phv_out_data_368; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_369 = pipe8_io_pipe_phv_out_data_369; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_370 = pipe8_io_pipe_phv_out_data_370; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_371 = pipe8_io_pipe_phv_out_data_371; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_372 = pipe8_io_pipe_phv_out_data_372; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_373 = pipe8_io_pipe_phv_out_data_373; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_374 = pipe8_io_pipe_phv_out_data_374; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_375 = pipe8_io_pipe_phv_out_data_375; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_376 = pipe8_io_pipe_phv_out_data_376; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_377 = pipe8_io_pipe_phv_out_data_377; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_378 = pipe8_io_pipe_phv_out_data_378; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_379 = pipe8_io_pipe_phv_out_data_379; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_380 = pipe8_io_pipe_phv_out_data_380; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_381 = pipe8_io_pipe_phv_out_data_381; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_382 = pipe8_io_pipe_phv_out_data_382; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_383 = pipe8_io_pipe_phv_out_data_383; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_384 = pipe8_io_pipe_phv_out_data_384; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_385 = pipe8_io_pipe_phv_out_data_385; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_386 = pipe8_io_pipe_phv_out_data_386; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_387 = pipe8_io_pipe_phv_out_data_387; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_388 = pipe8_io_pipe_phv_out_data_388; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_389 = pipe8_io_pipe_phv_out_data_389; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_390 = pipe8_io_pipe_phv_out_data_390; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_391 = pipe8_io_pipe_phv_out_data_391; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_392 = pipe8_io_pipe_phv_out_data_392; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_393 = pipe8_io_pipe_phv_out_data_393; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_394 = pipe8_io_pipe_phv_out_data_394; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_395 = pipe8_io_pipe_phv_out_data_395; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_396 = pipe8_io_pipe_phv_out_data_396; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_397 = pipe8_io_pipe_phv_out_data_397; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_398 = pipe8_io_pipe_phv_out_data_398; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_399 = pipe8_io_pipe_phv_out_data_399; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_400 = pipe8_io_pipe_phv_out_data_400; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_401 = pipe8_io_pipe_phv_out_data_401; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_402 = pipe8_io_pipe_phv_out_data_402; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_403 = pipe8_io_pipe_phv_out_data_403; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_404 = pipe8_io_pipe_phv_out_data_404; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_405 = pipe8_io_pipe_phv_out_data_405; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_406 = pipe8_io_pipe_phv_out_data_406; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_407 = pipe8_io_pipe_phv_out_data_407; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_408 = pipe8_io_pipe_phv_out_data_408; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_409 = pipe8_io_pipe_phv_out_data_409; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_410 = pipe8_io_pipe_phv_out_data_410; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_411 = pipe8_io_pipe_phv_out_data_411; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_412 = pipe8_io_pipe_phv_out_data_412; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_413 = pipe8_io_pipe_phv_out_data_413; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_414 = pipe8_io_pipe_phv_out_data_414; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_415 = pipe8_io_pipe_phv_out_data_415; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_416 = pipe8_io_pipe_phv_out_data_416; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_417 = pipe8_io_pipe_phv_out_data_417; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_418 = pipe8_io_pipe_phv_out_data_418; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_419 = pipe8_io_pipe_phv_out_data_419; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_420 = pipe8_io_pipe_phv_out_data_420; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_421 = pipe8_io_pipe_phv_out_data_421; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_422 = pipe8_io_pipe_phv_out_data_422; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_423 = pipe8_io_pipe_phv_out_data_423; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_424 = pipe8_io_pipe_phv_out_data_424; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_425 = pipe8_io_pipe_phv_out_data_425; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_426 = pipe8_io_pipe_phv_out_data_426; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_427 = pipe8_io_pipe_phv_out_data_427; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_428 = pipe8_io_pipe_phv_out_data_428; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_429 = pipe8_io_pipe_phv_out_data_429; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_430 = pipe8_io_pipe_phv_out_data_430; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_431 = pipe8_io_pipe_phv_out_data_431; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_432 = pipe8_io_pipe_phv_out_data_432; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_433 = pipe8_io_pipe_phv_out_data_433; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_434 = pipe8_io_pipe_phv_out_data_434; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_435 = pipe8_io_pipe_phv_out_data_435; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_436 = pipe8_io_pipe_phv_out_data_436; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_437 = pipe8_io_pipe_phv_out_data_437; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_438 = pipe8_io_pipe_phv_out_data_438; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_439 = pipe8_io_pipe_phv_out_data_439; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_440 = pipe8_io_pipe_phv_out_data_440; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_441 = pipe8_io_pipe_phv_out_data_441; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_442 = pipe8_io_pipe_phv_out_data_442; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_443 = pipe8_io_pipe_phv_out_data_443; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_444 = pipe8_io_pipe_phv_out_data_444; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_445 = pipe8_io_pipe_phv_out_data_445; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_446 = pipe8_io_pipe_phv_out_data_446; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_447 = pipe8_io_pipe_phv_out_data_447; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_448 = pipe8_io_pipe_phv_out_data_448; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_449 = pipe8_io_pipe_phv_out_data_449; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_450 = pipe8_io_pipe_phv_out_data_450; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_451 = pipe8_io_pipe_phv_out_data_451; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_452 = pipe8_io_pipe_phv_out_data_452; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_453 = pipe8_io_pipe_phv_out_data_453; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_454 = pipe8_io_pipe_phv_out_data_454; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_455 = pipe8_io_pipe_phv_out_data_455; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_456 = pipe8_io_pipe_phv_out_data_456; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_457 = pipe8_io_pipe_phv_out_data_457; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_458 = pipe8_io_pipe_phv_out_data_458; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_459 = pipe8_io_pipe_phv_out_data_459; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_460 = pipe8_io_pipe_phv_out_data_460; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_461 = pipe8_io_pipe_phv_out_data_461; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_462 = pipe8_io_pipe_phv_out_data_462; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_463 = pipe8_io_pipe_phv_out_data_463; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_464 = pipe8_io_pipe_phv_out_data_464; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_465 = pipe8_io_pipe_phv_out_data_465; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_466 = pipe8_io_pipe_phv_out_data_466; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_467 = pipe8_io_pipe_phv_out_data_467; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_468 = pipe8_io_pipe_phv_out_data_468; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_469 = pipe8_io_pipe_phv_out_data_469; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_470 = pipe8_io_pipe_phv_out_data_470; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_471 = pipe8_io_pipe_phv_out_data_471; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_472 = pipe8_io_pipe_phv_out_data_472; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_473 = pipe8_io_pipe_phv_out_data_473; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_474 = pipe8_io_pipe_phv_out_data_474; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_475 = pipe8_io_pipe_phv_out_data_475; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_476 = pipe8_io_pipe_phv_out_data_476; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_477 = pipe8_io_pipe_phv_out_data_477; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_478 = pipe8_io_pipe_phv_out_data_478; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_479 = pipe8_io_pipe_phv_out_data_479; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_480 = pipe8_io_pipe_phv_out_data_480; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_481 = pipe8_io_pipe_phv_out_data_481; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_482 = pipe8_io_pipe_phv_out_data_482; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_483 = pipe8_io_pipe_phv_out_data_483; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_484 = pipe8_io_pipe_phv_out_data_484; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_485 = pipe8_io_pipe_phv_out_data_485; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_486 = pipe8_io_pipe_phv_out_data_486; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_487 = pipe8_io_pipe_phv_out_data_487; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_488 = pipe8_io_pipe_phv_out_data_488; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_489 = pipe8_io_pipe_phv_out_data_489; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_490 = pipe8_io_pipe_phv_out_data_490; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_491 = pipe8_io_pipe_phv_out_data_491; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_492 = pipe8_io_pipe_phv_out_data_492; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_493 = pipe8_io_pipe_phv_out_data_493; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_494 = pipe8_io_pipe_phv_out_data_494; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_495 = pipe8_io_pipe_phv_out_data_495; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_496 = pipe8_io_pipe_phv_out_data_496; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_497 = pipe8_io_pipe_phv_out_data_497; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_498 = pipe8_io_pipe_phv_out_data_498; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_499 = pipe8_io_pipe_phv_out_data_499; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_500 = pipe8_io_pipe_phv_out_data_500; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_501 = pipe8_io_pipe_phv_out_data_501; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_502 = pipe8_io_pipe_phv_out_data_502; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_503 = pipe8_io_pipe_phv_out_data_503; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_504 = pipe8_io_pipe_phv_out_data_504; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_505 = pipe8_io_pipe_phv_out_data_505; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_506 = pipe8_io_pipe_phv_out_data_506; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_507 = pipe8_io_pipe_phv_out_data_507; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_508 = pipe8_io_pipe_phv_out_data_508; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_509 = pipe8_io_pipe_phv_out_data_509; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_510 = pipe8_io_pipe_phv_out_data_510; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_511 = pipe8_io_pipe_phv_out_data_511; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_0 = pipe8_io_pipe_phv_out_header_0; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_1 = pipe8_io_pipe_phv_out_header_1; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_2 = pipe8_io_pipe_phv_out_header_2; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_3 = pipe8_io_pipe_phv_out_header_3; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_4 = pipe8_io_pipe_phv_out_header_4; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_5 = pipe8_io_pipe_phv_out_header_5; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_6 = pipe8_io_pipe_phv_out_header_6; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_7 = pipe8_io_pipe_phv_out_header_7; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_8 = pipe8_io_pipe_phv_out_header_8; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_9 = pipe8_io_pipe_phv_out_header_9; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_10 = pipe8_io_pipe_phv_out_header_10; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_11 = pipe8_io_pipe_phv_out_header_11; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_12 = pipe8_io_pipe_phv_out_header_12; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_13 = pipe8_io_pipe_phv_out_header_13; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_14 = pipe8_io_pipe_phv_out_header_14; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_15 = pipe8_io_pipe_phv_out_header_15; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_current_state = pipe8_io_pipe_phv_out_parse_current_state; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_current_offset = pipe8_io_pipe_phv_out_parse_current_offset; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_transition_field = pipe8_io_pipe_phv_out_parse_transition_field; // @[hash.scala 176:27]
  assign io_pipe_phv_out_next_processor_id = pipe8_io_pipe_phv_out_next_processor_id; // @[hash.scala 176:27]
  assign io_pipe_phv_out_next_config_id = pipe8_io_pipe_phv_out_next_config_id; // @[hash.scala 176:27]
  assign io_pipe_phv_out_is_valid_processor = pipe8_io_pipe_phv_out_is_valid_processor; // @[hash.scala 176:27]
  assign io_key_out = pipe8_io_key_out; // @[hash.scala 177:27]
  assign io_hash_val = pipe8_io_sum_out[7:0]; // @[hash.scala 178:46]
  assign io_hash_val_cs = pipe8_io_val_out[15:12]; // @[hash.scala 179:46]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_256 = io_pipe_phv_in_data_256; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_257 = io_pipe_phv_in_data_257; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_258 = io_pipe_phv_in_data_258; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_259 = io_pipe_phv_in_data_259; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_260 = io_pipe_phv_in_data_260; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_261 = io_pipe_phv_in_data_261; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_262 = io_pipe_phv_in_data_262; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_263 = io_pipe_phv_in_data_263; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_264 = io_pipe_phv_in_data_264; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_265 = io_pipe_phv_in_data_265; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_266 = io_pipe_phv_in_data_266; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_267 = io_pipe_phv_in_data_267; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_268 = io_pipe_phv_in_data_268; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_269 = io_pipe_phv_in_data_269; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_270 = io_pipe_phv_in_data_270; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_271 = io_pipe_phv_in_data_271; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_272 = io_pipe_phv_in_data_272; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_273 = io_pipe_phv_in_data_273; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_274 = io_pipe_phv_in_data_274; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_275 = io_pipe_phv_in_data_275; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_276 = io_pipe_phv_in_data_276; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_277 = io_pipe_phv_in_data_277; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_278 = io_pipe_phv_in_data_278; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_279 = io_pipe_phv_in_data_279; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_280 = io_pipe_phv_in_data_280; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_281 = io_pipe_phv_in_data_281; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_282 = io_pipe_phv_in_data_282; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_283 = io_pipe_phv_in_data_283; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_284 = io_pipe_phv_in_data_284; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_285 = io_pipe_phv_in_data_285; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_286 = io_pipe_phv_in_data_286; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_287 = io_pipe_phv_in_data_287; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_288 = io_pipe_phv_in_data_288; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_289 = io_pipe_phv_in_data_289; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_290 = io_pipe_phv_in_data_290; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_291 = io_pipe_phv_in_data_291; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_292 = io_pipe_phv_in_data_292; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_293 = io_pipe_phv_in_data_293; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_294 = io_pipe_phv_in_data_294; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_295 = io_pipe_phv_in_data_295; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_296 = io_pipe_phv_in_data_296; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_297 = io_pipe_phv_in_data_297; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_298 = io_pipe_phv_in_data_298; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_299 = io_pipe_phv_in_data_299; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_300 = io_pipe_phv_in_data_300; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_301 = io_pipe_phv_in_data_301; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_302 = io_pipe_phv_in_data_302; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_303 = io_pipe_phv_in_data_303; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_304 = io_pipe_phv_in_data_304; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_305 = io_pipe_phv_in_data_305; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_306 = io_pipe_phv_in_data_306; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_307 = io_pipe_phv_in_data_307; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_308 = io_pipe_phv_in_data_308; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_309 = io_pipe_phv_in_data_309; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_310 = io_pipe_phv_in_data_310; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_311 = io_pipe_phv_in_data_311; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_312 = io_pipe_phv_in_data_312; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_313 = io_pipe_phv_in_data_313; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_314 = io_pipe_phv_in_data_314; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_315 = io_pipe_phv_in_data_315; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_316 = io_pipe_phv_in_data_316; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_317 = io_pipe_phv_in_data_317; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_318 = io_pipe_phv_in_data_318; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_319 = io_pipe_phv_in_data_319; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_320 = io_pipe_phv_in_data_320; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_321 = io_pipe_phv_in_data_321; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_322 = io_pipe_phv_in_data_322; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_323 = io_pipe_phv_in_data_323; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_324 = io_pipe_phv_in_data_324; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_325 = io_pipe_phv_in_data_325; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_326 = io_pipe_phv_in_data_326; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_327 = io_pipe_phv_in_data_327; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_328 = io_pipe_phv_in_data_328; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_329 = io_pipe_phv_in_data_329; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_330 = io_pipe_phv_in_data_330; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_331 = io_pipe_phv_in_data_331; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_332 = io_pipe_phv_in_data_332; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_333 = io_pipe_phv_in_data_333; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_334 = io_pipe_phv_in_data_334; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_335 = io_pipe_phv_in_data_335; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_336 = io_pipe_phv_in_data_336; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_337 = io_pipe_phv_in_data_337; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_338 = io_pipe_phv_in_data_338; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_339 = io_pipe_phv_in_data_339; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_340 = io_pipe_phv_in_data_340; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_341 = io_pipe_phv_in_data_341; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_342 = io_pipe_phv_in_data_342; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_343 = io_pipe_phv_in_data_343; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_344 = io_pipe_phv_in_data_344; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_345 = io_pipe_phv_in_data_345; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_346 = io_pipe_phv_in_data_346; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_347 = io_pipe_phv_in_data_347; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_348 = io_pipe_phv_in_data_348; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_349 = io_pipe_phv_in_data_349; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_350 = io_pipe_phv_in_data_350; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_351 = io_pipe_phv_in_data_351; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_352 = io_pipe_phv_in_data_352; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_353 = io_pipe_phv_in_data_353; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_354 = io_pipe_phv_in_data_354; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_355 = io_pipe_phv_in_data_355; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_356 = io_pipe_phv_in_data_356; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_357 = io_pipe_phv_in_data_357; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_358 = io_pipe_phv_in_data_358; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_359 = io_pipe_phv_in_data_359; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_360 = io_pipe_phv_in_data_360; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_361 = io_pipe_phv_in_data_361; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_362 = io_pipe_phv_in_data_362; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_363 = io_pipe_phv_in_data_363; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_364 = io_pipe_phv_in_data_364; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_365 = io_pipe_phv_in_data_365; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_366 = io_pipe_phv_in_data_366; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_367 = io_pipe_phv_in_data_367; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_368 = io_pipe_phv_in_data_368; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_369 = io_pipe_phv_in_data_369; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_370 = io_pipe_phv_in_data_370; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_371 = io_pipe_phv_in_data_371; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_372 = io_pipe_phv_in_data_372; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_373 = io_pipe_phv_in_data_373; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_374 = io_pipe_phv_in_data_374; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_375 = io_pipe_phv_in_data_375; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_376 = io_pipe_phv_in_data_376; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_377 = io_pipe_phv_in_data_377; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_378 = io_pipe_phv_in_data_378; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_379 = io_pipe_phv_in_data_379; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_380 = io_pipe_phv_in_data_380; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_381 = io_pipe_phv_in_data_381; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_382 = io_pipe_phv_in_data_382; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_383 = io_pipe_phv_in_data_383; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_384 = io_pipe_phv_in_data_384; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_385 = io_pipe_phv_in_data_385; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_386 = io_pipe_phv_in_data_386; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_387 = io_pipe_phv_in_data_387; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_388 = io_pipe_phv_in_data_388; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_389 = io_pipe_phv_in_data_389; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_390 = io_pipe_phv_in_data_390; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_391 = io_pipe_phv_in_data_391; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_392 = io_pipe_phv_in_data_392; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_393 = io_pipe_phv_in_data_393; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_394 = io_pipe_phv_in_data_394; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_395 = io_pipe_phv_in_data_395; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_396 = io_pipe_phv_in_data_396; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_397 = io_pipe_phv_in_data_397; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_398 = io_pipe_phv_in_data_398; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_399 = io_pipe_phv_in_data_399; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_400 = io_pipe_phv_in_data_400; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_401 = io_pipe_phv_in_data_401; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_402 = io_pipe_phv_in_data_402; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_403 = io_pipe_phv_in_data_403; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_404 = io_pipe_phv_in_data_404; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_405 = io_pipe_phv_in_data_405; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_406 = io_pipe_phv_in_data_406; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_407 = io_pipe_phv_in_data_407; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_408 = io_pipe_phv_in_data_408; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_409 = io_pipe_phv_in_data_409; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_410 = io_pipe_phv_in_data_410; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_411 = io_pipe_phv_in_data_411; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_412 = io_pipe_phv_in_data_412; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_413 = io_pipe_phv_in_data_413; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_414 = io_pipe_phv_in_data_414; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_415 = io_pipe_phv_in_data_415; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_416 = io_pipe_phv_in_data_416; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_417 = io_pipe_phv_in_data_417; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_418 = io_pipe_phv_in_data_418; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_419 = io_pipe_phv_in_data_419; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_420 = io_pipe_phv_in_data_420; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_421 = io_pipe_phv_in_data_421; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_422 = io_pipe_phv_in_data_422; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_423 = io_pipe_phv_in_data_423; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_424 = io_pipe_phv_in_data_424; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_425 = io_pipe_phv_in_data_425; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_426 = io_pipe_phv_in_data_426; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_427 = io_pipe_phv_in_data_427; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_428 = io_pipe_phv_in_data_428; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_429 = io_pipe_phv_in_data_429; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_430 = io_pipe_phv_in_data_430; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_431 = io_pipe_phv_in_data_431; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_432 = io_pipe_phv_in_data_432; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_433 = io_pipe_phv_in_data_433; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_434 = io_pipe_phv_in_data_434; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_435 = io_pipe_phv_in_data_435; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_436 = io_pipe_phv_in_data_436; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_437 = io_pipe_phv_in_data_437; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_438 = io_pipe_phv_in_data_438; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_439 = io_pipe_phv_in_data_439; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_440 = io_pipe_phv_in_data_440; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_441 = io_pipe_phv_in_data_441; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_442 = io_pipe_phv_in_data_442; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_443 = io_pipe_phv_in_data_443; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_444 = io_pipe_phv_in_data_444; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_445 = io_pipe_phv_in_data_445; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_446 = io_pipe_phv_in_data_446; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_447 = io_pipe_phv_in_data_447; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_448 = io_pipe_phv_in_data_448; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_449 = io_pipe_phv_in_data_449; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_450 = io_pipe_phv_in_data_450; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_451 = io_pipe_phv_in_data_451; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_452 = io_pipe_phv_in_data_452; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_453 = io_pipe_phv_in_data_453; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_454 = io_pipe_phv_in_data_454; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_455 = io_pipe_phv_in_data_455; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_456 = io_pipe_phv_in_data_456; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_457 = io_pipe_phv_in_data_457; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_458 = io_pipe_phv_in_data_458; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_459 = io_pipe_phv_in_data_459; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_460 = io_pipe_phv_in_data_460; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_461 = io_pipe_phv_in_data_461; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_462 = io_pipe_phv_in_data_462; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_463 = io_pipe_phv_in_data_463; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_464 = io_pipe_phv_in_data_464; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_465 = io_pipe_phv_in_data_465; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_466 = io_pipe_phv_in_data_466; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_467 = io_pipe_phv_in_data_467; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_468 = io_pipe_phv_in_data_468; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_469 = io_pipe_phv_in_data_469; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_470 = io_pipe_phv_in_data_470; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_471 = io_pipe_phv_in_data_471; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_472 = io_pipe_phv_in_data_472; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_473 = io_pipe_phv_in_data_473; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_474 = io_pipe_phv_in_data_474; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_475 = io_pipe_phv_in_data_475; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_476 = io_pipe_phv_in_data_476; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_477 = io_pipe_phv_in_data_477; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_478 = io_pipe_phv_in_data_478; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_479 = io_pipe_phv_in_data_479; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_480 = io_pipe_phv_in_data_480; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_481 = io_pipe_phv_in_data_481; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_482 = io_pipe_phv_in_data_482; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_483 = io_pipe_phv_in_data_483; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_484 = io_pipe_phv_in_data_484; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_485 = io_pipe_phv_in_data_485; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_486 = io_pipe_phv_in_data_486; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_487 = io_pipe_phv_in_data_487; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_488 = io_pipe_phv_in_data_488; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_489 = io_pipe_phv_in_data_489; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_490 = io_pipe_phv_in_data_490; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_491 = io_pipe_phv_in_data_491; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_492 = io_pipe_phv_in_data_492; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_493 = io_pipe_phv_in_data_493; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_494 = io_pipe_phv_in_data_494; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_495 = io_pipe_phv_in_data_495; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_496 = io_pipe_phv_in_data_496; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_497 = io_pipe_phv_in_data_497; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_498 = io_pipe_phv_in_data_498; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_499 = io_pipe_phv_in_data_499; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_500 = io_pipe_phv_in_data_500; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_501 = io_pipe_phv_in_data_501; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_502 = io_pipe_phv_in_data_502; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_503 = io_pipe_phv_in_data_503; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_504 = io_pipe_phv_in_data_504; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_505 = io_pipe_phv_in_data_505; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_506 = io_pipe_phv_in_data_506; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_507 = io_pipe_phv_in_data_507; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_508 = io_pipe_phv_in_data_508; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_509 = io_pipe_phv_in_data_509; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_510 = io_pipe_phv_in_data_510; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_511 = io_pipe_phv_in_data_511; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[hash.scala 136:27]
  assign pipe1_io_key_in = io_key_in; // @[hash.scala 137:27]
  assign pipe1_io_sum_in = pipe1_io_key_in; // @[hash.scala 138:27]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_256 = pipe1_io_pipe_phv_out_data_256; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_257 = pipe1_io_pipe_phv_out_data_257; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_258 = pipe1_io_pipe_phv_out_data_258; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_259 = pipe1_io_pipe_phv_out_data_259; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_260 = pipe1_io_pipe_phv_out_data_260; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_261 = pipe1_io_pipe_phv_out_data_261; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_262 = pipe1_io_pipe_phv_out_data_262; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_263 = pipe1_io_pipe_phv_out_data_263; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_264 = pipe1_io_pipe_phv_out_data_264; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_265 = pipe1_io_pipe_phv_out_data_265; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_266 = pipe1_io_pipe_phv_out_data_266; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_267 = pipe1_io_pipe_phv_out_data_267; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_268 = pipe1_io_pipe_phv_out_data_268; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_269 = pipe1_io_pipe_phv_out_data_269; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_270 = pipe1_io_pipe_phv_out_data_270; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_271 = pipe1_io_pipe_phv_out_data_271; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_272 = pipe1_io_pipe_phv_out_data_272; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_273 = pipe1_io_pipe_phv_out_data_273; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_274 = pipe1_io_pipe_phv_out_data_274; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_275 = pipe1_io_pipe_phv_out_data_275; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_276 = pipe1_io_pipe_phv_out_data_276; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_277 = pipe1_io_pipe_phv_out_data_277; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_278 = pipe1_io_pipe_phv_out_data_278; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_279 = pipe1_io_pipe_phv_out_data_279; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_280 = pipe1_io_pipe_phv_out_data_280; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_281 = pipe1_io_pipe_phv_out_data_281; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_282 = pipe1_io_pipe_phv_out_data_282; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_283 = pipe1_io_pipe_phv_out_data_283; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_284 = pipe1_io_pipe_phv_out_data_284; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_285 = pipe1_io_pipe_phv_out_data_285; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_286 = pipe1_io_pipe_phv_out_data_286; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_287 = pipe1_io_pipe_phv_out_data_287; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_288 = pipe1_io_pipe_phv_out_data_288; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_289 = pipe1_io_pipe_phv_out_data_289; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_290 = pipe1_io_pipe_phv_out_data_290; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_291 = pipe1_io_pipe_phv_out_data_291; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_292 = pipe1_io_pipe_phv_out_data_292; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_293 = pipe1_io_pipe_phv_out_data_293; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_294 = pipe1_io_pipe_phv_out_data_294; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_295 = pipe1_io_pipe_phv_out_data_295; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_296 = pipe1_io_pipe_phv_out_data_296; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_297 = pipe1_io_pipe_phv_out_data_297; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_298 = pipe1_io_pipe_phv_out_data_298; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_299 = pipe1_io_pipe_phv_out_data_299; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_300 = pipe1_io_pipe_phv_out_data_300; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_301 = pipe1_io_pipe_phv_out_data_301; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_302 = pipe1_io_pipe_phv_out_data_302; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_303 = pipe1_io_pipe_phv_out_data_303; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_304 = pipe1_io_pipe_phv_out_data_304; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_305 = pipe1_io_pipe_phv_out_data_305; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_306 = pipe1_io_pipe_phv_out_data_306; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_307 = pipe1_io_pipe_phv_out_data_307; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_308 = pipe1_io_pipe_phv_out_data_308; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_309 = pipe1_io_pipe_phv_out_data_309; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_310 = pipe1_io_pipe_phv_out_data_310; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_311 = pipe1_io_pipe_phv_out_data_311; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_312 = pipe1_io_pipe_phv_out_data_312; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_313 = pipe1_io_pipe_phv_out_data_313; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_314 = pipe1_io_pipe_phv_out_data_314; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_315 = pipe1_io_pipe_phv_out_data_315; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_316 = pipe1_io_pipe_phv_out_data_316; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_317 = pipe1_io_pipe_phv_out_data_317; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_318 = pipe1_io_pipe_phv_out_data_318; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_319 = pipe1_io_pipe_phv_out_data_319; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_320 = pipe1_io_pipe_phv_out_data_320; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_321 = pipe1_io_pipe_phv_out_data_321; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_322 = pipe1_io_pipe_phv_out_data_322; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_323 = pipe1_io_pipe_phv_out_data_323; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_324 = pipe1_io_pipe_phv_out_data_324; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_325 = pipe1_io_pipe_phv_out_data_325; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_326 = pipe1_io_pipe_phv_out_data_326; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_327 = pipe1_io_pipe_phv_out_data_327; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_328 = pipe1_io_pipe_phv_out_data_328; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_329 = pipe1_io_pipe_phv_out_data_329; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_330 = pipe1_io_pipe_phv_out_data_330; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_331 = pipe1_io_pipe_phv_out_data_331; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_332 = pipe1_io_pipe_phv_out_data_332; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_333 = pipe1_io_pipe_phv_out_data_333; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_334 = pipe1_io_pipe_phv_out_data_334; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_335 = pipe1_io_pipe_phv_out_data_335; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_336 = pipe1_io_pipe_phv_out_data_336; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_337 = pipe1_io_pipe_phv_out_data_337; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_338 = pipe1_io_pipe_phv_out_data_338; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_339 = pipe1_io_pipe_phv_out_data_339; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_340 = pipe1_io_pipe_phv_out_data_340; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_341 = pipe1_io_pipe_phv_out_data_341; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_342 = pipe1_io_pipe_phv_out_data_342; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_343 = pipe1_io_pipe_phv_out_data_343; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_344 = pipe1_io_pipe_phv_out_data_344; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_345 = pipe1_io_pipe_phv_out_data_345; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_346 = pipe1_io_pipe_phv_out_data_346; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_347 = pipe1_io_pipe_phv_out_data_347; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_348 = pipe1_io_pipe_phv_out_data_348; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_349 = pipe1_io_pipe_phv_out_data_349; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_350 = pipe1_io_pipe_phv_out_data_350; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_351 = pipe1_io_pipe_phv_out_data_351; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_352 = pipe1_io_pipe_phv_out_data_352; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_353 = pipe1_io_pipe_phv_out_data_353; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_354 = pipe1_io_pipe_phv_out_data_354; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_355 = pipe1_io_pipe_phv_out_data_355; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_356 = pipe1_io_pipe_phv_out_data_356; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_357 = pipe1_io_pipe_phv_out_data_357; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_358 = pipe1_io_pipe_phv_out_data_358; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_359 = pipe1_io_pipe_phv_out_data_359; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_360 = pipe1_io_pipe_phv_out_data_360; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_361 = pipe1_io_pipe_phv_out_data_361; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_362 = pipe1_io_pipe_phv_out_data_362; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_363 = pipe1_io_pipe_phv_out_data_363; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_364 = pipe1_io_pipe_phv_out_data_364; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_365 = pipe1_io_pipe_phv_out_data_365; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_366 = pipe1_io_pipe_phv_out_data_366; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_367 = pipe1_io_pipe_phv_out_data_367; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_368 = pipe1_io_pipe_phv_out_data_368; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_369 = pipe1_io_pipe_phv_out_data_369; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_370 = pipe1_io_pipe_phv_out_data_370; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_371 = pipe1_io_pipe_phv_out_data_371; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_372 = pipe1_io_pipe_phv_out_data_372; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_373 = pipe1_io_pipe_phv_out_data_373; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_374 = pipe1_io_pipe_phv_out_data_374; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_375 = pipe1_io_pipe_phv_out_data_375; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_376 = pipe1_io_pipe_phv_out_data_376; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_377 = pipe1_io_pipe_phv_out_data_377; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_378 = pipe1_io_pipe_phv_out_data_378; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_379 = pipe1_io_pipe_phv_out_data_379; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_380 = pipe1_io_pipe_phv_out_data_380; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_381 = pipe1_io_pipe_phv_out_data_381; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_382 = pipe1_io_pipe_phv_out_data_382; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_383 = pipe1_io_pipe_phv_out_data_383; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_384 = pipe1_io_pipe_phv_out_data_384; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_385 = pipe1_io_pipe_phv_out_data_385; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_386 = pipe1_io_pipe_phv_out_data_386; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_387 = pipe1_io_pipe_phv_out_data_387; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_388 = pipe1_io_pipe_phv_out_data_388; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_389 = pipe1_io_pipe_phv_out_data_389; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_390 = pipe1_io_pipe_phv_out_data_390; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_391 = pipe1_io_pipe_phv_out_data_391; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_392 = pipe1_io_pipe_phv_out_data_392; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_393 = pipe1_io_pipe_phv_out_data_393; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_394 = pipe1_io_pipe_phv_out_data_394; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_395 = pipe1_io_pipe_phv_out_data_395; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_396 = pipe1_io_pipe_phv_out_data_396; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_397 = pipe1_io_pipe_phv_out_data_397; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_398 = pipe1_io_pipe_phv_out_data_398; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_399 = pipe1_io_pipe_phv_out_data_399; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_400 = pipe1_io_pipe_phv_out_data_400; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_401 = pipe1_io_pipe_phv_out_data_401; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_402 = pipe1_io_pipe_phv_out_data_402; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_403 = pipe1_io_pipe_phv_out_data_403; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_404 = pipe1_io_pipe_phv_out_data_404; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_405 = pipe1_io_pipe_phv_out_data_405; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_406 = pipe1_io_pipe_phv_out_data_406; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_407 = pipe1_io_pipe_phv_out_data_407; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_408 = pipe1_io_pipe_phv_out_data_408; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_409 = pipe1_io_pipe_phv_out_data_409; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_410 = pipe1_io_pipe_phv_out_data_410; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_411 = pipe1_io_pipe_phv_out_data_411; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_412 = pipe1_io_pipe_phv_out_data_412; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_413 = pipe1_io_pipe_phv_out_data_413; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_414 = pipe1_io_pipe_phv_out_data_414; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_415 = pipe1_io_pipe_phv_out_data_415; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_416 = pipe1_io_pipe_phv_out_data_416; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_417 = pipe1_io_pipe_phv_out_data_417; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_418 = pipe1_io_pipe_phv_out_data_418; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_419 = pipe1_io_pipe_phv_out_data_419; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_420 = pipe1_io_pipe_phv_out_data_420; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_421 = pipe1_io_pipe_phv_out_data_421; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_422 = pipe1_io_pipe_phv_out_data_422; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_423 = pipe1_io_pipe_phv_out_data_423; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_424 = pipe1_io_pipe_phv_out_data_424; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_425 = pipe1_io_pipe_phv_out_data_425; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_426 = pipe1_io_pipe_phv_out_data_426; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_427 = pipe1_io_pipe_phv_out_data_427; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_428 = pipe1_io_pipe_phv_out_data_428; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_429 = pipe1_io_pipe_phv_out_data_429; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_430 = pipe1_io_pipe_phv_out_data_430; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_431 = pipe1_io_pipe_phv_out_data_431; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_432 = pipe1_io_pipe_phv_out_data_432; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_433 = pipe1_io_pipe_phv_out_data_433; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_434 = pipe1_io_pipe_phv_out_data_434; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_435 = pipe1_io_pipe_phv_out_data_435; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_436 = pipe1_io_pipe_phv_out_data_436; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_437 = pipe1_io_pipe_phv_out_data_437; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_438 = pipe1_io_pipe_phv_out_data_438; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_439 = pipe1_io_pipe_phv_out_data_439; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_440 = pipe1_io_pipe_phv_out_data_440; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_441 = pipe1_io_pipe_phv_out_data_441; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_442 = pipe1_io_pipe_phv_out_data_442; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_443 = pipe1_io_pipe_phv_out_data_443; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_444 = pipe1_io_pipe_phv_out_data_444; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_445 = pipe1_io_pipe_phv_out_data_445; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_446 = pipe1_io_pipe_phv_out_data_446; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_447 = pipe1_io_pipe_phv_out_data_447; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_448 = pipe1_io_pipe_phv_out_data_448; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_449 = pipe1_io_pipe_phv_out_data_449; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_450 = pipe1_io_pipe_phv_out_data_450; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_451 = pipe1_io_pipe_phv_out_data_451; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_452 = pipe1_io_pipe_phv_out_data_452; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_453 = pipe1_io_pipe_phv_out_data_453; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_454 = pipe1_io_pipe_phv_out_data_454; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_455 = pipe1_io_pipe_phv_out_data_455; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_456 = pipe1_io_pipe_phv_out_data_456; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_457 = pipe1_io_pipe_phv_out_data_457; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_458 = pipe1_io_pipe_phv_out_data_458; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_459 = pipe1_io_pipe_phv_out_data_459; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_460 = pipe1_io_pipe_phv_out_data_460; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_461 = pipe1_io_pipe_phv_out_data_461; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_462 = pipe1_io_pipe_phv_out_data_462; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_463 = pipe1_io_pipe_phv_out_data_463; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_464 = pipe1_io_pipe_phv_out_data_464; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_465 = pipe1_io_pipe_phv_out_data_465; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_466 = pipe1_io_pipe_phv_out_data_466; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_467 = pipe1_io_pipe_phv_out_data_467; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_468 = pipe1_io_pipe_phv_out_data_468; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_469 = pipe1_io_pipe_phv_out_data_469; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_470 = pipe1_io_pipe_phv_out_data_470; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_471 = pipe1_io_pipe_phv_out_data_471; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_472 = pipe1_io_pipe_phv_out_data_472; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_473 = pipe1_io_pipe_phv_out_data_473; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_474 = pipe1_io_pipe_phv_out_data_474; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_475 = pipe1_io_pipe_phv_out_data_475; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_476 = pipe1_io_pipe_phv_out_data_476; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_477 = pipe1_io_pipe_phv_out_data_477; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_478 = pipe1_io_pipe_phv_out_data_478; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_479 = pipe1_io_pipe_phv_out_data_479; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_480 = pipe1_io_pipe_phv_out_data_480; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_481 = pipe1_io_pipe_phv_out_data_481; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_482 = pipe1_io_pipe_phv_out_data_482; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_483 = pipe1_io_pipe_phv_out_data_483; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_484 = pipe1_io_pipe_phv_out_data_484; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_485 = pipe1_io_pipe_phv_out_data_485; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_486 = pipe1_io_pipe_phv_out_data_486; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_487 = pipe1_io_pipe_phv_out_data_487; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_488 = pipe1_io_pipe_phv_out_data_488; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_489 = pipe1_io_pipe_phv_out_data_489; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_490 = pipe1_io_pipe_phv_out_data_490; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_491 = pipe1_io_pipe_phv_out_data_491; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_492 = pipe1_io_pipe_phv_out_data_492; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_493 = pipe1_io_pipe_phv_out_data_493; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_494 = pipe1_io_pipe_phv_out_data_494; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_495 = pipe1_io_pipe_phv_out_data_495; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_496 = pipe1_io_pipe_phv_out_data_496; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_497 = pipe1_io_pipe_phv_out_data_497; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_498 = pipe1_io_pipe_phv_out_data_498; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_499 = pipe1_io_pipe_phv_out_data_499; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_500 = pipe1_io_pipe_phv_out_data_500; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_501 = pipe1_io_pipe_phv_out_data_501; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_502 = pipe1_io_pipe_phv_out_data_502; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_503 = pipe1_io_pipe_phv_out_data_503; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_504 = pipe1_io_pipe_phv_out_data_504; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_505 = pipe1_io_pipe_phv_out_data_505; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_506 = pipe1_io_pipe_phv_out_data_506; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_507 = pipe1_io_pipe_phv_out_data_507; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_508 = pipe1_io_pipe_phv_out_data_508; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_509 = pipe1_io_pipe_phv_out_data_509; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_510 = pipe1_io_pipe_phv_out_data_510; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_511 = pipe1_io_pipe_phv_out_data_511; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 140:27]
  assign pipe2_io_key_in = pipe1_io_key_out; // @[hash.scala 141:27]
  assign pipe2_io_sum_in = pipe1_io_sum_out; // @[hash.scala 142:27]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_256 = pipe2_io_pipe_phv_out_data_256; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_257 = pipe2_io_pipe_phv_out_data_257; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_258 = pipe2_io_pipe_phv_out_data_258; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_259 = pipe2_io_pipe_phv_out_data_259; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_260 = pipe2_io_pipe_phv_out_data_260; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_261 = pipe2_io_pipe_phv_out_data_261; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_262 = pipe2_io_pipe_phv_out_data_262; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_263 = pipe2_io_pipe_phv_out_data_263; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_264 = pipe2_io_pipe_phv_out_data_264; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_265 = pipe2_io_pipe_phv_out_data_265; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_266 = pipe2_io_pipe_phv_out_data_266; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_267 = pipe2_io_pipe_phv_out_data_267; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_268 = pipe2_io_pipe_phv_out_data_268; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_269 = pipe2_io_pipe_phv_out_data_269; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_270 = pipe2_io_pipe_phv_out_data_270; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_271 = pipe2_io_pipe_phv_out_data_271; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_272 = pipe2_io_pipe_phv_out_data_272; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_273 = pipe2_io_pipe_phv_out_data_273; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_274 = pipe2_io_pipe_phv_out_data_274; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_275 = pipe2_io_pipe_phv_out_data_275; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_276 = pipe2_io_pipe_phv_out_data_276; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_277 = pipe2_io_pipe_phv_out_data_277; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_278 = pipe2_io_pipe_phv_out_data_278; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_279 = pipe2_io_pipe_phv_out_data_279; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_280 = pipe2_io_pipe_phv_out_data_280; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_281 = pipe2_io_pipe_phv_out_data_281; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_282 = pipe2_io_pipe_phv_out_data_282; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_283 = pipe2_io_pipe_phv_out_data_283; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_284 = pipe2_io_pipe_phv_out_data_284; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_285 = pipe2_io_pipe_phv_out_data_285; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_286 = pipe2_io_pipe_phv_out_data_286; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_287 = pipe2_io_pipe_phv_out_data_287; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_288 = pipe2_io_pipe_phv_out_data_288; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_289 = pipe2_io_pipe_phv_out_data_289; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_290 = pipe2_io_pipe_phv_out_data_290; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_291 = pipe2_io_pipe_phv_out_data_291; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_292 = pipe2_io_pipe_phv_out_data_292; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_293 = pipe2_io_pipe_phv_out_data_293; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_294 = pipe2_io_pipe_phv_out_data_294; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_295 = pipe2_io_pipe_phv_out_data_295; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_296 = pipe2_io_pipe_phv_out_data_296; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_297 = pipe2_io_pipe_phv_out_data_297; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_298 = pipe2_io_pipe_phv_out_data_298; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_299 = pipe2_io_pipe_phv_out_data_299; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_300 = pipe2_io_pipe_phv_out_data_300; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_301 = pipe2_io_pipe_phv_out_data_301; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_302 = pipe2_io_pipe_phv_out_data_302; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_303 = pipe2_io_pipe_phv_out_data_303; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_304 = pipe2_io_pipe_phv_out_data_304; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_305 = pipe2_io_pipe_phv_out_data_305; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_306 = pipe2_io_pipe_phv_out_data_306; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_307 = pipe2_io_pipe_phv_out_data_307; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_308 = pipe2_io_pipe_phv_out_data_308; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_309 = pipe2_io_pipe_phv_out_data_309; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_310 = pipe2_io_pipe_phv_out_data_310; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_311 = pipe2_io_pipe_phv_out_data_311; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_312 = pipe2_io_pipe_phv_out_data_312; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_313 = pipe2_io_pipe_phv_out_data_313; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_314 = pipe2_io_pipe_phv_out_data_314; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_315 = pipe2_io_pipe_phv_out_data_315; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_316 = pipe2_io_pipe_phv_out_data_316; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_317 = pipe2_io_pipe_phv_out_data_317; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_318 = pipe2_io_pipe_phv_out_data_318; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_319 = pipe2_io_pipe_phv_out_data_319; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_320 = pipe2_io_pipe_phv_out_data_320; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_321 = pipe2_io_pipe_phv_out_data_321; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_322 = pipe2_io_pipe_phv_out_data_322; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_323 = pipe2_io_pipe_phv_out_data_323; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_324 = pipe2_io_pipe_phv_out_data_324; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_325 = pipe2_io_pipe_phv_out_data_325; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_326 = pipe2_io_pipe_phv_out_data_326; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_327 = pipe2_io_pipe_phv_out_data_327; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_328 = pipe2_io_pipe_phv_out_data_328; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_329 = pipe2_io_pipe_phv_out_data_329; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_330 = pipe2_io_pipe_phv_out_data_330; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_331 = pipe2_io_pipe_phv_out_data_331; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_332 = pipe2_io_pipe_phv_out_data_332; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_333 = pipe2_io_pipe_phv_out_data_333; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_334 = pipe2_io_pipe_phv_out_data_334; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_335 = pipe2_io_pipe_phv_out_data_335; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_336 = pipe2_io_pipe_phv_out_data_336; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_337 = pipe2_io_pipe_phv_out_data_337; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_338 = pipe2_io_pipe_phv_out_data_338; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_339 = pipe2_io_pipe_phv_out_data_339; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_340 = pipe2_io_pipe_phv_out_data_340; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_341 = pipe2_io_pipe_phv_out_data_341; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_342 = pipe2_io_pipe_phv_out_data_342; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_343 = pipe2_io_pipe_phv_out_data_343; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_344 = pipe2_io_pipe_phv_out_data_344; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_345 = pipe2_io_pipe_phv_out_data_345; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_346 = pipe2_io_pipe_phv_out_data_346; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_347 = pipe2_io_pipe_phv_out_data_347; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_348 = pipe2_io_pipe_phv_out_data_348; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_349 = pipe2_io_pipe_phv_out_data_349; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_350 = pipe2_io_pipe_phv_out_data_350; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_351 = pipe2_io_pipe_phv_out_data_351; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_352 = pipe2_io_pipe_phv_out_data_352; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_353 = pipe2_io_pipe_phv_out_data_353; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_354 = pipe2_io_pipe_phv_out_data_354; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_355 = pipe2_io_pipe_phv_out_data_355; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_356 = pipe2_io_pipe_phv_out_data_356; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_357 = pipe2_io_pipe_phv_out_data_357; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_358 = pipe2_io_pipe_phv_out_data_358; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_359 = pipe2_io_pipe_phv_out_data_359; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_360 = pipe2_io_pipe_phv_out_data_360; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_361 = pipe2_io_pipe_phv_out_data_361; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_362 = pipe2_io_pipe_phv_out_data_362; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_363 = pipe2_io_pipe_phv_out_data_363; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_364 = pipe2_io_pipe_phv_out_data_364; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_365 = pipe2_io_pipe_phv_out_data_365; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_366 = pipe2_io_pipe_phv_out_data_366; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_367 = pipe2_io_pipe_phv_out_data_367; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_368 = pipe2_io_pipe_phv_out_data_368; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_369 = pipe2_io_pipe_phv_out_data_369; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_370 = pipe2_io_pipe_phv_out_data_370; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_371 = pipe2_io_pipe_phv_out_data_371; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_372 = pipe2_io_pipe_phv_out_data_372; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_373 = pipe2_io_pipe_phv_out_data_373; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_374 = pipe2_io_pipe_phv_out_data_374; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_375 = pipe2_io_pipe_phv_out_data_375; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_376 = pipe2_io_pipe_phv_out_data_376; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_377 = pipe2_io_pipe_phv_out_data_377; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_378 = pipe2_io_pipe_phv_out_data_378; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_379 = pipe2_io_pipe_phv_out_data_379; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_380 = pipe2_io_pipe_phv_out_data_380; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_381 = pipe2_io_pipe_phv_out_data_381; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_382 = pipe2_io_pipe_phv_out_data_382; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_383 = pipe2_io_pipe_phv_out_data_383; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_384 = pipe2_io_pipe_phv_out_data_384; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_385 = pipe2_io_pipe_phv_out_data_385; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_386 = pipe2_io_pipe_phv_out_data_386; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_387 = pipe2_io_pipe_phv_out_data_387; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_388 = pipe2_io_pipe_phv_out_data_388; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_389 = pipe2_io_pipe_phv_out_data_389; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_390 = pipe2_io_pipe_phv_out_data_390; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_391 = pipe2_io_pipe_phv_out_data_391; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_392 = pipe2_io_pipe_phv_out_data_392; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_393 = pipe2_io_pipe_phv_out_data_393; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_394 = pipe2_io_pipe_phv_out_data_394; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_395 = pipe2_io_pipe_phv_out_data_395; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_396 = pipe2_io_pipe_phv_out_data_396; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_397 = pipe2_io_pipe_phv_out_data_397; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_398 = pipe2_io_pipe_phv_out_data_398; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_399 = pipe2_io_pipe_phv_out_data_399; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_400 = pipe2_io_pipe_phv_out_data_400; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_401 = pipe2_io_pipe_phv_out_data_401; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_402 = pipe2_io_pipe_phv_out_data_402; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_403 = pipe2_io_pipe_phv_out_data_403; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_404 = pipe2_io_pipe_phv_out_data_404; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_405 = pipe2_io_pipe_phv_out_data_405; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_406 = pipe2_io_pipe_phv_out_data_406; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_407 = pipe2_io_pipe_phv_out_data_407; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_408 = pipe2_io_pipe_phv_out_data_408; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_409 = pipe2_io_pipe_phv_out_data_409; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_410 = pipe2_io_pipe_phv_out_data_410; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_411 = pipe2_io_pipe_phv_out_data_411; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_412 = pipe2_io_pipe_phv_out_data_412; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_413 = pipe2_io_pipe_phv_out_data_413; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_414 = pipe2_io_pipe_phv_out_data_414; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_415 = pipe2_io_pipe_phv_out_data_415; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_416 = pipe2_io_pipe_phv_out_data_416; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_417 = pipe2_io_pipe_phv_out_data_417; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_418 = pipe2_io_pipe_phv_out_data_418; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_419 = pipe2_io_pipe_phv_out_data_419; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_420 = pipe2_io_pipe_phv_out_data_420; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_421 = pipe2_io_pipe_phv_out_data_421; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_422 = pipe2_io_pipe_phv_out_data_422; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_423 = pipe2_io_pipe_phv_out_data_423; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_424 = pipe2_io_pipe_phv_out_data_424; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_425 = pipe2_io_pipe_phv_out_data_425; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_426 = pipe2_io_pipe_phv_out_data_426; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_427 = pipe2_io_pipe_phv_out_data_427; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_428 = pipe2_io_pipe_phv_out_data_428; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_429 = pipe2_io_pipe_phv_out_data_429; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_430 = pipe2_io_pipe_phv_out_data_430; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_431 = pipe2_io_pipe_phv_out_data_431; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_432 = pipe2_io_pipe_phv_out_data_432; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_433 = pipe2_io_pipe_phv_out_data_433; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_434 = pipe2_io_pipe_phv_out_data_434; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_435 = pipe2_io_pipe_phv_out_data_435; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_436 = pipe2_io_pipe_phv_out_data_436; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_437 = pipe2_io_pipe_phv_out_data_437; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_438 = pipe2_io_pipe_phv_out_data_438; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_439 = pipe2_io_pipe_phv_out_data_439; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_440 = pipe2_io_pipe_phv_out_data_440; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_441 = pipe2_io_pipe_phv_out_data_441; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_442 = pipe2_io_pipe_phv_out_data_442; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_443 = pipe2_io_pipe_phv_out_data_443; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_444 = pipe2_io_pipe_phv_out_data_444; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_445 = pipe2_io_pipe_phv_out_data_445; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_446 = pipe2_io_pipe_phv_out_data_446; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_447 = pipe2_io_pipe_phv_out_data_447; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_448 = pipe2_io_pipe_phv_out_data_448; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_449 = pipe2_io_pipe_phv_out_data_449; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_450 = pipe2_io_pipe_phv_out_data_450; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_451 = pipe2_io_pipe_phv_out_data_451; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_452 = pipe2_io_pipe_phv_out_data_452; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_453 = pipe2_io_pipe_phv_out_data_453; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_454 = pipe2_io_pipe_phv_out_data_454; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_455 = pipe2_io_pipe_phv_out_data_455; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_456 = pipe2_io_pipe_phv_out_data_456; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_457 = pipe2_io_pipe_phv_out_data_457; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_458 = pipe2_io_pipe_phv_out_data_458; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_459 = pipe2_io_pipe_phv_out_data_459; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_460 = pipe2_io_pipe_phv_out_data_460; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_461 = pipe2_io_pipe_phv_out_data_461; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_462 = pipe2_io_pipe_phv_out_data_462; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_463 = pipe2_io_pipe_phv_out_data_463; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_464 = pipe2_io_pipe_phv_out_data_464; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_465 = pipe2_io_pipe_phv_out_data_465; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_466 = pipe2_io_pipe_phv_out_data_466; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_467 = pipe2_io_pipe_phv_out_data_467; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_468 = pipe2_io_pipe_phv_out_data_468; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_469 = pipe2_io_pipe_phv_out_data_469; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_470 = pipe2_io_pipe_phv_out_data_470; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_471 = pipe2_io_pipe_phv_out_data_471; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_472 = pipe2_io_pipe_phv_out_data_472; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_473 = pipe2_io_pipe_phv_out_data_473; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_474 = pipe2_io_pipe_phv_out_data_474; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_475 = pipe2_io_pipe_phv_out_data_475; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_476 = pipe2_io_pipe_phv_out_data_476; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_477 = pipe2_io_pipe_phv_out_data_477; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_478 = pipe2_io_pipe_phv_out_data_478; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_479 = pipe2_io_pipe_phv_out_data_479; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_480 = pipe2_io_pipe_phv_out_data_480; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_481 = pipe2_io_pipe_phv_out_data_481; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_482 = pipe2_io_pipe_phv_out_data_482; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_483 = pipe2_io_pipe_phv_out_data_483; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_484 = pipe2_io_pipe_phv_out_data_484; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_485 = pipe2_io_pipe_phv_out_data_485; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_486 = pipe2_io_pipe_phv_out_data_486; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_487 = pipe2_io_pipe_phv_out_data_487; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_488 = pipe2_io_pipe_phv_out_data_488; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_489 = pipe2_io_pipe_phv_out_data_489; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_490 = pipe2_io_pipe_phv_out_data_490; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_491 = pipe2_io_pipe_phv_out_data_491; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_492 = pipe2_io_pipe_phv_out_data_492; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_493 = pipe2_io_pipe_phv_out_data_493; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_494 = pipe2_io_pipe_phv_out_data_494; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_495 = pipe2_io_pipe_phv_out_data_495; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_496 = pipe2_io_pipe_phv_out_data_496; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_497 = pipe2_io_pipe_phv_out_data_497; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_498 = pipe2_io_pipe_phv_out_data_498; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_499 = pipe2_io_pipe_phv_out_data_499; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_500 = pipe2_io_pipe_phv_out_data_500; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_501 = pipe2_io_pipe_phv_out_data_501; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_502 = pipe2_io_pipe_phv_out_data_502; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_503 = pipe2_io_pipe_phv_out_data_503; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_504 = pipe2_io_pipe_phv_out_data_504; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_505 = pipe2_io_pipe_phv_out_data_505; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_506 = pipe2_io_pipe_phv_out_data_506; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_507 = pipe2_io_pipe_phv_out_data_507; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_508 = pipe2_io_pipe_phv_out_data_508; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_509 = pipe2_io_pipe_phv_out_data_509; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_510 = pipe2_io_pipe_phv_out_data_510; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_511 = pipe2_io_pipe_phv_out_data_511; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 144:27]
  assign pipe3_io_key_in = pipe2_io_key_out; // @[hash.scala 145:27]
  assign pipe3_io_sum_in = pipe2_io_sum_out; // @[hash.scala 146:27]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_160 = pipe3_io_pipe_phv_out_data_160; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_161 = pipe3_io_pipe_phv_out_data_161; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_162 = pipe3_io_pipe_phv_out_data_162; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_163 = pipe3_io_pipe_phv_out_data_163; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_164 = pipe3_io_pipe_phv_out_data_164; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_165 = pipe3_io_pipe_phv_out_data_165; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_166 = pipe3_io_pipe_phv_out_data_166; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_167 = pipe3_io_pipe_phv_out_data_167; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_168 = pipe3_io_pipe_phv_out_data_168; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_169 = pipe3_io_pipe_phv_out_data_169; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_170 = pipe3_io_pipe_phv_out_data_170; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_171 = pipe3_io_pipe_phv_out_data_171; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_172 = pipe3_io_pipe_phv_out_data_172; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_173 = pipe3_io_pipe_phv_out_data_173; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_174 = pipe3_io_pipe_phv_out_data_174; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_175 = pipe3_io_pipe_phv_out_data_175; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_176 = pipe3_io_pipe_phv_out_data_176; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_177 = pipe3_io_pipe_phv_out_data_177; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_178 = pipe3_io_pipe_phv_out_data_178; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_179 = pipe3_io_pipe_phv_out_data_179; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_180 = pipe3_io_pipe_phv_out_data_180; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_181 = pipe3_io_pipe_phv_out_data_181; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_182 = pipe3_io_pipe_phv_out_data_182; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_183 = pipe3_io_pipe_phv_out_data_183; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_184 = pipe3_io_pipe_phv_out_data_184; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_185 = pipe3_io_pipe_phv_out_data_185; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_186 = pipe3_io_pipe_phv_out_data_186; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_187 = pipe3_io_pipe_phv_out_data_187; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_188 = pipe3_io_pipe_phv_out_data_188; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_189 = pipe3_io_pipe_phv_out_data_189; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_190 = pipe3_io_pipe_phv_out_data_190; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_191 = pipe3_io_pipe_phv_out_data_191; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_192 = pipe3_io_pipe_phv_out_data_192; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_193 = pipe3_io_pipe_phv_out_data_193; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_194 = pipe3_io_pipe_phv_out_data_194; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_195 = pipe3_io_pipe_phv_out_data_195; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_196 = pipe3_io_pipe_phv_out_data_196; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_197 = pipe3_io_pipe_phv_out_data_197; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_198 = pipe3_io_pipe_phv_out_data_198; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_199 = pipe3_io_pipe_phv_out_data_199; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_200 = pipe3_io_pipe_phv_out_data_200; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_201 = pipe3_io_pipe_phv_out_data_201; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_202 = pipe3_io_pipe_phv_out_data_202; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_203 = pipe3_io_pipe_phv_out_data_203; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_204 = pipe3_io_pipe_phv_out_data_204; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_205 = pipe3_io_pipe_phv_out_data_205; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_206 = pipe3_io_pipe_phv_out_data_206; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_207 = pipe3_io_pipe_phv_out_data_207; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_208 = pipe3_io_pipe_phv_out_data_208; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_209 = pipe3_io_pipe_phv_out_data_209; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_210 = pipe3_io_pipe_phv_out_data_210; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_211 = pipe3_io_pipe_phv_out_data_211; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_212 = pipe3_io_pipe_phv_out_data_212; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_213 = pipe3_io_pipe_phv_out_data_213; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_214 = pipe3_io_pipe_phv_out_data_214; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_215 = pipe3_io_pipe_phv_out_data_215; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_216 = pipe3_io_pipe_phv_out_data_216; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_217 = pipe3_io_pipe_phv_out_data_217; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_218 = pipe3_io_pipe_phv_out_data_218; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_219 = pipe3_io_pipe_phv_out_data_219; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_220 = pipe3_io_pipe_phv_out_data_220; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_221 = pipe3_io_pipe_phv_out_data_221; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_222 = pipe3_io_pipe_phv_out_data_222; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_223 = pipe3_io_pipe_phv_out_data_223; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_224 = pipe3_io_pipe_phv_out_data_224; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_225 = pipe3_io_pipe_phv_out_data_225; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_226 = pipe3_io_pipe_phv_out_data_226; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_227 = pipe3_io_pipe_phv_out_data_227; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_228 = pipe3_io_pipe_phv_out_data_228; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_229 = pipe3_io_pipe_phv_out_data_229; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_230 = pipe3_io_pipe_phv_out_data_230; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_231 = pipe3_io_pipe_phv_out_data_231; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_232 = pipe3_io_pipe_phv_out_data_232; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_233 = pipe3_io_pipe_phv_out_data_233; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_234 = pipe3_io_pipe_phv_out_data_234; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_235 = pipe3_io_pipe_phv_out_data_235; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_236 = pipe3_io_pipe_phv_out_data_236; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_237 = pipe3_io_pipe_phv_out_data_237; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_238 = pipe3_io_pipe_phv_out_data_238; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_239 = pipe3_io_pipe_phv_out_data_239; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_240 = pipe3_io_pipe_phv_out_data_240; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_241 = pipe3_io_pipe_phv_out_data_241; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_242 = pipe3_io_pipe_phv_out_data_242; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_243 = pipe3_io_pipe_phv_out_data_243; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_244 = pipe3_io_pipe_phv_out_data_244; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_245 = pipe3_io_pipe_phv_out_data_245; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_246 = pipe3_io_pipe_phv_out_data_246; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_247 = pipe3_io_pipe_phv_out_data_247; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_248 = pipe3_io_pipe_phv_out_data_248; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_249 = pipe3_io_pipe_phv_out_data_249; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_250 = pipe3_io_pipe_phv_out_data_250; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_251 = pipe3_io_pipe_phv_out_data_251; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_252 = pipe3_io_pipe_phv_out_data_252; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_253 = pipe3_io_pipe_phv_out_data_253; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_254 = pipe3_io_pipe_phv_out_data_254; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_255 = pipe3_io_pipe_phv_out_data_255; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_256 = pipe3_io_pipe_phv_out_data_256; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_257 = pipe3_io_pipe_phv_out_data_257; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_258 = pipe3_io_pipe_phv_out_data_258; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_259 = pipe3_io_pipe_phv_out_data_259; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_260 = pipe3_io_pipe_phv_out_data_260; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_261 = pipe3_io_pipe_phv_out_data_261; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_262 = pipe3_io_pipe_phv_out_data_262; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_263 = pipe3_io_pipe_phv_out_data_263; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_264 = pipe3_io_pipe_phv_out_data_264; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_265 = pipe3_io_pipe_phv_out_data_265; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_266 = pipe3_io_pipe_phv_out_data_266; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_267 = pipe3_io_pipe_phv_out_data_267; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_268 = pipe3_io_pipe_phv_out_data_268; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_269 = pipe3_io_pipe_phv_out_data_269; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_270 = pipe3_io_pipe_phv_out_data_270; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_271 = pipe3_io_pipe_phv_out_data_271; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_272 = pipe3_io_pipe_phv_out_data_272; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_273 = pipe3_io_pipe_phv_out_data_273; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_274 = pipe3_io_pipe_phv_out_data_274; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_275 = pipe3_io_pipe_phv_out_data_275; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_276 = pipe3_io_pipe_phv_out_data_276; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_277 = pipe3_io_pipe_phv_out_data_277; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_278 = pipe3_io_pipe_phv_out_data_278; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_279 = pipe3_io_pipe_phv_out_data_279; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_280 = pipe3_io_pipe_phv_out_data_280; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_281 = pipe3_io_pipe_phv_out_data_281; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_282 = pipe3_io_pipe_phv_out_data_282; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_283 = pipe3_io_pipe_phv_out_data_283; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_284 = pipe3_io_pipe_phv_out_data_284; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_285 = pipe3_io_pipe_phv_out_data_285; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_286 = pipe3_io_pipe_phv_out_data_286; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_287 = pipe3_io_pipe_phv_out_data_287; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_288 = pipe3_io_pipe_phv_out_data_288; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_289 = pipe3_io_pipe_phv_out_data_289; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_290 = pipe3_io_pipe_phv_out_data_290; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_291 = pipe3_io_pipe_phv_out_data_291; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_292 = pipe3_io_pipe_phv_out_data_292; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_293 = pipe3_io_pipe_phv_out_data_293; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_294 = pipe3_io_pipe_phv_out_data_294; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_295 = pipe3_io_pipe_phv_out_data_295; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_296 = pipe3_io_pipe_phv_out_data_296; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_297 = pipe3_io_pipe_phv_out_data_297; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_298 = pipe3_io_pipe_phv_out_data_298; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_299 = pipe3_io_pipe_phv_out_data_299; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_300 = pipe3_io_pipe_phv_out_data_300; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_301 = pipe3_io_pipe_phv_out_data_301; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_302 = pipe3_io_pipe_phv_out_data_302; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_303 = pipe3_io_pipe_phv_out_data_303; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_304 = pipe3_io_pipe_phv_out_data_304; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_305 = pipe3_io_pipe_phv_out_data_305; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_306 = pipe3_io_pipe_phv_out_data_306; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_307 = pipe3_io_pipe_phv_out_data_307; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_308 = pipe3_io_pipe_phv_out_data_308; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_309 = pipe3_io_pipe_phv_out_data_309; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_310 = pipe3_io_pipe_phv_out_data_310; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_311 = pipe3_io_pipe_phv_out_data_311; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_312 = pipe3_io_pipe_phv_out_data_312; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_313 = pipe3_io_pipe_phv_out_data_313; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_314 = pipe3_io_pipe_phv_out_data_314; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_315 = pipe3_io_pipe_phv_out_data_315; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_316 = pipe3_io_pipe_phv_out_data_316; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_317 = pipe3_io_pipe_phv_out_data_317; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_318 = pipe3_io_pipe_phv_out_data_318; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_319 = pipe3_io_pipe_phv_out_data_319; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_320 = pipe3_io_pipe_phv_out_data_320; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_321 = pipe3_io_pipe_phv_out_data_321; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_322 = pipe3_io_pipe_phv_out_data_322; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_323 = pipe3_io_pipe_phv_out_data_323; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_324 = pipe3_io_pipe_phv_out_data_324; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_325 = pipe3_io_pipe_phv_out_data_325; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_326 = pipe3_io_pipe_phv_out_data_326; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_327 = pipe3_io_pipe_phv_out_data_327; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_328 = pipe3_io_pipe_phv_out_data_328; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_329 = pipe3_io_pipe_phv_out_data_329; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_330 = pipe3_io_pipe_phv_out_data_330; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_331 = pipe3_io_pipe_phv_out_data_331; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_332 = pipe3_io_pipe_phv_out_data_332; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_333 = pipe3_io_pipe_phv_out_data_333; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_334 = pipe3_io_pipe_phv_out_data_334; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_335 = pipe3_io_pipe_phv_out_data_335; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_336 = pipe3_io_pipe_phv_out_data_336; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_337 = pipe3_io_pipe_phv_out_data_337; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_338 = pipe3_io_pipe_phv_out_data_338; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_339 = pipe3_io_pipe_phv_out_data_339; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_340 = pipe3_io_pipe_phv_out_data_340; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_341 = pipe3_io_pipe_phv_out_data_341; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_342 = pipe3_io_pipe_phv_out_data_342; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_343 = pipe3_io_pipe_phv_out_data_343; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_344 = pipe3_io_pipe_phv_out_data_344; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_345 = pipe3_io_pipe_phv_out_data_345; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_346 = pipe3_io_pipe_phv_out_data_346; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_347 = pipe3_io_pipe_phv_out_data_347; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_348 = pipe3_io_pipe_phv_out_data_348; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_349 = pipe3_io_pipe_phv_out_data_349; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_350 = pipe3_io_pipe_phv_out_data_350; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_351 = pipe3_io_pipe_phv_out_data_351; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_352 = pipe3_io_pipe_phv_out_data_352; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_353 = pipe3_io_pipe_phv_out_data_353; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_354 = pipe3_io_pipe_phv_out_data_354; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_355 = pipe3_io_pipe_phv_out_data_355; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_356 = pipe3_io_pipe_phv_out_data_356; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_357 = pipe3_io_pipe_phv_out_data_357; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_358 = pipe3_io_pipe_phv_out_data_358; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_359 = pipe3_io_pipe_phv_out_data_359; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_360 = pipe3_io_pipe_phv_out_data_360; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_361 = pipe3_io_pipe_phv_out_data_361; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_362 = pipe3_io_pipe_phv_out_data_362; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_363 = pipe3_io_pipe_phv_out_data_363; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_364 = pipe3_io_pipe_phv_out_data_364; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_365 = pipe3_io_pipe_phv_out_data_365; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_366 = pipe3_io_pipe_phv_out_data_366; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_367 = pipe3_io_pipe_phv_out_data_367; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_368 = pipe3_io_pipe_phv_out_data_368; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_369 = pipe3_io_pipe_phv_out_data_369; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_370 = pipe3_io_pipe_phv_out_data_370; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_371 = pipe3_io_pipe_phv_out_data_371; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_372 = pipe3_io_pipe_phv_out_data_372; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_373 = pipe3_io_pipe_phv_out_data_373; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_374 = pipe3_io_pipe_phv_out_data_374; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_375 = pipe3_io_pipe_phv_out_data_375; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_376 = pipe3_io_pipe_phv_out_data_376; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_377 = pipe3_io_pipe_phv_out_data_377; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_378 = pipe3_io_pipe_phv_out_data_378; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_379 = pipe3_io_pipe_phv_out_data_379; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_380 = pipe3_io_pipe_phv_out_data_380; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_381 = pipe3_io_pipe_phv_out_data_381; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_382 = pipe3_io_pipe_phv_out_data_382; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_383 = pipe3_io_pipe_phv_out_data_383; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_384 = pipe3_io_pipe_phv_out_data_384; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_385 = pipe3_io_pipe_phv_out_data_385; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_386 = pipe3_io_pipe_phv_out_data_386; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_387 = pipe3_io_pipe_phv_out_data_387; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_388 = pipe3_io_pipe_phv_out_data_388; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_389 = pipe3_io_pipe_phv_out_data_389; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_390 = pipe3_io_pipe_phv_out_data_390; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_391 = pipe3_io_pipe_phv_out_data_391; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_392 = pipe3_io_pipe_phv_out_data_392; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_393 = pipe3_io_pipe_phv_out_data_393; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_394 = pipe3_io_pipe_phv_out_data_394; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_395 = pipe3_io_pipe_phv_out_data_395; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_396 = pipe3_io_pipe_phv_out_data_396; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_397 = pipe3_io_pipe_phv_out_data_397; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_398 = pipe3_io_pipe_phv_out_data_398; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_399 = pipe3_io_pipe_phv_out_data_399; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_400 = pipe3_io_pipe_phv_out_data_400; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_401 = pipe3_io_pipe_phv_out_data_401; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_402 = pipe3_io_pipe_phv_out_data_402; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_403 = pipe3_io_pipe_phv_out_data_403; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_404 = pipe3_io_pipe_phv_out_data_404; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_405 = pipe3_io_pipe_phv_out_data_405; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_406 = pipe3_io_pipe_phv_out_data_406; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_407 = pipe3_io_pipe_phv_out_data_407; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_408 = pipe3_io_pipe_phv_out_data_408; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_409 = pipe3_io_pipe_phv_out_data_409; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_410 = pipe3_io_pipe_phv_out_data_410; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_411 = pipe3_io_pipe_phv_out_data_411; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_412 = pipe3_io_pipe_phv_out_data_412; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_413 = pipe3_io_pipe_phv_out_data_413; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_414 = pipe3_io_pipe_phv_out_data_414; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_415 = pipe3_io_pipe_phv_out_data_415; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_416 = pipe3_io_pipe_phv_out_data_416; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_417 = pipe3_io_pipe_phv_out_data_417; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_418 = pipe3_io_pipe_phv_out_data_418; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_419 = pipe3_io_pipe_phv_out_data_419; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_420 = pipe3_io_pipe_phv_out_data_420; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_421 = pipe3_io_pipe_phv_out_data_421; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_422 = pipe3_io_pipe_phv_out_data_422; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_423 = pipe3_io_pipe_phv_out_data_423; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_424 = pipe3_io_pipe_phv_out_data_424; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_425 = pipe3_io_pipe_phv_out_data_425; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_426 = pipe3_io_pipe_phv_out_data_426; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_427 = pipe3_io_pipe_phv_out_data_427; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_428 = pipe3_io_pipe_phv_out_data_428; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_429 = pipe3_io_pipe_phv_out_data_429; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_430 = pipe3_io_pipe_phv_out_data_430; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_431 = pipe3_io_pipe_phv_out_data_431; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_432 = pipe3_io_pipe_phv_out_data_432; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_433 = pipe3_io_pipe_phv_out_data_433; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_434 = pipe3_io_pipe_phv_out_data_434; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_435 = pipe3_io_pipe_phv_out_data_435; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_436 = pipe3_io_pipe_phv_out_data_436; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_437 = pipe3_io_pipe_phv_out_data_437; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_438 = pipe3_io_pipe_phv_out_data_438; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_439 = pipe3_io_pipe_phv_out_data_439; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_440 = pipe3_io_pipe_phv_out_data_440; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_441 = pipe3_io_pipe_phv_out_data_441; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_442 = pipe3_io_pipe_phv_out_data_442; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_443 = pipe3_io_pipe_phv_out_data_443; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_444 = pipe3_io_pipe_phv_out_data_444; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_445 = pipe3_io_pipe_phv_out_data_445; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_446 = pipe3_io_pipe_phv_out_data_446; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_447 = pipe3_io_pipe_phv_out_data_447; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_448 = pipe3_io_pipe_phv_out_data_448; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_449 = pipe3_io_pipe_phv_out_data_449; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_450 = pipe3_io_pipe_phv_out_data_450; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_451 = pipe3_io_pipe_phv_out_data_451; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_452 = pipe3_io_pipe_phv_out_data_452; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_453 = pipe3_io_pipe_phv_out_data_453; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_454 = pipe3_io_pipe_phv_out_data_454; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_455 = pipe3_io_pipe_phv_out_data_455; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_456 = pipe3_io_pipe_phv_out_data_456; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_457 = pipe3_io_pipe_phv_out_data_457; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_458 = pipe3_io_pipe_phv_out_data_458; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_459 = pipe3_io_pipe_phv_out_data_459; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_460 = pipe3_io_pipe_phv_out_data_460; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_461 = pipe3_io_pipe_phv_out_data_461; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_462 = pipe3_io_pipe_phv_out_data_462; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_463 = pipe3_io_pipe_phv_out_data_463; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_464 = pipe3_io_pipe_phv_out_data_464; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_465 = pipe3_io_pipe_phv_out_data_465; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_466 = pipe3_io_pipe_phv_out_data_466; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_467 = pipe3_io_pipe_phv_out_data_467; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_468 = pipe3_io_pipe_phv_out_data_468; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_469 = pipe3_io_pipe_phv_out_data_469; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_470 = pipe3_io_pipe_phv_out_data_470; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_471 = pipe3_io_pipe_phv_out_data_471; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_472 = pipe3_io_pipe_phv_out_data_472; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_473 = pipe3_io_pipe_phv_out_data_473; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_474 = pipe3_io_pipe_phv_out_data_474; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_475 = pipe3_io_pipe_phv_out_data_475; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_476 = pipe3_io_pipe_phv_out_data_476; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_477 = pipe3_io_pipe_phv_out_data_477; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_478 = pipe3_io_pipe_phv_out_data_478; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_479 = pipe3_io_pipe_phv_out_data_479; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_480 = pipe3_io_pipe_phv_out_data_480; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_481 = pipe3_io_pipe_phv_out_data_481; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_482 = pipe3_io_pipe_phv_out_data_482; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_483 = pipe3_io_pipe_phv_out_data_483; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_484 = pipe3_io_pipe_phv_out_data_484; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_485 = pipe3_io_pipe_phv_out_data_485; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_486 = pipe3_io_pipe_phv_out_data_486; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_487 = pipe3_io_pipe_phv_out_data_487; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_488 = pipe3_io_pipe_phv_out_data_488; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_489 = pipe3_io_pipe_phv_out_data_489; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_490 = pipe3_io_pipe_phv_out_data_490; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_491 = pipe3_io_pipe_phv_out_data_491; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_492 = pipe3_io_pipe_phv_out_data_492; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_493 = pipe3_io_pipe_phv_out_data_493; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_494 = pipe3_io_pipe_phv_out_data_494; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_495 = pipe3_io_pipe_phv_out_data_495; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_496 = pipe3_io_pipe_phv_out_data_496; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_497 = pipe3_io_pipe_phv_out_data_497; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_498 = pipe3_io_pipe_phv_out_data_498; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_499 = pipe3_io_pipe_phv_out_data_499; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_500 = pipe3_io_pipe_phv_out_data_500; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_501 = pipe3_io_pipe_phv_out_data_501; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_502 = pipe3_io_pipe_phv_out_data_502; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_503 = pipe3_io_pipe_phv_out_data_503; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_504 = pipe3_io_pipe_phv_out_data_504; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_505 = pipe3_io_pipe_phv_out_data_505; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_506 = pipe3_io_pipe_phv_out_data_506; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_507 = pipe3_io_pipe_phv_out_data_507; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_508 = pipe3_io_pipe_phv_out_data_508; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_509 = pipe3_io_pipe_phv_out_data_509; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_510 = pipe3_io_pipe_phv_out_data_510; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_511 = pipe3_io_pipe_phv_out_data_511; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 148:27]
  assign pipe4_io_key_in = pipe3_io_key_out; // @[hash.scala 149:27]
  assign pipe4_io_sum_in = pipe3_io_sum_out; // @[hash.scala 150:27]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_96 = pipe4_io_pipe_phv_out_data_96; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_97 = pipe4_io_pipe_phv_out_data_97; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_98 = pipe4_io_pipe_phv_out_data_98; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_99 = pipe4_io_pipe_phv_out_data_99; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_100 = pipe4_io_pipe_phv_out_data_100; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_101 = pipe4_io_pipe_phv_out_data_101; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_102 = pipe4_io_pipe_phv_out_data_102; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_103 = pipe4_io_pipe_phv_out_data_103; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_104 = pipe4_io_pipe_phv_out_data_104; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_105 = pipe4_io_pipe_phv_out_data_105; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_106 = pipe4_io_pipe_phv_out_data_106; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_107 = pipe4_io_pipe_phv_out_data_107; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_108 = pipe4_io_pipe_phv_out_data_108; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_109 = pipe4_io_pipe_phv_out_data_109; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_110 = pipe4_io_pipe_phv_out_data_110; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_111 = pipe4_io_pipe_phv_out_data_111; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_112 = pipe4_io_pipe_phv_out_data_112; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_113 = pipe4_io_pipe_phv_out_data_113; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_114 = pipe4_io_pipe_phv_out_data_114; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_115 = pipe4_io_pipe_phv_out_data_115; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_116 = pipe4_io_pipe_phv_out_data_116; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_117 = pipe4_io_pipe_phv_out_data_117; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_118 = pipe4_io_pipe_phv_out_data_118; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_119 = pipe4_io_pipe_phv_out_data_119; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_120 = pipe4_io_pipe_phv_out_data_120; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_121 = pipe4_io_pipe_phv_out_data_121; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_122 = pipe4_io_pipe_phv_out_data_122; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_123 = pipe4_io_pipe_phv_out_data_123; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_124 = pipe4_io_pipe_phv_out_data_124; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_125 = pipe4_io_pipe_phv_out_data_125; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_126 = pipe4_io_pipe_phv_out_data_126; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_127 = pipe4_io_pipe_phv_out_data_127; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_128 = pipe4_io_pipe_phv_out_data_128; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_129 = pipe4_io_pipe_phv_out_data_129; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_130 = pipe4_io_pipe_phv_out_data_130; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_131 = pipe4_io_pipe_phv_out_data_131; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_132 = pipe4_io_pipe_phv_out_data_132; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_133 = pipe4_io_pipe_phv_out_data_133; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_134 = pipe4_io_pipe_phv_out_data_134; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_135 = pipe4_io_pipe_phv_out_data_135; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_136 = pipe4_io_pipe_phv_out_data_136; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_137 = pipe4_io_pipe_phv_out_data_137; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_138 = pipe4_io_pipe_phv_out_data_138; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_139 = pipe4_io_pipe_phv_out_data_139; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_140 = pipe4_io_pipe_phv_out_data_140; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_141 = pipe4_io_pipe_phv_out_data_141; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_142 = pipe4_io_pipe_phv_out_data_142; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_143 = pipe4_io_pipe_phv_out_data_143; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_144 = pipe4_io_pipe_phv_out_data_144; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_145 = pipe4_io_pipe_phv_out_data_145; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_146 = pipe4_io_pipe_phv_out_data_146; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_147 = pipe4_io_pipe_phv_out_data_147; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_148 = pipe4_io_pipe_phv_out_data_148; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_149 = pipe4_io_pipe_phv_out_data_149; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_150 = pipe4_io_pipe_phv_out_data_150; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_151 = pipe4_io_pipe_phv_out_data_151; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_152 = pipe4_io_pipe_phv_out_data_152; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_153 = pipe4_io_pipe_phv_out_data_153; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_154 = pipe4_io_pipe_phv_out_data_154; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_155 = pipe4_io_pipe_phv_out_data_155; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_156 = pipe4_io_pipe_phv_out_data_156; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_157 = pipe4_io_pipe_phv_out_data_157; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_158 = pipe4_io_pipe_phv_out_data_158; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_159 = pipe4_io_pipe_phv_out_data_159; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_160 = pipe4_io_pipe_phv_out_data_160; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_161 = pipe4_io_pipe_phv_out_data_161; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_162 = pipe4_io_pipe_phv_out_data_162; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_163 = pipe4_io_pipe_phv_out_data_163; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_164 = pipe4_io_pipe_phv_out_data_164; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_165 = pipe4_io_pipe_phv_out_data_165; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_166 = pipe4_io_pipe_phv_out_data_166; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_167 = pipe4_io_pipe_phv_out_data_167; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_168 = pipe4_io_pipe_phv_out_data_168; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_169 = pipe4_io_pipe_phv_out_data_169; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_170 = pipe4_io_pipe_phv_out_data_170; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_171 = pipe4_io_pipe_phv_out_data_171; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_172 = pipe4_io_pipe_phv_out_data_172; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_173 = pipe4_io_pipe_phv_out_data_173; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_174 = pipe4_io_pipe_phv_out_data_174; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_175 = pipe4_io_pipe_phv_out_data_175; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_176 = pipe4_io_pipe_phv_out_data_176; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_177 = pipe4_io_pipe_phv_out_data_177; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_178 = pipe4_io_pipe_phv_out_data_178; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_179 = pipe4_io_pipe_phv_out_data_179; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_180 = pipe4_io_pipe_phv_out_data_180; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_181 = pipe4_io_pipe_phv_out_data_181; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_182 = pipe4_io_pipe_phv_out_data_182; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_183 = pipe4_io_pipe_phv_out_data_183; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_184 = pipe4_io_pipe_phv_out_data_184; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_185 = pipe4_io_pipe_phv_out_data_185; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_186 = pipe4_io_pipe_phv_out_data_186; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_187 = pipe4_io_pipe_phv_out_data_187; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_188 = pipe4_io_pipe_phv_out_data_188; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_189 = pipe4_io_pipe_phv_out_data_189; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_190 = pipe4_io_pipe_phv_out_data_190; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_191 = pipe4_io_pipe_phv_out_data_191; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_192 = pipe4_io_pipe_phv_out_data_192; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_193 = pipe4_io_pipe_phv_out_data_193; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_194 = pipe4_io_pipe_phv_out_data_194; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_195 = pipe4_io_pipe_phv_out_data_195; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_196 = pipe4_io_pipe_phv_out_data_196; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_197 = pipe4_io_pipe_phv_out_data_197; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_198 = pipe4_io_pipe_phv_out_data_198; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_199 = pipe4_io_pipe_phv_out_data_199; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_200 = pipe4_io_pipe_phv_out_data_200; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_201 = pipe4_io_pipe_phv_out_data_201; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_202 = pipe4_io_pipe_phv_out_data_202; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_203 = pipe4_io_pipe_phv_out_data_203; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_204 = pipe4_io_pipe_phv_out_data_204; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_205 = pipe4_io_pipe_phv_out_data_205; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_206 = pipe4_io_pipe_phv_out_data_206; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_207 = pipe4_io_pipe_phv_out_data_207; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_208 = pipe4_io_pipe_phv_out_data_208; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_209 = pipe4_io_pipe_phv_out_data_209; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_210 = pipe4_io_pipe_phv_out_data_210; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_211 = pipe4_io_pipe_phv_out_data_211; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_212 = pipe4_io_pipe_phv_out_data_212; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_213 = pipe4_io_pipe_phv_out_data_213; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_214 = pipe4_io_pipe_phv_out_data_214; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_215 = pipe4_io_pipe_phv_out_data_215; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_216 = pipe4_io_pipe_phv_out_data_216; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_217 = pipe4_io_pipe_phv_out_data_217; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_218 = pipe4_io_pipe_phv_out_data_218; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_219 = pipe4_io_pipe_phv_out_data_219; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_220 = pipe4_io_pipe_phv_out_data_220; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_221 = pipe4_io_pipe_phv_out_data_221; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_222 = pipe4_io_pipe_phv_out_data_222; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_223 = pipe4_io_pipe_phv_out_data_223; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_224 = pipe4_io_pipe_phv_out_data_224; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_225 = pipe4_io_pipe_phv_out_data_225; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_226 = pipe4_io_pipe_phv_out_data_226; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_227 = pipe4_io_pipe_phv_out_data_227; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_228 = pipe4_io_pipe_phv_out_data_228; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_229 = pipe4_io_pipe_phv_out_data_229; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_230 = pipe4_io_pipe_phv_out_data_230; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_231 = pipe4_io_pipe_phv_out_data_231; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_232 = pipe4_io_pipe_phv_out_data_232; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_233 = pipe4_io_pipe_phv_out_data_233; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_234 = pipe4_io_pipe_phv_out_data_234; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_235 = pipe4_io_pipe_phv_out_data_235; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_236 = pipe4_io_pipe_phv_out_data_236; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_237 = pipe4_io_pipe_phv_out_data_237; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_238 = pipe4_io_pipe_phv_out_data_238; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_239 = pipe4_io_pipe_phv_out_data_239; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_240 = pipe4_io_pipe_phv_out_data_240; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_241 = pipe4_io_pipe_phv_out_data_241; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_242 = pipe4_io_pipe_phv_out_data_242; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_243 = pipe4_io_pipe_phv_out_data_243; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_244 = pipe4_io_pipe_phv_out_data_244; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_245 = pipe4_io_pipe_phv_out_data_245; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_246 = pipe4_io_pipe_phv_out_data_246; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_247 = pipe4_io_pipe_phv_out_data_247; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_248 = pipe4_io_pipe_phv_out_data_248; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_249 = pipe4_io_pipe_phv_out_data_249; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_250 = pipe4_io_pipe_phv_out_data_250; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_251 = pipe4_io_pipe_phv_out_data_251; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_252 = pipe4_io_pipe_phv_out_data_252; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_253 = pipe4_io_pipe_phv_out_data_253; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_254 = pipe4_io_pipe_phv_out_data_254; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_255 = pipe4_io_pipe_phv_out_data_255; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_256 = pipe4_io_pipe_phv_out_data_256; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_257 = pipe4_io_pipe_phv_out_data_257; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_258 = pipe4_io_pipe_phv_out_data_258; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_259 = pipe4_io_pipe_phv_out_data_259; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_260 = pipe4_io_pipe_phv_out_data_260; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_261 = pipe4_io_pipe_phv_out_data_261; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_262 = pipe4_io_pipe_phv_out_data_262; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_263 = pipe4_io_pipe_phv_out_data_263; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_264 = pipe4_io_pipe_phv_out_data_264; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_265 = pipe4_io_pipe_phv_out_data_265; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_266 = pipe4_io_pipe_phv_out_data_266; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_267 = pipe4_io_pipe_phv_out_data_267; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_268 = pipe4_io_pipe_phv_out_data_268; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_269 = pipe4_io_pipe_phv_out_data_269; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_270 = pipe4_io_pipe_phv_out_data_270; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_271 = pipe4_io_pipe_phv_out_data_271; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_272 = pipe4_io_pipe_phv_out_data_272; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_273 = pipe4_io_pipe_phv_out_data_273; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_274 = pipe4_io_pipe_phv_out_data_274; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_275 = pipe4_io_pipe_phv_out_data_275; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_276 = pipe4_io_pipe_phv_out_data_276; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_277 = pipe4_io_pipe_phv_out_data_277; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_278 = pipe4_io_pipe_phv_out_data_278; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_279 = pipe4_io_pipe_phv_out_data_279; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_280 = pipe4_io_pipe_phv_out_data_280; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_281 = pipe4_io_pipe_phv_out_data_281; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_282 = pipe4_io_pipe_phv_out_data_282; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_283 = pipe4_io_pipe_phv_out_data_283; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_284 = pipe4_io_pipe_phv_out_data_284; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_285 = pipe4_io_pipe_phv_out_data_285; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_286 = pipe4_io_pipe_phv_out_data_286; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_287 = pipe4_io_pipe_phv_out_data_287; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_288 = pipe4_io_pipe_phv_out_data_288; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_289 = pipe4_io_pipe_phv_out_data_289; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_290 = pipe4_io_pipe_phv_out_data_290; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_291 = pipe4_io_pipe_phv_out_data_291; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_292 = pipe4_io_pipe_phv_out_data_292; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_293 = pipe4_io_pipe_phv_out_data_293; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_294 = pipe4_io_pipe_phv_out_data_294; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_295 = pipe4_io_pipe_phv_out_data_295; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_296 = pipe4_io_pipe_phv_out_data_296; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_297 = pipe4_io_pipe_phv_out_data_297; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_298 = pipe4_io_pipe_phv_out_data_298; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_299 = pipe4_io_pipe_phv_out_data_299; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_300 = pipe4_io_pipe_phv_out_data_300; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_301 = pipe4_io_pipe_phv_out_data_301; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_302 = pipe4_io_pipe_phv_out_data_302; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_303 = pipe4_io_pipe_phv_out_data_303; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_304 = pipe4_io_pipe_phv_out_data_304; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_305 = pipe4_io_pipe_phv_out_data_305; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_306 = pipe4_io_pipe_phv_out_data_306; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_307 = pipe4_io_pipe_phv_out_data_307; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_308 = pipe4_io_pipe_phv_out_data_308; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_309 = pipe4_io_pipe_phv_out_data_309; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_310 = pipe4_io_pipe_phv_out_data_310; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_311 = pipe4_io_pipe_phv_out_data_311; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_312 = pipe4_io_pipe_phv_out_data_312; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_313 = pipe4_io_pipe_phv_out_data_313; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_314 = pipe4_io_pipe_phv_out_data_314; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_315 = pipe4_io_pipe_phv_out_data_315; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_316 = pipe4_io_pipe_phv_out_data_316; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_317 = pipe4_io_pipe_phv_out_data_317; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_318 = pipe4_io_pipe_phv_out_data_318; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_319 = pipe4_io_pipe_phv_out_data_319; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_320 = pipe4_io_pipe_phv_out_data_320; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_321 = pipe4_io_pipe_phv_out_data_321; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_322 = pipe4_io_pipe_phv_out_data_322; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_323 = pipe4_io_pipe_phv_out_data_323; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_324 = pipe4_io_pipe_phv_out_data_324; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_325 = pipe4_io_pipe_phv_out_data_325; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_326 = pipe4_io_pipe_phv_out_data_326; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_327 = pipe4_io_pipe_phv_out_data_327; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_328 = pipe4_io_pipe_phv_out_data_328; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_329 = pipe4_io_pipe_phv_out_data_329; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_330 = pipe4_io_pipe_phv_out_data_330; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_331 = pipe4_io_pipe_phv_out_data_331; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_332 = pipe4_io_pipe_phv_out_data_332; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_333 = pipe4_io_pipe_phv_out_data_333; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_334 = pipe4_io_pipe_phv_out_data_334; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_335 = pipe4_io_pipe_phv_out_data_335; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_336 = pipe4_io_pipe_phv_out_data_336; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_337 = pipe4_io_pipe_phv_out_data_337; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_338 = pipe4_io_pipe_phv_out_data_338; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_339 = pipe4_io_pipe_phv_out_data_339; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_340 = pipe4_io_pipe_phv_out_data_340; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_341 = pipe4_io_pipe_phv_out_data_341; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_342 = pipe4_io_pipe_phv_out_data_342; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_343 = pipe4_io_pipe_phv_out_data_343; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_344 = pipe4_io_pipe_phv_out_data_344; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_345 = pipe4_io_pipe_phv_out_data_345; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_346 = pipe4_io_pipe_phv_out_data_346; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_347 = pipe4_io_pipe_phv_out_data_347; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_348 = pipe4_io_pipe_phv_out_data_348; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_349 = pipe4_io_pipe_phv_out_data_349; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_350 = pipe4_io_pipe_phv_out_data_350; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_351 = pipe4_io_pipe_phv_out_data_351; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_352 = pipe4_io_pipe_phv_out_data_352; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_353 = pipe4_io_pipe_phv_out_data_353; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_354 = pipe4_io_pipe_phv_out_data_354; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_355 = pipe4_io_pipe_phv_out_data_355; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_356 = pipe4_io_pipe_phv_out_data_356; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_357 = pipe4_io_pipe_phv_out_data_357; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_358 = pipe4_io_pipe_phv_out_data_358; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_359 = pipe4_io_pipe_phv_out_data_359; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_360 = pipe4_io_pipe_phv_out_data_360; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_361 = pipe4_io_pipe_phv_out_data_361; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_362 = pipe4_io_pipe_phv_out_data_362; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_363 = pipe4_io_pipe_phv_out_data_363; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_364 = pipe4_io_pipe_phv_out_data_364; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_365 = pipe4_io_pipe_phv_out_data_365; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_366 = pipe4_io_pipe_phv_out_data_366; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_367 = pipe4_io_pipe_phv_out_data_367; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_368 = pipe4_io_pipe_phv_out_data_368; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_369 = pipe4_io_pipe_phv_out_data_369; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_370 = pipe4_io_pipe_phv_out_data_370; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_371 = pipe4_io_pipe_phv_out_data_371; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_372 = pipe4_io_pipe_phv_out_data_372; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_373 = pipe4_io_pipe_phv_out_data_373; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_374 = pipe4_io_pipe_phv_out_data_374; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_375 = pipe4_io_pipe_phv_out_data_375; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_376 = pipe4_io_pipe_phv_out_data_376; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_377 = pipe4_io_pipe_phv_out_data_377; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_378 = pipe4_io_pipe_phv_out_data_378; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_379 = pipe4_io_pipe_phv_out_data_379; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_380 = pipe4_io_pipe_phv_out_data_380; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_381 = pipe4_io_pipe_phv_out_data_381; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_382 = pipe4_io_pipe_phv_out_data_382; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_383 = pipe4_io_pipe_phv_out_data_383; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_384 = pipe4_io_pipe_phv_out_data_384; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_385 = pipe4_io_pipe_phv_out_data_385; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_386 = pipe4_io_pipe_phv_out_data_386; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_387 = pipe4_io_pipe_phv_out_data_387; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_388 = pipe4_io_pipe_phv_out_data_388; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_389 = pipe4_io_pipe_phv_out_data_389; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_390 = pipe4_io_pipe_phv_out_data_390; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_391 = pipe4_io_pipe_phv_out_data_391; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_392 = pipe4_io_pipe_phv_out_data_392; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_393 = pipe4_io_pipe_phv_out_data_393; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_394 = pipe4_io_pipe_phv_out_data_394; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_395 = pipe4_io_pipe_phv_out_data_395; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_396 = pipe4_io_pipe_phv_out_data_396; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_397 = pipe4_io_pipe_phv_out_data_397; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_398 = pipe4_io_pipe_phv_out_data_398; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_399 = pipe4_io_pipe_phv_out_data_399; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_400 = pipe4_io_pipe_phv_out_data_400; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_401 = pipe4_io_pipe_phv_out_data_401; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_402 = pipe4_io_pipe_phv_out_data_402; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_403 = pipe4_io_pipe_phv_out_data_403; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_404 = pipe4_io_pipe_phv_out_data_404; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_405 = pipe4_io_pipe_phv_out_data_405; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_406 = pipe4_io_pipe_phv_out_data_406; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_407 = pipe4_io_pipe_phv_out_data_407; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_408 = pipe4_io_pipe_phv_out_data_408; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_409 = pipe4_io_pipe_phv_out_data_409; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_410 = pipe4_io_pipe_phv_out_data_410; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_411 = pipe4_io_pipe_phv_out_data_411; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_412 = pipe4_io_pipe_phv_out_data_412; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_413 = pipe4_io_pipe_phv_out_data_413; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_414 = pipe4_io_pipe_phv_out_data_414; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_415 = pipe4_io_pipe_phv_out_data_415; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_416 = pipe4_io_pipe_phv_out_data_416; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_417 = pipe4_io_pipe_phv_out_data_417; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_418 = pipe4_io_pipe_phv_out_data_418; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_419 = pipe4_io_pipe_phv_out_data_419; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_420 = pipe4_io_pipe_phv_out_data_420; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_421 = pipe4_io_pipe_phv_out_data_421; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_422 = pipe4_io_pipe_phv_out_data_422; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_423 = pipe4_io_pipe_phv_out_data_423; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_424 = pipe4_io_pipe_phv_out_data_424; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_425 = pipe4_io_pipe_phv_out_data_425; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_426 = pipe4_io_pipe_phv_out_data_426; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_427 = pipe4_io_pipe_phv_out_data_427; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_428 = pipe4_io_pipe_phv_out_data_428; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_429 = pipe4_io_pipe_phv_out_data_429; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_430 = pipe4_io_pipe_phv_out_data_430; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_431 = pipe4_io_pipe_phv_out_data_431; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_432 = pipe4_io_pipe_phv_out_data_432; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_433 = pipe4_io_pipe_phv_out_data_433; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_434 = pipe4_io_pipe_phv_out_data_434; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_435 = pipe4_io_pipe_phv_out_data_435; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_436 = pipe4_io_pipe_phv_out_data_436; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_437 = pipe4_io_pipe_phv_out_data_437; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_438 = pipe4_io_pipe_phv_out_data_438; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_439 = pipe4_io_pipe_phv_out_data_439; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_440 = pipe4_io_pipe_phv_out_data_440; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_441 = pipe4_io_pipe_phv_out_data_441; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_442 = pipe4_io_pipe_phv_out_data_442; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_443 = pipe4_io_pipe_phv_out_data_443; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_444 = pipe4_io_pipe_phv_out_data_444; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_445 = pipe4_io_pipe_phv_out_data_445; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_446 = pipe4_io_pipe_phv_out_data_446; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_447 = pipe4_io_pipe_phv_out_data_447; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_448 = pipe4_io_pipe_phv_out_data_448; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_449 = pipe4_io_pipe_phv_out_data_449; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_450 = pipe4_io_pipe_phv_out_data_450; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_451 = pipe4_io_pipe_phv_out_data_451; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_452 = pipe4_io_pipe_phv_out_data_452; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_453 = pipe4_io_pipe_phv_out_data_453; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_454 = pipe4_io_pipe_phv_out_data_454; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_455 = pipe4_io_pipe_phv_out_data_455; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_456 = pipe4_io_pipe_phv_out_data_456; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_457 = pipe4_io_pipe_phv_out_data_457; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_458 = pipe4_io_pipe_phv_out_data_458; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_459 = pipe4_io_pipe_phv_out_data_459; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_460 = pipe4_io_pipe_phv_out_data_460; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_461 = pipe4_io_pipe_phv_out_data_461; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_462 = pipe4_io_pipe_phv_out_data_462; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_463 = pipe4_io_pipe_phv_out_data_463; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_464 = pipe4_io_pipe_phv_out_data_464; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_465 = pipe4_io_pipe_phv_out_data_465; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_466 = pipe4_io_pipe_phv_out_data_466; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_467 = pipe4_io_pipe_phv_out_data_467; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_468 = pipe4_io_pipe_phv_out_data_468; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_469 = pipe4_io_pipe_phv_out_data_469; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_470 = pipe4_io_pipe_phv_out_data_470; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_471 = pipe4_io_pipe_phv_out_data_471; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_472 = pipe4_io_pipe_phv_out_data_472; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_473 = pipe4_io_pipe_phv_out_data_473; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_474 = pipe4_io_pipe_phv_out_data_474; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_475 = pipe4_io_pipe_phv_out_data_475; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_476 = pipe4_io_pipe_phv_out_data_476; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_477 = pipe4_io_pipe_phv_out_data_477; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_478 = pipe4_io_pipe_phv_out_data_478; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_479 = pipe4_io_pipe_phv_out_data_479; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_480 = pipe4_io_pipe_phv_out_data_480; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_481 = pipe4_io_pipe_phv_out_data_481; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_482 = pipe4_io_pipe_phv_out_data_482; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_483 = pipe4_io_pipe_phv_out_data_483; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_484 = pipe4_io_pipe_phv_out_data_484; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_485 = pipe4_io_pipe_phv_out_data_485; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_486 = pipe4_io_pipe_phv_out_data_486; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_487 = pipe4_io_pipe_phv_out_data_487; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_488 = pipe4_io_pipe_phv_out_data_488; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_489 = pipe4_io_pipe_phv_out_data_489; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_490 = pipe4_io_pipe_phv_out_data_490; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_491 = pipe4_io_pipe_phv_out_data_491; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_492 = pipe4_io_pipe_phv_out_data_492; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_493 = pipe4_io_pipe_phv_out_data_493; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_494 = pipe4_io_pipe_phv_out_data_494; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_495 = pipe4_io_pipe_phv_out_data_495; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_496 = pipe4_io_pipe_phv_out_data_496; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_497 = pipe4_io_pipe_phv_out_data_497; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_498 = pipe4_io_pipe_phv_out_data_498; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_499 = pipe4_io_pipe_phv_out_data_499; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_500 = pipe4_io_pipe_phv_out_data_500; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_501 = pipe4_io_pipe_phv_out_data_501; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_502 = pipe4_io_pipe_phv_out_data_502; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_503 = pipe4_io_pipe_phv_out_data_503; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_504 = pipe4_io_pipe_phv_out_data_504; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_505 = pipe4_io_pipe_phv_out_data_505; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_506 = pipe4_io_pipe_phv_out_data_506; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_507 = pipe4_io_pipe_phv_out_data_507; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_508 = pipe4_io_pipe_phv_out_data_508; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_509 = pipe4_io_pipe_phv_out_data_509; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_510 = pipe4_io_pipe_phv_out_data_510; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_511 = pipe4_io_pipe_phv_out_data_511; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 152:27]
  assign pipe5_io_hash_depth_0 = hash_depth_0; // @[hash.scala 156:27]
  assign pipe5_io_hash_depth_1 = hash_depth_1; // @[hash.scala 156:27]
  assign pipe5_io_key_in = pipe4_io_key_out; // @[hash.scala 153:27]
  assign pipe5_io_sum_in = pipe4_io_sum_out[15:0]; // @[hash.scala 154:27]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_96 = pipe5_io_pipe_phv_out_data_96; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_97 = pipe5_io_pipe_phv_out_data_97; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_98 = pipe5_io_pipe_phv_out_data_98; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_99 = pipe5_io_pipe_phv_out_data_99; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_100 = pipe5_io_pipe_phv_out_data_100; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_101 = pipe5_io_pipe_phv_out_data_101; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_102 = pipe5_io_pipe_phv_out_data_102; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_103 = pipe5_io_pipe_phv_out_data_103; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_104 = pipe5_io_pipe_phv_out_data_104; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_105 = pipe5_io_pipe_phv_out_data_105; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_106 = pipe5_io_pipe_phv_out_data_106; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_107 = pipe5_io_pipe_phv_out_data_107; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_108 = pipe5_io_pipe_phv_out_data_108; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_109 = pipe5_io_pipe_phv_out_data_109; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_110 = pipe5_io_pipe_phv_out_data_110; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_111 = pipe5_io_pipe_phv_out_data_111; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_112 = pipe5_io_pipe_phv_out_data_112; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_113 = pipe5_io_pipe_phv_out_data_113; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_114 = pipe5_io_pipe_phv_out_data_114; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_115 = pipe5_io_pipe_phv_out_data_115; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_116 = pipe5_io_pipe_phv_out_data_116; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_117 = pipe5_io_pipe_phv_out_data_117; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_118 = pipe5_io_pipe_phv_out_data_118; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_119 = pipe5_io_pipe_phv_out_data_119; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_120 = pipe5_io_pipe_phv_out_data_120; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_121 = pipe5_io_pipe_phv_out_data_121; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_122 = pipe5_io_pipe_phv_out_data_122; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_123 = pipe5_io_pipe_phv_out_data_123; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_124 = pipe5_io_pipe_phv_out_data_124; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_125 = pipe5_io_pipe_phv_out_data_125; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_126 = pipe5_io_pipe_phv_out_data_126; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_127 = pipe5_io_pipe_phv_out_data_127; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_128 = pipe5_io_pipe_phv_out_data_128; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_129 = pipe5_io_pipe_phv_out_data_129; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_130 = pipe5_io_pipe_phv_out_data_130; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_131 = pipe5_io_pipe_phv_out_data_131; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_132 = pipe5_io_pipe_phv_out_data_132; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_133 = pipe5_io_pipe_phv_out_data_133; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_134 = pipe5_io_pipe_phv_out_data_134; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_135 = pipe5_io_pipe_phv_out_data_135; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_136 = pipe5_io_pipe_phv_out_data_136; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_137 = pipe5_io_pipe_phv_out_data_137; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_138 = pipe5_io_pipe_phv_out_data_138; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_139 = pipe5_io_pipe_phv_out_data_139; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_140 = pipe5_io_pipe_phv_out_data_140; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_141 = pipe5_io_pipe_phv_out_data_141; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_142 = pipe5_io_pipe_phv_out_data_142; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_143 = pipe5_io_pipe_phv_out_data_143; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_144 = pipe5_io_pipe_phv_out_data_144; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_145 = pipe5_io_pipe_phv_out_data_145; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_146 = pipe5_io_pipe_phv_out_data_146; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_147 = pipe5_io_pipe_phv_out_data_147; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_148 = pipe5_io_pipe_phv_out_data_148; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_149 = pipe5_io_pipe_phv_out_data_149; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_150 = pipe5_io_pipe_phv_out_data_150; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_151 = pipe5_io_pipe_phv_out_data_151; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_152 = pipe5_io_pipe_phv_out_data_152; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_153 = pipe5_io_pipe_phv_out_data_153; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_154 = pipe5_io_pipe_phv_out_data_154; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_155 = pipe5_io_pipe_phv_out_data_155; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_156 = pipe5_io_pipe_phv_out_data_156; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_157 = pipe5_io_pipe_phv_out_data_157; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_158 = pipe5_io_pipe_phv_out_data_158; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_159 = pipe5_io_pipe_phv_out_data_159; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_160 = pipe5_io_pipe_phv_out_data_160; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_161 = pipe5_io_pipe_phv_out_data_161; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_162 = pipe5_io_pipe_phv_out_data_162; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_163 = pipe5_io_pipe_phv_out_data_163; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_164 = pipe5_io_pipe_phv_out_data_164; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_165 = pipe5_io_pipe_phv_out_data_165; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_166 = pipe5_io_pipe_phv_out_data_166; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_167 = pipe5_io_pipe_phv_out_data_167; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_168 = pipe5_io_pipe_phv_out_data_168; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_169 = pipe5_io_pipe_phv_out_data_169; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_170 = pipe5_io_pipe_phv_out_data_170; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_171 = pipe5_io_pipe_phv_out_data_171; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_172 = pipe5_io_pipe_phv_out_data_172; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_173 = pipe5_io_pipe_phv_out_data_173; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_174 = pipe5_io_pipe_phv_out_data_174; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_175 = pipe5_io_pipe_phv_out_data_175; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_176 = pipe5_io_pipe_phv_out_data_176; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_177 = pipe5_io_pipe_phv_out_data_177; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_178 = pipe5_io_pipe_phv_out_data_178; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_179 = pipe5_io_pipe_phv_out_data_179; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_180 = pipe5_io_pipe_phv_out_data_180; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_181 = pipe5_io_pipe_phv_out_data_181; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_182 = pipe5_io_pipe_phv_out_data_182; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_183 = pipe5_io_pipe_phv_out_data_183; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_184 = pipe5_io_pipe_phv_out_data_184; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_185 = pipe5_io_pipe_phv_out_data_185; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_186 = pipe5_io_pipe_phv_out_data_186; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_187 = pipe5_io_pipe_phv_out_data_187; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_188 = pipe5_io_pipe_phv_out_data_188; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_189 = pipe5_io_pipe_phv_out_data_189; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_190 = pipe5_io_pipe_phv_out_data_190; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_191 = pipe5_io_pipe_phv_out_data_191; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_192 = pipe5_io_pipe_phv_out_data_192; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_193 = pipe5_io_pipe_phv_out_data_193; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_194 = pipe5_io_pipe_phv_out_data_194; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_195 = pipe5_io_pipe_phv_out_data_195; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_196 = pipe5_io_pipe_phv_out_data_196; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_197 = pipe5_io_pipe_phv_out_data_197; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_198 = pipe5_io_pipe_phv_out_data_198; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_199 = pipe5_io_pipe_phv_out_data_199; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_200 = pipe5_io_pipe_phv_out_data_200; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_201 = pipe5_io_pipe_phv_out_data_201; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_202 = pipe5_io_pipe_phv_out_data_202; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_203 = pipe5_io_pipe_phv_out_data_203; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_204 = pipe5_io_pipe_phv_out_data_204; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_205 = pipe5_io_pipe_phv_out_data_205; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_206 = pipe5_io_pipe_phv_out_data_206; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_207 = pipe5_io_pipe_phv_out_data_207; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_208 = pipe5_io_pipe_phv_out_data_208; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_209 = pipe5_io_pipe_phv_out_data_209; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_210 = pipe5_io_pipe_phv_out_data_210; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_211 = pipe5_io_pipe_phv_out_data_211; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_212 = pipe5_io_pipe_phv_out_data_212; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_213 = pipe5_io_pipe_phv_out_data_213; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_214 = pipe5_io_pipe_phv_out_data_214; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_215 = pipe5_io_pipe_phv_out_data_215; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_216 = pipe5_io_pipe_phv_out_data_216; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_217 = pipe5_io_pipe_phv_out_data_217; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_218 = pipe5_io_pipe_phv_out_data_218; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_219 = pipe5_io_pipe_phv_out_data_219; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_220 = pipe5_io_pipe_phv_out_data_220; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_221 = pipe5_io_pipe_phv_out_data_221; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_222 = pipe5_io_pipe_phv_out_data_222; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_223 = pipe5_io_pipe_phv_out_data_223; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_224 = pipe5_io_pipe_phv_out_data_224; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_225 = pipe5_io_pipe_phv_out_data_225; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_226 = pipe5_io_pipe_phv_out_data_226; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_227 = pipe5_io_pipe_phv_out_data_227; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_228 = pipe5_io_pipe_phv_out_data_228; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_229 = pipe5_io_pipe_phv_out_data_229; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_230 = pipe5_io_pipe_phv_out_data_230; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_231 = pipe5_io_pipe_phv_out_data_231; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_232 = pipe5_io_pipe_phv_out_data_232; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_233 = pipe5_io_pipe_phv_out_data_233; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_234 = pipe5_io_pipe_phv_out_data_234; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_235 = pipe5_io_pipe_phv_out_data_235; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_236 = pipe5_io_pipe_phv_out_data_236; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_237 = pipe5_io_pipe_phv_out_data_237; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_238 = pipe5_io_pipe_phv_out_data_238; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_239 = pipe5_io_pipe_phv_out_data_239; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_240 = pipe5_io_pipe_phv_out_data_240; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_241 = pipe5_io_pipe_phv_out_data_241; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_242 = pipe5_io_pipe_phv_out_data_242; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_243 = pipe5_io_pipe_phv_out_data_243; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_244 = pipe5_io_pipe_phv_out_data_244; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_245 = pipe5_io_pipe_phv_out_data_245; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_246 = pipe5_io_pipe_phv_out_data_246; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_247 = pipe5_io_pipe_phv_out_data_247; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_248 = pipe5_io_pipe_phv_out_data_248; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_249 = pipe5_io_pipe_phv_out_data_249; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_250 = pipe5_io_pipe_phv_out_data_250; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_251 = pipe5_io_pipe_phv_out_data_251; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_252 = pipe5_io_pipe_phv_out_data_252; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_253 = pipe5_io_pipe_phv_out_data_253; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_254 = pipe5_io_pipe_phv_out_data_254; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_255 = pipe5_io_pipe_phv_out_data_255; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_256 = pipe5_io_pipe_phv_out_data_256; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_257 = pipe5_io_pipe_phv_out_data_257; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_258 = pipe5_io_pipe_phv_out_data_258; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_259 = pipe5_io_pipe_phv_out_data_259; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_260 = pipe5_io_pipe_phv_out_data_260; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_261 = pipe5_io_pipe_phv_out_data_261; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_262 = pipe5_io_pipe_phv_out_data_262; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_263 = pipe5_io_pipe_phv_out_data_263; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_264 = pipe5_io_pipe_phv_out_data_264; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_265 = pipe5_io_pipe_phv_out_data_265; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_266 = pipe5_io_pipe_phv_out_data_266; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_267 = pipe5_io_pipe_phv_out_data_267; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_268 = pipe5_io_pipe_phv_out_data_268; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_269 = pipe5_io_pipe_phv_out_data_269; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_270 = pipe5_io_pipe_phv_out_data_270; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_271 = pipe5_io_pipe_phv_out_data_271; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_272 = pipe5_io_pipe_phv_out_data_272; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_273 = pipe5_io_pipe_phv_out_data_273; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_274 = pipe5_io_pipe_phv_out_data_274; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_275 = pipe5_io_pipe_phv_out_data_275; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_276 = pipe5_io_pipe_phv_out_data_276; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_277 = pipe5_io_pipe_phv_out_data_277; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_278 = pipe5_io_pipe_phv_out_data_278; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_279 = pipe5_io_pipe_phv_out_data_279; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_280 = pipe5_io_pipe_phv_out_data_280; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_281 = pipe5_io_pipe_phv_out_data_281; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_282 = pipe5_io_pipe_phv_out_data_282; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_283 = pipe5_io_pipe_phv_out_data_283; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_284 = pipe5_io_pipe_phv_out_data_284; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_285 = pipe5_io_pipe_phv_out_data_285; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_286 = pipe5_io_pipe_phv_out_data_286; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_287 = pipe5_io_pipe_phv_out_data_287; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_288 = pipe5_io_pipe_phv_out_data_288; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_289 = pipe5_io_pipe_phv_out_data_289; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_290 = pipe5_io_pipe_phv_out_data_290; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_291 = pipe5_io_pipe_phv_out_data_291; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_292 = pipe5_io_pipe_phv_out_data_292; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_293 = pipe5_io_pipe_phv_out_data_293; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_294 = pipe5_io_pipe_phv_out_data_294; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_295 = pipe5_io_pipe_phv_out_data_295; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_296 = pipe5_io_pipe_phv_out_data_296; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_297 = pipe5_io_pipe_phv_out_data_297; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_298 = pipe5_io_pipe_phv_out_data_298; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_299 = pipe5_io_pipe_phv_out_data_299; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_300 = pipe5_io_pipe_phv_out_data_300; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_301 = pipe5_io_pipe_phv_out_data_301; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_302 = pipe5_io_pipe_phv_out_data_302; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_303 = pipe5_io_pipe_phv_out_data_303; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_304 = pipe5_io_pipe_phv_out_data_304; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_305 = pipe5_io_pipe_phv_out_data_305; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_306 = pipe5_io_pipe_phv_out_data_306; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_307 = pipe5_io_pipe_phv_out_data_307; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_308 = pipe5_io_pipe_phv_out_data_308; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_309 = pipe5_io_pipe_phv_out_data_309; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_310 = pipe5_io_pipe_phv_out_data_310; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_311 = pipe5_io_pipe_phv_out_data_311; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_312 = pipe5_io_pipe_phv_out_data_312; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_313 = pipe5_io_pipe_phv_out_data_313; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_314 = pipe5_io_pipe_phv_out_data_314; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_315 = pipe5_io_pipe_phv_out_data_315; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_316 = pipe5_io_pipe_phv_out_data_316; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_317 = pipe5_io_pipe_phv_out_data_317; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_318 = pipe5_io_pipe_phv_out_data_318; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_319 = pipe5_io_pipe_phv_out_data_319; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_320 = pipe5_io_pipe_phv_out_data_320; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_321 = pipe5_io_pipe_phv_out_data_321; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_322 = pipe5_io_pipe_phv_out_data_322; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_323 = pipe5_io_pipe_phv_out_data_323; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_324 = pipe5_io_pipe_phv_out_data_324; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_325 = pipe5_io_pipe_phv_out_data_325; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_326 = pipe5_io_pipe_phv_out_data_326; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_327 = pipe5_io_pipe_phv_out_data_327; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_328 = pipe5_io_pipe_phv_out_data_328; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_329 = pipe5_io_pipe_phv_out_data_329; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_330 = pipe5_io_pipe_phv_out_data_330; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_331 = pipe5_io_pipe_phv_out_data_331; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_332 = pipe5_io_pipe_phv_out_data_332; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_333 = pipe5_io_pipe_phv_out_data_333; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_334 = pipe5_io_pipe_phv_out_data_334; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_335 = pipe5_io_pipe_phv_out_data_335; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_336 = pipe5_io_pipe_phv_out_data_336; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_337 = pipe5_io_pipe_phv_out_data_337; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_338 = pipe5_io_pipe_phv_out_data_338; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_339 = pipe5_io_pipe_phv_out_data_339; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_340 = pipe5_io_pipe_phv_out_data_340; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_341 = pipe5_io_pipe_phv_out_data_341; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_342 = pipe5_io_pipe_phv_out_data_342; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_343 = pipe5_io_pipe_phv_out_data_343; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_344 = pipe5_io_pipe_phv_out_data_344; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_345 = pipe5_io_pipe_phv_out_data_345; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_346 = pipe5_io_pipe_phv_out_data_346; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_347 = pipe5_io_pipe_phv_out_data_347; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_348 = pipe5_io_pipe_phv_out_data_348; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_349 = pipe5_io_pipe_phv_out_data_349; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_350 = pipe5_io_pipe_phv_out_data_350; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_351 = pipe5_io_pipe_phv_out_data_351; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_352 = pipe5_io_pipe_phv_out_data_352; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_353 = pipe5_io_pipe_phv_out_data_353; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_354 = pipe5_io_pipe_phv_out_data_354; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_355 = pipe5_io_pipe_phv_out_data_355; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_356 = pipe5_io_pipe_phv_out_data_356; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_357 = pipe5_io_pipe_phv_out_data_357; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_358 = pipe5_io_pipe_phv_out_data_358; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_359 = pipe5_io_pipe_phv_out_data_359; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_360 = pipe5_io_pipe_phv_out_data_360; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_361 = pipe5_io_pipe_phv_out_data_361; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_362 = pipe5_io_pipe_phv_out_data_362; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_363 = pipe5_io_pipe_phv_out_data_363; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_364 = pipe5_io_pipe_phv_out_data_364; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_365 = pipe5_io_pipe_phv_out_data_365; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_366 = pipe5_io_pipe_phv_out_data_366; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_367 = pipe5_io_pipe_phv_out_data_367; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_368 = pipe5_io_pipe_phv_out_data_368; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_369 = pipe5_io_pipe_phv_out_data_369; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_370 = pipe5_io_pipe_phv_out_data_370; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_371 = pipe5_io_pipe_phv_out_data_371; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_372 = pipe5_io_pipe_phv_out_data_372; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_373 = pipe5_io_pipe_phv_out_data_373; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_374 = pipe5_io_pipe_phv_out_data_374; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_375 = pipe5_io_pipe_phv_out_data_375; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_376 = pipe5_io_pipe_phv_out_data_376; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_377 = pipe5_io_pipe_phv_out_data_377; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_378 = pipe5_io_pipe_phv_out_data_378; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_379 = pipe5_io_pipe_phv_out_data_379; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_380 = pipe5_io_pipe_phv_out_data_380; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_381 = pipe5_io_pipe_phv_out_data_381; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_382 = pipe5_io_pipe_phv_out_data_382; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_383 = pipe5_io_pipe_phv_out_data_383; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_384 = pipe5_io_pipe_phv_out_data_384; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_385 = pipe5_io_pipe_phv_out_data_385; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_386 = pipe5_io_pipe_phv_out_data_386; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_387 = pipe5_io_pipe_phv_out_data_387; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_388 = pipe5_io_pipe_phv_out_data_388; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_389 = pipe5_io_pipe_phv_out_data_389; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_390 = pipe5_io_pipe_phv_out_data_390; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_391 = pipe5_io_pipe_phv_out_data_391; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_392 = pipe5_io_pipe_phv_out_data_392; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_393 = pipe5_io_pipe_phv_out_data_393; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_394 = pipe5_io_pipe_phv_out_data_394; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_395 = pipe5_io_pipe_phv_out_data_395; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_396 = pipe5_io_pipe_phv_out_data_396; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_397 = pipe5_io_pipe_phv_out_data_397; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_398 = pipe5_io_pipe_phv_out_data_398; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_399 = pipe5_io_pipe_phv_out_data_399; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_400 = pipe5_io_pipe_phv_out_data_400; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_401 = pipe5_io_pipe_phv_out_data_401; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_402 = pipe5_io_pipe_phv_out_data_402; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_403 = pipe5_io_pipe_phv_out_data_403; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_404 = pipe5_io_pipe_phv_out_data_404; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_405 = pipe5_io_pipe_phv_out_data_405; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_406 = pipe5_io_pipe_phv_out_data_406; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_407 = pipe5_io_pipe_phv_out_data_407; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_408 = pipe5_io_pipe_phv_out_data_408; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_409 = pipe5_io_pipe_phv_out_data_409; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_410 = pipe5_io_pipe_phv_out_data_410; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_411 = pipe5_io_pipe_phv_out_data_411; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_412 = pipe5_io_pipe_phv_out_data_412; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_413 = pipe5_io_pipe_phv_out_data_413; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_414 = pipe5_io_pipe_phv_out_data_414; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_415 = pipe5_io_pipe_phv_out_data_415; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_416 = pipe5_io_pipe_phv_out_data_416; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_417 = pipe5_io_pipe_phv_out_data_417; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_418 = pipe5_io_pipe_phv_out_data_418; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_419 = pipe5_io_pipe_phv_out_data_419; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_420 = pipe5_io_pipe_phv_out_data_420; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_421 = pipe5_io_pipe_phv_out_data_421; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_422 = pipe5_io_pipe_phv_out_data_422; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_423 = pipe5_io_pipe_phv_out_data_423; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_424 = pipe5_io_pipe_phv_out_data_424; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_425 = pipe5_io_pipe_phv_out_data_425; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_426 = pipe5_io_pipe_phv_out_data_426; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_427 = pipe5_io_pipe_phv_out_data_427; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_428 = pipe5_io_pipe_phv_out_data_428; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_429 = pipe5_io_pipe_phv_out_data_429; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_430 = pipe5_io_pipe_phv_out_data_430; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_431 = pipe5_io_pipe_phv_out_data_431; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_432 = pipe5_io_pipe_phv_out_data_432; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_433 = pipe5_io_pipe_phv_out_data_433; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_434 = pipe5_io_pipe_phv_out_data_434; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_435 = pipe5_io_pipe_phv_out_data_435; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_436 = pipe5_io_pipe_phv_out_data_436; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_437 = pipe5_io_pipe_phv_out_data_437; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_438 = pipe5_io_pipe_phv_out_data_438; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_439 = pipe5_io_pipe_phv_out_data_439; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_440 = pipe5_io_pipe_phv_out_data_440; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_441 = pipe5_io_pipe_phv_out_data_441; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_442 = pipe5_io_pipe_phv_out_data_442; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_443 = pipe5_io_pipe_phv_out_data_443; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_444 = pipe5_io_pipe_phv_out_data_444; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_445 = pipe5_io_pipe_phv_out_data_445; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_446 = pipe5_io_pipe_phv_out_data_446; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_447 = pipe5_io_pipe_phv_out_data_447; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_448 = pipe5_io_pipe_phv_out_data_448; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_449 = pipe5_io_pipe_phv_out_data_449; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_450 = pipe5_io_pipe_phv_out_data_450; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_451 = pipe5_io_pipe_phv_out_data_451; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_452 = pipe5_io_pipe_phv_out_data_452; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_453 = pipe5_io_pipe_phv_out_data_453; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_454 = pipe5_io_pipe_phv_out_data_454; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_455 = pipe5_io_pipe_phv_out_data_455; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_456 = pipe5_io_pipe_phv_out_data_456; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_457 = pipe5_io_pipe_phv_out_data_457; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_458 = pipe5_io_pipe_phv_out_data_458; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_459 = pipe5_io_pipe_phv_out_data_459; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_460 = pipe5_io_pipe_phv_out_data_460; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_461 = pipe5_io_pipe_phv_out_data_461; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_462 = pipe5_io_pipe_phv_out_data_462; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_463 = pipe5_io_pipe_phv_out_data_463; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_464 = pipe5_io_pipe_phv_out_data_464; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_465 = pipe5_io_pipe_phv_out_data_465; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_466 = pipe5_io_pipe_phv_out_data_466; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_467 = pipe5_io_pipe_phv_out_data_467; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_468 = pipe5_io_pipe_phv_out_data_468; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_469 = pipe5_io_pipe_phv_out_data_469; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_470 = pipe5_io_pipe_phv_out_data_470; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_471 = pipe5_io_pipe_phv_out_data_471; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_472 = pipe5_io_pipe_phv_out_data_472; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_473 = pipe5_io_pipe_phv_out_data_473; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_474 = pipe5_io_pipe_phv_out_data_474; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_475 = pipe5_io_pipe_phv_out_data_475; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_476 = pipe5_io_pipe_phv_out_data_476; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_477 = pipe5_io_pipe_phv_out_data_477; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_478 = pipe5_io_pipe_phv_out_data_478; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_479 = pipe5_io_pipe_phv_out_data_479; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_480 = pipe5_io_pipe_phv_out_data_480; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_481 = pipe5_io_pipe_phv_out_data_481; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_482 = pipe5_io_pipe_phv_out_data_482; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_483 = pipe5_io_pipe_phv_out_data_483; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_484 = pipe5_io_pipe_phv_out_data_484; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_485 = pipe5_io_pipe_phv_out_data_485; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_486 = pipe5_io_pipe_phv_out_data_486; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_487 = pipe5_io_pipe_phv_out_data_487; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_488 = pipe5_io_pipe_phv_out_data_488; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_489 = pipe5_io_pipe_phv_out_data_489; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_490 = pipe5_io_pipe_phv_out_data_490; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_491 = pipe5_io_pipe_phv_out_data_491; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_492 = pipe5_io_pipe_phv_out_data_492; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_493 = pipe5_io_pipe_phv_out_data_493; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_494 = pipe5_io_pipe_phv_out_data_494; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_495 = pipe5_io_pipe_phv_out_data_495; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_496 = pipe5_io_pipe_phv_out_data_496; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_497 = pipe5_io_pipe_phv_out_data_497; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_498 = pipe5_io_pipe_phv_out_data_498; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_499 = pipe5_io_pipe_phv_out_data_499; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_500 = pipe5_io_pipe_phv_out_data_500; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_501 = pipe5_io_pipe_phv_out_data_501; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_502 = pipe5_io_pipe_phv_out_data_502; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_503 = pipe5_io_pipe_phv_out_data_503; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_504 = pipe5_io_pipe_phv_out_data_504; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_505 = pipe5_io_pipe_phv_out_data_505; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_506 = pipe5_io_pipe_phv_out_data_506; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_507 = pipe5_io_pipe_phv_out_data_507; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_508 = pipe5_io_pipe_phv_out_data_508; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_509 = pipe5_io_pipe_phv_out_data_509; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_510 = pipe5_io_pipe_phv_out_data_510; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_511 = pipe5_io_pipe_phv_out_data_511; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 158:27]
  assign pipe6_io_hash_depth_0 = hash_depth_0; // @[hash.scala 162:27]
  assign pipe6_io_hash_depth_1 = hash_depth_1; // @[hash.scala 162:27]
  assign pipe6_io_key_in = pipe5_io_key_out; // @[hash.scala 159:27]
  assign pipe6_io_sum_in = pipe5_io_sum_out; // @[hash.scala 160:27]
  assign pipe6_io_val_in = pipe5_io_val_out; // @[hash.scala 161:27]
  assign pipe7_clock = clock;
  assign pipe7_io_pipe_phv_in_data_0 = pipe6_io_pipe_phv_out_data_0; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_1 = pipe6_io_pipe_phv_out_data_1; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_2 = pipe6_io_pipe_phv_out_data_2; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_3 = pipe6_io_pipe_phv_out_data_3; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_4 = pipe6_io_pipe_phv_out_data_4; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_5 = pipe6_io_pipe_phv_out_data_5; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_6 = pipe6_io_pipe_phv_out_data_6; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_7 = pipe6_io_pipe_phv_out_data_7; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_8 = pipe6_io_pipe_phv_out_data_8; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_9 = pipe6_io_pipe_phv_out_data_9; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_10 = pipe6_io_pipe_phv_out_data_10; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_11 = pipe6_io_pipe_phv_out_data_11; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_12 = pipe6_io_pipe_phv_out_data_12; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_13 = pipe6_io_pipe_phv_out_data_13; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_14 = pipe6_io_pipe_phv_out_data_14; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_15 = pipe6_io_pipe_phv_out_data_15; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_16 = pipe6_io_pipe_phv_out_data_16; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_17 = pipe6_io_pipe_phv_out_data_17; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_18 = pipe6_io_pipe_phv_out_data_18; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_19 = pipe6_io_pipe_phv_out_data_19; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_20 = pipe6_io_pipe_phv_out_data_20; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_21 = pipe6_io_pipe_phv_out_data_21; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_22 = pipe6_io_pipe_phv_out_data_22; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_23 = pipe6_io_pipe_phv_out_data_23; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_24 = pipe6_io_pipe_phv_out_data_24; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_25 = pipe6_io_pipe_phv_out_data_25; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_26 = pipe6_io_pipe_phv_out_data_26; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_27 = pipe6_io_pipe_phv_out_data_27; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_28 = pipe6_io_pipe_phv_out_data_28; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_29 = pipe6_io_pipe_phv_out_data_29; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_30 = pipe6_io_pipe_phv_out_data_30; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_31 = pipe6_io_pipe_phv_out_data_31; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_32 = pipe6_io_pipe_phv_out_data_32; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_33 = pipe6_io_pipe_phv_out_data_33; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_34 = pipe6_io_pipe_phv_out_data_34; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_35 = pipe6_io_pipe_phv_out_data_35; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_36 = pipe6_io_pipe_phv_out_data_36; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_37 = pipe6_io_pipe_phv_out_data_37; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_38 = pipe6_io_pipe_phv_out_data_38; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_39 = pipe6_io_pipe_phv_out_data_39; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_40 = pipe6_io_pipe_phv_out_data_40; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_41 = pipe6_io_pipe_phv_out_data_41; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_42 = pipe6_io_pipe_phv_out_data_42; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_43 = pipe6_io_pipe_phv_out_data_43; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_44 = pipe6_io_pipe_phv_out_data_44; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_45 = pipe6_io_pipe_phv_out_data_45; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_46 = pipe6_io_pipe_phv_out_data_46; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_47 = pipe6_io_pipe_phv_out_data_47; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_48 = pipe6_io_pipe_phv_out_data_48; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_49 = pipe6_io_pipe_phv_out_data_49; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_50 = pipe6_io_pipe_phv_out_data_50; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_51 = pipe6_io_pipe_phv_out_data_51; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_52 = pipe6_io_pipe_phv_out_data_52; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_53 = pipe6_io_pipe_phv_out_data_53; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_54 = pipe6_io_pipe_phv_out_data_54; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_55 = pipe6_io_pipe_phv_out_data_55; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_56 = pipe6_io_pipe_phv_out_data_56; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_57 = pipe6_io_pipe_phv_out_data_57; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_58 = pipe6_io_pipe_phv_out_data_58; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_59 = pipe6_io_pipe_phv_out_data_59; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_60 = pipe6_io_pipe_phv_out_data_60; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_61 = pipe6_io_pipe_phv_out_data_61; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_62 = pipe6_io_pipe_phv_out_data_62; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_63 = pipe6_io_pipe_phv_out_data_63; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_64 = pipe6_io_pipe_phv_out_data_64; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_65 = pipe6_io_pipe_phv_out_data_65; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_66 = pipe6_io_pipe_phv_out_data_66; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_67 = pipe6_io_pipe_phv_out_data_67; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_68 = pipe6_io_pipe_phv_out_data_68; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_69 = pipe6_io_pipe_phv_out_data_69; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_70 = pipe6_io_pipe_phv_out_data_70; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_71 = pipe6_io_pipe_phv_out_data_71; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_72 = pipe6_io_pipe_phv_out_data_72; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_73 = pipe6_io_pipe_phv_out_data_73; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_74 = pipe6_io_pipe_phv_out_data_74; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_75 = pipe6_io_pipe_phv_out_data_75; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_76 = pipe6_io_pipe_phv_out_data_76; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_77 = pipe6_io_pipe_phv_out_data_77; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_78 = pipe6_io_pipe_phv_out_data_78; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_79 = pipe6_io_pipe_phv_out_data_79; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_80 = pipe6_io_pipe_phv_out_data_80; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_81 = pipe6_io_pipe_phv_out_data_81; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_82 = pipe6_io_pipe_phv_out_data_82; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_83 = pipe6_io_pipe_phv_out_data_83; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_84 = pipe6_io_pipe_phv_out_data_84; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_85 = pipe6_io_pipe_phv_out_data_85; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_86 = pipe6_io_pipe_phv_out_data_86; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_87 = pipe6_io_pipe_phv_out_data_87; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_88 = pipe6_io_pipe_phv_out_data_88; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_89 = pipe6_io_pipe_phv_out_data_89; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_90 = pipe6_io_pipe_phv_out_data_90; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_91 = pipe6_io_pipe_phv_out_data_91; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_92 = pipe6_io_pipe_phv_out_data_92; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_93 = pipe6_io_pipe_phv_out_data_93; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_94 = pipe6_io_pipe_phv_out_data_94; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_95 = pipe6_io_pipe_phv_out_data_95; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_96 = pipe6_io_pipe_phv_out_data_96; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_97 = pipe6_io_pipe_phv_out_data_97; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_98 = pipe6_io_pipe_phv_out_data_98; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_99 = pipe6_io_pipe_phv_out_data_99; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_100 = pipe6_io_pipe_phv_out_data_100; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_101 = pipe6_io_pipe_phv_out_data_101; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_102 = pipe6_io_pipe_phv_out_data_102; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_103 = pipe6_io_pipe_phv_out_data_103; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_104 = pipe6_io_pipe_phv_out_data_104; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_105 = pipe6_io_pipe_phv_out_data_105; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_106 = pipe6_io_pipe_phv_out_data_106; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_107 = pipe6_io_pipe_phv_out_data_107; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_108 = pipe6_io_pipe_phv_out_data_108; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_109 = pipe6_io_pipe_phv_out_data_109; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_110 = pipe6_io_pipe_phv_out_data_110; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_111 = pipe6_io_pipe_phv_out_data_111; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_112 = pipe6_io_pipe_phv_out_data_112; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_113 = pipe6_io_pipe_phv_out_data_113; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_114 = pipe6_io_pipe_phv_out_data_114; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_115 = pipe6_io_pipe_phv_out_data_115; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_116 = pipe6_io_pipe_phv_out_data_116; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_117 = pipe6_io_pipe_phv_out_data_117; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_118 = pipe6_io_pipe_phv_out_data_118; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_119 = pipe6_io_pipe_phv_out_data_119; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_120 = pipe6_io_pipe_phv_out_data_120; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_121 = pipe6_io_pipe_phv_out_data_121; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_122 = pipe6_io_pipe_phv_out_data_122; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_123 = pipe6_io_pipe_phv_out_data_123; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_124 = pipe6_io_pipe_phv_out_data_124; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_125 = pipe6_io_pipe_phv_out_data_125; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_126 = pipe6_io_pipe_phv_out_data_126; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_127 = pipe6_io_pipe_phv_out_data_127; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_128 = pipe6_io_pipe_phv_out_data_128; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_129 = pipe6_io_pipe_phv_out_data_129; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_130 = pipe6_io_pipe_phv_out_data_130; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_131 = pipe6_io_pipe_phv_out_data_131; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_132 = pipe6_io_pipe_phv_out_data_132; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_133 = pipe6_io_pipe_phv_out_data_133; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_134 = pipe6_io_pipe_phv_out_data_134; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_135 = pipe6_io_pipe_phv_out_data_135; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_136 = pipe6_io_pipe_phv_out_data_136; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_137 = pipe6_io_pipe_phv_out_data_137; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_138 = pipe6_io_pipe_phv_out_data_138; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_139 = pipe6_io_pipe_phv_out_data_139; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_140 = pipe6_io_pipe_phv_out_data_140; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_141 = pipe6_io_pipe_phv_out_data_141; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_142 = pipe6_io_pipe_phv_out_data_142; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_143 = pipe6_io_pipe_phv_out_data_143; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_144 = pipe6_io_pipe_phv_out_data_144; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_145 = pipe6_io_pipe_phv_out_data_145; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_146 = pipe6_io_pipe_phv_out_data_146; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_147 = pipe6_io_pipe_phv_out_data_147; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_148 = pipe6_io_pipe_phv_out_data_148; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_149 = pipe6_io_pipe_phv_out_data_149; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_150 = pipe6_io_pipe_phv_out_data_150; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_151 = pipe6_io_pipe_phv_out_data_151; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_152 = pipe6_io_pipe_phv_out_data_152; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_153 = pipe6_io_pipe_phv_out_data_153; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_154 = pipe6_io_pipe_phv_out_data_154; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_155 = pipe6_io_pipe_phv_out_data_155; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_156 = pipe6_io_pipe_phv_out_data_156; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_157 = pipe6_io_pipe_phv_out_data_157; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_158 = pipe6_io_pipe_phv_out_data_158; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_159 = pipe6_io_pipe_phv_out_data_159; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_160 = pipe6_io_pipe_phv_out_data_160; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_161 = pipe6_io_pipe_phv_out_data_161; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_162 = pipe6_io_pipe_phv_out_data_162; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_163 = pipe6_io_pipe_phv_out_data_163; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_164 = pipe6_io_pipe_phv_out_data_164; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_165 = pipe6_io_pipe_phv_out_data_165; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_166 = pipe6_io_pipe_phv_out_data_166; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_167 = pipe6_io_pipe_phv_out_data_167; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_168 = pipe6_io_pipe_phv_out_data_168; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_169 = pipe6_io_pipe_phv_out_data_169; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_170 = pipe6_io_pipe_phv_out_data_170; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_171 = pipe6_io_pipe_phv_out_data_171; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_172 = pipe6_io_pipe_phv_out_data_172; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_173 = pipe6_io_pipe_phv_out_data_173; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_174 = pipe6_io_pipe_phv_out_data_174; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_175 = pipe6_io_pipe_phv_out_data_175; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_176 = pipe6_io_pipe_phv_out_data_176; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_177 = pipe6_io_pipe_phv_out_data_177; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_178 = pipe6_io_pipe_phv_out_data_178; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_179 = pipe6_io_pipe_phv_out_data_179; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_180 = pipe6_io_pipe_phv_out_data_180; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_181 = pipe6_io_pipe_phv_out_data_181; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_182 = pipe6_io_pipe_phv_out_data_182; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_183 = pipe6_io_pipe_phv_out_data_183; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_184 = pipe6_io_pipe_phv_out_data_184; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_185 = pipe6_io_pipe_phv_out_data_185; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_186 = pipe6_io_pipe_phv_out_data_186; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_187 = pipe6_io_pipe_phv_out_data_187; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_188 = pipe6_io_pipe_phv_out_data_188; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_189 = pipe6_io_pipe_phv_out_data_189; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_190 = pipe6_io_pipe_phv_out_data_190; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_191 = pipe6_io_pipe_phv_out_data_191; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_192 = pipe6_io_pipe_phv_out_data_192; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_193 = pipe6_io_pipe_phv_out_data_193; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_194 = pipe6_io_pipe_phv_out_data_194; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_195 = pipe6_io_pipe_phv_out_data_195; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_196 = pipe6_io_pipe_phv_out_data_196; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_197 = pipe6_io_pipe_phv_out_data_197; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_198 = pipe6_io_pipe_phv_out_data_198; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_199 = pipe6_io_pipe_phv_out_data_199; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_200 = pipe6_io_pipe_phv_out_data_200; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_201 = pipe6_io_pipe_phv_out_data_201; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_202 = pipe6_io_pipe_phv_out_data_202; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_203 = pipe6_io_pipe_phv_out_data_203; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_204 = pipe6_io_pipe_phv_out_data_204; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_205 = pipe6_io_pipe_phv_out_data_205; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_206 = pipe6_io_pipe_phv_out_data_206; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_207 = pipe6_io_pipe_phv_out_data_207; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_208 = pipe6_io_pipe_phv_out_data_208; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_209 = pipe6_io_pipe_phv_out_data_209; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_210 = pipe6_io_pipe_phv_out_data_210; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_211 = pipe6_io_pipe_phv_out_data_211; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_212 = pipe6_io_pipe_phv_out_data_212; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_213 = pipe6_io_pipe_phv_out_data_213; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_214 = pipe6_io_pipe_phv_out_data_214; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_215 = pipe6_io_pipe_phv_out_data_215; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_216 = pipe6_io_pipe_phv_out_data_216; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_217 = pipe6_io_pipe_phv_out_data_217; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_218 = pipe6_io_pipe_phv_out_data_218; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_219 = pipe6_io_pipe_phv_out_data_219; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_220 = pipe6_io_pipe_phv_out_data_220; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_221 = pipe6_io_pipe_phv_out_data_221; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_222 = pipe6_io_pipe_phv_out_data_222; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_223 = pipe6_io_pipe_phv_out_data_223; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_224 = pipe6_io_pipe_phv_out_data_224; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_225 = pipe6_io_pipe_phv_out_data_225; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_226 = pipe6_io_pipe_phv_out_data_226; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_227 = pipe6_io_pipe_phv_out_data_227; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_228 = pipe6_io_pipe_phv_out_data_228; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_229 = pipe6_io_pipe_phv_out_data_229; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_230 = pipe6_io_pipe_phv_out_data_230; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_231 = pipe6_io_pipe_phv_out_data_231; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_232 = pipe6_io_pipe_phv_out_data_232; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_233 = pipe6_io_pipe_phv_out_data_233; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_234 = pipe6_io_pipe_phv_out_data_234; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_235 = pipe6_io_pipe_phv_out_data_235; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_236 = pipe6_io_pipe_phv_out_data_236; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_237 = pipe6_io_pipe_phv_out_data_237; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_238 = pipe6_io_pipe_phv_out_data_238; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_239 = pipe6_io_pipe_phv_out_data_239; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_240 = pipe6_io_pipe_phv_out_data_240; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_241 = pipe6_io_pipe_phv_out_data_241; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_242 = pipe6_io_pipe_phv_out_data_242; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_243 = pipe6_io_pipe_phv_out_data_243; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_244 = pipe6_io_pipe_phv_out_data_244; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_245 = pipe6_io_pipe_phv_out_data_245; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_246 = pipe6_io_pipe_phv_out_data_246; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_247 = pipe6_io_pipe_phv_out_data_247; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_248 = pipe6_io_pipe_phv_out_data_248; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_249 = pipe6_io_pipe_phv_out_data_249; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_250 = pipe6_io_pipe_phv_out_data_250; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_251 = pipe6_io_pipe_phv_out_data_251; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_252 = pipe6_io_pipe_phv_out_data_252; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_253 = pipe6_io_pipe_phv_out_data_253; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_254 = pipe6_io_pipe_phv_out_data_254; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_255 = pipe6_io_pipe_phv_out_data_255; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_256 = pipe6_io_pipe_phv_out_data_256; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_257 = pipe6_io_pipe_phv_out_data_257; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_258 = pipe6_io_pipe_phv_out_data_258; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_259 = pipe6_io_pipe_phv_out_data_259; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_260 = pipe6_io_pipe_phv_out_data_260; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_261 = pipe6_io_pipe_phv_out_data_261; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_262 = pipe6_io_pipe_phv_out_data_262; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_263 = pipe6_io_pipe_phv_out_data_263; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_264 = pipe6_io_pipe_phv_out_data_264; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_265 = pipe6_io_pipe_phv_out_data_265; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_266 = pipe6_io_pipe_phv_out_data_266; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_267 = pipe6_io_pipe_phv_out_data_267; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_268 = pipe6_io_pipe_phv_out_data_268; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_269 = pipe6_io_pipe_phv_out_data_269; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_270 = pipe6_io_pipe_phv_out_data_270; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_271 = pipe6_io_pipe_phv_out_data_271; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_272 = pipe6_io_pipe_phv_out_data_272; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_273 = pipe6_io_pipe_phv_out_data_273; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_274 = pipe6_io_pipe_phv_out_data_274; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_275 = pipe6_io_pipe_phv_out_data_275; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_276 = pipe6_io_pipe_phv_out_data_276; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_277 = pipe6_io_pipe_phv_out_data_277; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_278 = pipe6_io_pipe_phv_out_data_278; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_279 = pipe6_io_pipe_phv_out_data_279; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_280 = pipe6_io_pipe_phv_out_data_280; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_281 = pipe6_io_pipe_phv_out_data_281; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_282 = pipe6_io_pipe_phv_out_data_282; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_283 = pipe6_io_pipe_phv_out_data_283; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_284 = pipe6_io_pipe_phv_out_data_284; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_285 = pipe6_io_pipe_phv_out_data_285; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_286 = pipe6_io_pipe_phv_out_data_286; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_287 = pipe6_io_pipe_phv_out_data_287; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_288 = pipe6_io_pipe_phv_out_data_288; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_289 = pipe6_io_pipe_phv_out_data_289; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_290 = pipe6_io_pipe_phv_out_data_290; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_291 = pipe6_io_pipe_phv_out_data_291; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_292 = pipe6_io_pipe_phv_out_data_292; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_293 = pipe6_io_pipe_phv_out_data_293; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_294 = pipe6_io_pipe_phv_out_data_294; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_295 = pipe6_io_pipe_phv_out_data_295; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_296 = pipe6_io_pipe_phv_out_data_296; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_297 = pipe6_io_pipe_phv_out_data_297; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_298 = pipe6_io_pipe_phv_out_data_298; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_299 = pipe6_io_pipe_phv_out_data_299; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_300 = pipe6_io_pipe_phv_out_data_300; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_301 = pipe6_io_pipe_phv_out_data_301; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_302 = pipe6_io_pipe_phv_out_data_302; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_303 = pipe6_io_pipe_phv_out_data_303; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_304 = pipe6_io_pipe_phv_out_data_304; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_305 = pipe6_io_pipe_phv_out_data_305; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_306 = pipe6_io_pipe_phv_out_data_306; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_307 = pipe6_io_pipe_phv_out_data_307; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_308 = pipe6_io_pipe_phv_out_data_308; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_309 = pipe6_io_pipe_phv_out_data_309; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_310 = pipe6_io_pipe_phv_out_data_310; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_311 = pipe6_io_pipe_phv_out_data_311; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_312 = pipe6_io_pipe_phv_out_data_312; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_313 = pipe6_io_pipe_phv_out_data_313; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_314 = pipe6_io_pipe_phv_out_data_314; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_315 = pipe6_io_pipe_phv_out_data_315; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_316 = pipe6_io_pipe_phv_out_data_316; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_317 = pipe6_io_pipe_phv_out_data_317; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_318 = pipe6_io_pipe_phv_out_data_318; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_319 = pipe6_io_pipe_phv_out_data_319; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_320 = pipe6_io_pipe_phv_out_data_320; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_321 = pipe6_io_pipe_phv_out_data_321; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_322 = pipe6_io_pipe_phv_out_data_322; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_323 = pipe6_io_pipe_phv_out_data_323; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_324 = pipe6_io_pipe_phv_out_data_324; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_325 = pipe6_io_pipe_phv_out_data_325; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_326 = pipe6_io_pipe_phv_out_data_326; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_327 = pipe6_io_pipe_phv_out_data_327; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_328 = pipe6_io_pipe_phv_out_data_328; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_329 = pipe6_io_pipe_phv_out_data_329; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_330 = pipe6_io_pipe_phv_out_data_330; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_331 = pipe6_io_pipe_phv_out_data_331; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_332 = pipe6_io_pipe_phv_out_data_332; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_333 = pipe6_io_pipe_phv_out_data_333; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_334 = pipe6_io_pipe_phv_out_data_334; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_335 = pipe6_io_pipe_phv_out_data_335; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_336 = pipe6_io_pipe_phv_out_data_336; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_337 = pipe6_io_pipe_phv_out_data_337; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_338 = pipe6_io_pipe_phv_out_data_338; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_339 = pipe6_io_pipe_phv_out_data_339; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_340 = pipe6_io_pipe_phv_out_data_340; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_341 = pipe6_io_pipe_phv_out_data_341; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_342 = pipe6_io_pipe_phv_out_data_342; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_343 = pipe6_io_pipe_phv_out_data_343; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_344 = pipe6_io_pipe_phv_out_data_344; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_345 = pipe6_io_pipe_phv_out_data_345; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_346 = pipe6_io_pipe_phv_out_data_346; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_347 = pipe6_io_pipe_phv_out_data_347; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_348 = pipe6_io_pipe_phv_out_data_348; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_349 = pipe6_io_pipe_phv_out_data_349; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_350 = pipe6_io_pipe_phv_out_data_350; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_351 = pipe6_io_pipe_phv_out_data_351; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_352 = pipe6_io_pipe_phv_out_data_352; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_353 = pipe6_io_pipe_phv_out_data_353; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_354 = pipe6_io_pipe_phv_out_data_354; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_355 = pipe6_io_pipe_phv_out_data_355; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_356 = pipe6_io_pipe_phv_out_data_356; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_357 = pipe6_io_pipe_phv_out_data_357; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_358 = pipe6_io_pipe_phv_out_data_358; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_359 = pipe6_io_pipe_phv_out_data_359; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_360 = pipe6_io_pipe_phv_out_data_360; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_361 = pipe6_io_pipe_phv_out_data_361; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_362 = pipe6_io_pipe_phv_out_data_362; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_363 = pipe6_io_pipe_phv_out_data_363; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_364 = pipe6_io_pipe_phv_out_data_364; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_365 = pipe6_io_pipe_phv_out_data_365; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_366 = pipe6_io_pipe_phv_out_data_366; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_367 = pipe6_io_pipe_phv_out_data_367; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_368 = pipe6_io_pipe_phv_out_data_368; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_369 = pipe6_io_pipe_phv_out_data_369; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_370 = pipe6_io_pipe_phv_out_data_370; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_371 = pipe6_io_pipe_phv_out_data_371; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_372 = pipe6_io_pipe_phv_out_data_372; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_373 = pipe6_io_pipe_phv_out_data_373; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_374 = pipe6_io_pipe_phv_out_data_374; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_375 = pipe6_io_pipe_phv_out_data_375; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_376 = pipe6_io_pipe_phv_out_data_376; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_377 = pipe6_io_pipe_phv_out_data_377; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_378 = pipe6_io_pipe_phv_out_data_378; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_379 = pipe6_io_pipe_phv_out_data_379; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_380 = pipe6_io_pipe_phv_out_data_380; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_381 = pipe6_io_pipe_phv_out_data_381; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_382 = pipe6_io_pipe_phv_out_data_382; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_383 = pipe6_io_pipe_phv_out_data_383; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_384 = pipe6_io_pipe_phv_out_data_384; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_385 = pipe6_io_pipe_phv_out_data_385; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_386 = pipe6_io_pipe_phv_out_data_386; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_387 = pipe6_io_pipe_phv_out_data_387; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_388 = pipe6_io_pipe_phv_out_data_388; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_389 = pipe6_io_pipe_phv_out_data_389; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_390 = pipe6_io_pipe_phv_out_data_390; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_391 = pipe6_io_pipe_phv_out_data_391; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_392 = pipe6_io_pipe_phv_out_data_392; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_393 = pipe6_io_pipe_phv_out_data_393; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_394 = pipe6_io_pipe_phv_out_data_394; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_395 = pipe6_io_pipe_phv_out_data_395; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_396 = pipe6_io_pipe_phv_out_data_396; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_397 = pipe6_io_pipe_phv_out_data_397; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_398 = pipe6_io_pipe_phv_out_data_398; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_399 = pipe6_io_pipe_phv_out_data_399; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_400 = pipe6_io_pipe_phv_out_data_400; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_401 = pipe6_io_pipe_phv_out_data_401; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_402 = pipe6_io_pipe_phv_out_data_402; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_403 = pipe6_io_pipe_phv_out_data_403; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_404 = pipe6_io_pipe_phv_out_data_404; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_405 = pipe6_io_pipe_phv_out_data_405; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_406 = pipe6_io_pipe_phv_out_data_406; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_407 = pipe6_io_pipe_phv_out_data_407; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_408 = pipe6_io_pipe_phv_out_data_408; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_409 = pipe6_io_pipe_phv_out_data_409; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_410 = pipe6_io_pipe_phv_out_data_410; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_411 = pipe6_io_pipe_phv_out_data_411; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_412 = pipe6_io_pipe_phv_out_data_412; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_413 = pipe6_io_pipe_phv_out_data_413; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_414 = pipe6_io_pipe_phv_out_data_414; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_415 = pipe6_io_pipe_phv_out_data_415; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_416 = pipe6_io_pipe_phv_out_data_416; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_417 = pipe6_io_pipe_phv_out_data_417; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_418 = pipe6_io_pipe_phv_out_data_418; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_419 = pipe6_io_pipe_phv_out_data_419; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_420 = pipe6_io_pipe_phv_out_data_420; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_421 = pipe6_io_pipe_phv_out_data_421; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_422 = pipe6_io_pipe_phv_out_data_422; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_423 = pipe6_io_pipe_phv_out_data_423; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_424 = pipe6_io_pipe_phv_out_data_424; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_425 = pipe6_io_pipe_phv_out_data_425; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_426 = pipe6_io_pipe_phv_out_data_426; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_427 = pipe6_io_pipe_phv_out_data_427; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_428 = pipe6_io_pipe_phv_out_data_428; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_429 = pipe6_io_pipe_phv_out_data_429; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_430 = pipe6_io_pipe_phv_out_data_430; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_431 = pipe6_io_pipe_phv_out_data_431; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_432 = pipe6_io_pipe_phv_out_data_432; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_433 = pipe6_io_pipe_phv_out_data_433; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_434 = pipe6_io_pipe_phv_out_data_434; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_435 = pipe6_io_pipe_phv_out_data_435; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_436 = pipe6_io_pipe_phv_out_data_436; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_437 = pipe6_io_pipe_phv_out_data_437; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_438 = pipe6_io_pipe_phv_out_data_438; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_439 = pipe6_io_pipe_phv_out_data_439; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_440 = pipe6_io_pipe_phv_out_data_440; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_441 = pipe6_io_pipe_phv_out_data_441; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_442 = pipe6_io_pipe_phv_out_data_442; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_443 = pipe6_io_pipe_phv_out_data_443; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_444 = pipe6_io_pipe_phv_out_data_444; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_445 = pipe6_io_pipe_phv_out_data_445; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_446 = pipe6_io_pipe_phv_out_data_446; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_447 = pipe6_io_pipe_phv_out_data_447; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_448 = pipe6_io_pipe_phv_out_data_448; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_449 = pipe6_io_pipe_phv_out_data_449; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_450 = pipe6_io_pipe_phv_out_data_450; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_451 = pipe6_io_pipe_phv_out_data_451; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_452 = pipe6_io_pipe_phv_out_data_452; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_453 = pipe6_io_pipe_phv_out_data_453; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_454 = pipe6_io_pipe_phv_out_data_454; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_455 = pipe6_io_pipe_phv_out_data_455; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_456 = pipe6_io_pipe_phv_out_data_456; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_457 = pipe6_io_pipe_phv_out_data_457; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_458 = pipe6_io_pipe_phv_out_data_458; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_459 = pipe6_io_pipe_phv_out_data_459; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_460 = pipe6_io_pipe_phv_out_data_460; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_461 = pipe6_io_pipe_phv_out_data_461; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_462 = pipe6_io_pipe_phv_out_data_462; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_463 = pipe6_io_pipe_phv_out_data_463; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_464 = pipe6_io_pipe_phv_out_data_464; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_465 = pipe6_io_pipe_phv_out_data_465; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_466 = pipe6_io_pipe_phv_out_data_466; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_467 = pipe6_io_pipe_phv_out_data_467; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_468 = pipe6_io_pipe_phv_out_data_468; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_469 = pipe6_io_pipe_phv_out_data_469; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_470 = pipe6_io_pipe_phv_out_data_470; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_471 = pipe6_io_pipe_phv_out_data_471; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_472 = pipe6_io_pipe_phv_out_data_472; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_473 = pipe6_io_pipe_phv_out_data_473; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_474 = pipe6_io_pipe_phv_out_data_474; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_475 = pipe6_io_pipe_phv_out_data_475; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_476 = pipe6_io_pipe_phv_out_data_476; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_477 = pipe6_io_pipe_phv_out_data_477; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_478 = pipe6_io_pipe_phv_out_data_478; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_479 = pipe6_io_pipe_phv_out_data_479; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_480 = pipe6_io_pipe_phv_out_data_480; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_481 = pipe6_io_pipe_phv_out_data_481; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_482 = pipe6_io_pipe_phv_out_data_482; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_483 = pipe6_io_pipe_phv_out_data_483; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_484 = pipe6_io_pipe_phv_out_data_484; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_485 = pipe6_io_pipe_phv_out_data_485; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_486 = pipe6_io_pipe_phv_out_data_486; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_487 = pipe6_io_pipe_phv_out_data_487; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_488 = pipe6_io_pipe_phv_out_data_488; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_489 = pipe6_io_pipe_phv_out_data_489; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_490 = pipe6_io_pipe_phv_out_data_490; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_491 = pipe6_io_pipe_phv_out_data_491; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_492 = pipe6_io_pipe_phv_out_data_492; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_493 = pipe6_io_pipe_phv_out_data_493; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_494 = pipe6_io_pipe_phv_out_data_494; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_495 = pipe6_io_pipe_phv_out_data_495; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_496 = pipe6_io_pipe_phv_out_data_496; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_497 = pipe6_io_pipe_phv_out_data_497; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_498 = pipe6_io_pipe_phv_out_data_498; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_499 = pipe6_io_pipe_phv_out_data_499; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_500 = pipe6_io_pipe_phv_out_data_500; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_501 = pipe6_io_pipe_phv_out_data_501; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_502 = pipe6_io_pipe_phv_out_data_502; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_503 = pipe6_io_pipe_phv_out_data_503; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_504 = pipe6_io_pipe_phv_out_data_504; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_505 = pipe6_io_pipe_phv_out_data_505; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_506 = pipe6_io_pipe_phv_out_data_506; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_507 = pipe6_io_pipe_phv_out_data_507; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_508 = pipe6_io_pipe_phv_out_data_508; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_509 = pipe6_io_pipe_phv_out_data_509; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_510 = pipe6_io_pipe_phv_out_data_510; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_511 = pipe6_io_pipe_phv_out_data_511; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_0 = pipe6_io_pipe_phv_out_header_0; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_1 = pipe6_io_pipe_phv_out_header_1; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_2 = pipe6_io_pipe_phv_out_header_2; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_3 = pipe6_io_pipe_phv_out_header_3; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_4 = pipe6_io_pipe_phv_out_header_4; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_5 = pipe6_io_pipe_phv_out_header_5; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_6 = pipe6_io_pipe_phv_out_header_6; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_7 = pipe6_io_pipe_phv_out_header_7; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_8 = pipe6_io_pipe_phv_out_header_8; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_9 = pipe6_io_pipe_phv_out_header_9; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_10 = pipe6_io_pipe_phv_out_header_10; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_11 = pipe6_io_pipe_phv_out_header_11; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_12 = pipe6_io_pipe_phv_out_header_12; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_13 = pipe6_io_pipe_phv_out_header_13; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_14 = pipe6_io_pipe_phv_out_header_14; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_15 = pipe6_io_pipe_phv_out_header_15; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_is_valid_processor = pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 164:27]
  assign pipe7_io_hash_depth_0 = hash_depth_0; // @[hash.scala 168:27]
  assign pipe7_io_hash_depth_1 = hash_depth_1; // @[hash.scala 168:27]
  assign pipe7_io_key_in = pipe6_io_key_out; // @[hash.scala 165:27]
  assign pipe7_io_sum_in = pipe6_io_sum_out; // @[hash.scala 166:27]
  assign pipe7_io_val_in = pipe6_io_val_out; // @[hash.scala 167:27]
  assign pipe8_clock = clock;
  assign pipe8_io_pipe_phv_in_data_0 = pipe7_io_pipe_phv_out_data_0; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_1 = pipe7_io_pipe_phv_out_data_1; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_2 = pipe7_io_pipe_phv_out_data_2; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_3 = pipe7_io_pipe_phv_out_data_3; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_4 = pipe7_io_pipe_phv_out_data_4; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_5 = pipe7_io_pipe_phv_out_data_5; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_6 = pipe7_io_pipe_phv_out_data_6; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_7 = pipe7_io_pipe_phv_out_data_7; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_8 = pipe7_io_pipe_phv_out_data_8; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_9 = pipe7_io_pipe_phv_out_data_9; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_10 = pipe7_io_pipe_phv_out_data_10; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_11 = pipe7_io_pipe_phv_out_data_11; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_12 = pipe7_io_pipe_phv_out_data_12; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_13 = pipe7_io_pipe_phv_out_data_13; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_14 = pipe7_io_pipe_phv_out_data_14; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_15 = pipe7_io_pipe_phv_out_data_15; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_16 = pipe7_io_pipe_phv_out_data_16; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_17 = pipe7_io_pipe_phv_out_data_17; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_18 = pipe7_io_pipe_phv_out_data_18; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_19 = pipe7_io_pipe_phv_out_data_19; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_20 = pipe7_io_pipe_phv_out_data_20; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_21 = pipe7_io_pipe_phv_out_data_21; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_22 = pipe7_io_pipe_phv_out_data_22; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_23 = pipe7_io_pipe_phv_out_data_23; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_24 = pipe7_io_pipe_phv_out_data_24; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_25 = pipe7_io_pipe_phv_out_data_25; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_26 = pipe7_io_pipe_phv_out_data_26; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_27 = pipe7_io_pipe_phv_out_data_27; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_28 = pipe7_io_pipe_phv_out_data_28; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_29 = pipe7_io_pipe_phv_out_data_29; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_30 = pipe7_io_pipe_phv_out_data_30; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_31 = pipe7_io_pipe_phv_out_data_31; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_32 = pipe7_io_pipe_phv_out_data_32; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_33 = pipe7_io_pipe_phv_out_data_33; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_34 = pipe7_io_pipe_phv_out_data_34; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_35 = pipe7_io_pipe_phv_out_data_35; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_36 = pipe7_io_pipe_phv_out_data_36; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_37 = pipe7_io_pipe_phv_out_data_37; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_38 = pipe7_io_pipe_phv_out_data_38; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_39 = pipe7_io_pipe_phv_out_data_39; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_40 = pipe7_io_pipe_phv_out_data_40; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_41 = pipe7_io_pipe_phv_out_data_41; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_42 = pipe7_io_pipe_phv_out_data_42; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_43 = pipe7_io_pipe_phv_out_data_43; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_44 = pipe7_io_pipe_phv_out_data_44; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_45 = pipe7_io_pipe_phv_out_data_45; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_46 = pipe7_io_pipe_phv_out_data_46; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_47 = pipe7_io_pipe_phv_out_data_47; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_48 = pipe7_io_pipe_phv_out_data_48; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_49 = pipe7_io_pipe_phv_out_data_49; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_50 = pipe7_io_pipe_phv_out_data_50; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_51 = pipe7_io_pipe_phv_out_data_51; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_52 = pipe7_io_pipe_phv_out_data_52; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_53 = pipe7_io_pipe_phv_out_data_53; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_54 = pipe7_io_pipe_phv_out_data_54; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_55 = pipe7_io_pipe_phv_out_data_55; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_56 = pipe7_io_pipe_phv_out_data_56; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_57 = pipe7_io_pipe_phv_out_data_57; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_58 = pipe7_io_pipe_phv_out_data_58; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_59 = pipe7_io_pipe_phv_out_data_59; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_60 = pipe7_io_pipe_phv_out_data_60; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_61 = pipe7_io_pipe_phv_out_data_61; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_62 = pipe7_io_pipe_phv_out_data_62; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_63 = pipe7_io_pipe_phv_out_data_63; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_64 = pipe7_io_pipe_phv_out_data_64; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_65 = pipe7_io_pipe_phv_out_data_65; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_66 = pipe7_io_pipe_phv_out_data_66; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_67 = pipe7_io_pipe_phv_out_data_67; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_68 = pipe7_io_pipe_phv_out_data_68; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_69 = pipe7_io_pipe_phv_out_data_69; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_70 = pipe7_io_pipe_phv_out_data_70; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_71 = pipe7_io_pipe_phv_out_data_71; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_72 = pipe7_io_pipe_phv_out_data_72; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_73 = pipe7_io_pipe_phv_out_data_73; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_74 = pipe7_io_pipe_phv_out_data_74; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_75 = pipe7_io_pipe_phv_out_data_75; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_76 = pipe7_io_pipe_phv_out_data_76; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_77 = pipe7_io_pipe_phv_out_data_77; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_78 = pipe7_io_pipe_phv_out_data_78; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_79 = pipe7_io_pipe_phv_out_data_79; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_80 = pipe7_io_pipe_phv_out_data_80; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_81 = pipe7_io_pipe_phv_out_data_81; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_82 = pipe7_io_pipe_phv_out_data_82; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_83 = pipe7_io_pipe_phv_out_data_83; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_84 = pipe7_io_pipe_phv_out_data_84; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_85 = pipe7_io_pipe_phv_out_data_85; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_86 = pipe7_io_pipe_phv_out_data_86; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_87 = pipe7_io_pipe_phv_out_data_87; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_88 = pipe7_io_pipe_phv_out_data_88; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_89 = pipe7_io_pipe_phv_out_data_89; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_90 = pipe7_io_pipe_phv_out_data_90; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_91 = pipe7_io_pipe_phv_out_data_91; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_92 = pipe7_io_pipe_phv_out_data_92; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_93 = pipe7_io_pipe_phv_out_data_93; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_94 = pipe7_io_pipe_phv_out_data_94; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_95 = pipe7_io_pipe_phv_out_data_95; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_96 = pipe7_io_pipe_phv_out_data_96; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_97 = pipe7_io_pipe_phv_out_data_97; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_98 = pipe7_io_pipe_phv_out_data_98; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_99 = pipe7_io_pipe_phv_out_data_99; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_100 = pipe7_io_pipe_phv_out_data_100; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_101 = pipe7_io_pipe_phv_out_data_101; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_102 = pipe7_io_pipe_phv_out_data_102; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_103 = pipe7_io_pipe_phv_out_data_103; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_104 = pipe7_io_pipe_phv_out_data_104; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_105 = pipe7_io_pipe_phv_out_data_105; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_106 = pipe7_io_pipe_phv_out_data_106; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_107 = pipe7_io_pipe_phv_out_data_107; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_108 = pipe7_io_pipe_phv_out_data_108; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_109 = pipe7_io_pipe_phv_out_data_109; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_110 = pipe7_io_pipe_phv_out_data_110; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_111 = pipe7_io_pipe_phv_out_data_111; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_112 = pipe7_io_pipe_phv_out_data_112; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_113 = pipe7_io_pipe_phv_out_data_113; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_114 = pipe7_io_pipe_phv_out_data_114; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_115 = pipe7_io_pipe_phv_out_data_115; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_116 = pipe7_io_pipe_phv_out_data_116; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_117 = pipe7_io_pipe_phv_out_data_117; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_118 = pipe7_io_pipe_phv_out_data_118; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_119 = pipe7_io_pipe_phv_out_data_119; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_120 = pipe7_io_pipe_phv_out_data_120; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_121 = pipe7_io_pipe_phv_out_data_121; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_122 = pipe7_io_pipe_phv_out_data_122; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_123 = pipe7_io_pipe_phv_out_data_123; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_124 = pipe7_io_pipe_phv_out_data_124; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_125 = pipe7_io_pipe_phv_out_data_125; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_126 = pipe7_io_pipe_phv_out_data_126; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_127 = pipe7_io_pipe_phv_out_data_127; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_128 = pipe7_io_pipe_phv_out_data_128; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_129 = pipe7_io_pipe_phv_out_data_129; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_130 = pipe7_io_pipe_phv_out_data_130; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_131 = pipe7_io_pipe_phv_out_data_131; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_132 = pipe7_io_pipe_phv_out_data_132; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_133 = pipe7_io_pipe_phv_out_data_133; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_134 = pipe7_io_pipe_phv_out_data_134; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_135 = pipe7_io_pipe_phv_out_data_135; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_136 = pipe7_io_pipe_phv_out_data_136; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_137 = pipe7_io_pipe_phv_out_data_137; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_138 = pipe7_io_pipe_phv_out_data_138; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_139 = pipe7_io_pipe_phv_out_data_139; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_140 = pipe7_io_pipe_phv_out_data_140; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_141 = pipe7_io_pipe_phv_out_data_141; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_142 = pipe7_io_pipe_phv_out_data_142; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_143 = pipe7_io_pipe_phv_out_data_143; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_144 = pipe7_io_pipe_phv_out_data_144; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_145 = pipe7_io_pipe_phv_out_data_145; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_146 = pipe7_io_pipe_phv_out_data_146; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_147 = pipe7_io_pipe_phv_out_data_147; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_148 = pipe7_io_pipe_phv_out_data_148; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_149 = pipe7_io_pipe_phv_out_data_149; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_150 = pipe7_io_pipe_phv_out_data_150; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_151 = pipe7_io_pipe_phv_out_data_151; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_152 = pipe7_io_pipe_phv_out_data_152; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_153 = pipe7_io_pipe_phv_out_data_153; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_154 = pipe7_io_pipe_phv_out_data_154; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_155 = pipe7_io_pipe_phv_out_data_155; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_156 = pipe7_io_pipe_phv_out_data_156; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_157 = pipe7_io_pipe_phv_out_data_157; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_158 = pipe7_io_pipe_phv_out_data_158; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_159 = pipe7_io_pipe_phv_out_data_159; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_160 = pipe7_io_pipe_phv_out_data_160; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_161 = pipe7_io_pipe_phv_out_data_161; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_162 = pipe7_io_pipe_phv_out_data_162; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_163 = pipe7_io_pipe_phv_out_data_163; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_164 = pipe7_io_pipe_phv_out_data_164; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_165 = pipe7_io_pipe_phv_out_data_165; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_166 = pipe7_io_pipe_phv_out_data_166; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_167 = pipe7_io_pipe_phv_out_data_167; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_168 = pipe7_io_pipe_phv_out_data_168; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_169 = pipe7_io_pipe_phv_out_data_169; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_170 = pipe7_io_pipe_phv_out_data_170; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_171 = pipe7_io_pipe_phv_out_data_171; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_172 = pipe7_io_pipe_phv_out_data_172; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_173 = pipe7_io_pipe_phv_out_data_173; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_174 = pipe7_io_pipe_phv_out_data_174; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_175 = pipe7_io_pipe_phv_out_data_175; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_176 = pipe7_io_pipe_phv_out_data_176; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_177 = pipe7_io_pipe_phv_out_data_177; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_178 = pipe7_io_pipe_phv_out_data_178; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_179 = pipe7_io_pipe_phv_out_data_179; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_180 = pipe7_io_pipe_phv_out_data_180; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_181 = pipe7_io_pipe_phv_out_data_181; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_182 = pipe7_io_pipe_phv_out_data_182; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_183 = pipe7_io_pipe_phv_out_data_183; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_184 = pipe7_io_pipe_phv_out_data_184; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_185 = pipe7_io_pipe_phv_out_data_185; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_186 = pipe7_io_pipe_phv_out_data_186; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_187 = pipe7_io_pipe_phv_out_data_187; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_188 = pipe7_io_pipe_phv_out_data_188; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_189 = pipe7_io_pipe_phv_out_data_189; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_190 = pipe7_io_pipe_phv_out_data_190; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_191 = pipe7_io_pipe_phv_out_data_191; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_192 = pipe7_io_pipe_phv_out_data_192; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_193 = pipe7_io_pipe_phv_out_data_193; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_194 = pipe7_io_pipe_phv_out_data_194; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_195 = pipe7_io_pipe_phv_out_data_195; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_196 = pipe7_io_pipe_phv_out_data_196; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_197 = pipe7_io_pipe_phv_out_data_197; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_198 = pipe7_io_pipe_phv_out_data_198; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_199 = pipe7_io_pipe_phv_out_data_199; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_200 = pipe7_io_pipe_phv_out_data_200; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_201 = pipe7_io_pipe_phv_out_data_201; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_202 = pipe7_io_pipe_phv_out_data_202; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_203 = pipe7_io_pipe_phv_out_data_203; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_204 = pipe7_io_pipe_phv_out_data_204; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_205 = pipe7_io_pipe_phv_out_data_205; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_206 = pipe7_io_pipe_phv_out_data_206; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_207 = pipe7_io_pipe_phv_out_data_207; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_208 = pipe7_io_pipe_phv_out_data_208; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_209 = pipe7_io_pipe_phv_out_data_209; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_210 = pipe7_io_pipe_phv_out_data_210; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_211 = pipe7_io_pipe_phv_out_data_211; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_212 = pipe7_io_pipe_phv_out_data_212; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_213 = pipe7_io_pipe_phv_out_data_213; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_214 = pipe7_io_pipe_phv_out_data_214; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_215 = pipe7_io_pipe_phv_out_data_215; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_216 = pipe7_io_pipe_phv_out_data_216; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_217 = pipe7_io_pipe_phv_out_data_217; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_218 = pipe7_io_pipe_phv_out_data_218; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_219 = pipe7_io_pipe_phv_out_data_219; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_220 = pipe7_io_pipe_phv_out_data_220; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_221 = pipe7_io_pipe_phv_out_data_221; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_222 = pipe7_io_pipe_phv_out_data_222; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_223 = pipe7_io_pipe_phv_out_data_223; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_224 = pipe7_io_pipe_phv_out_data_224; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_225 = pipe7_io_pipe_phv_out_data_225; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_226 = pipe7_io_pipe_phv_out_data_226; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_227 = pipe7_io_pipe_phv_out_data_227; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_228 = pipe7_io_pipe_phv_out_data_228; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_229 = pipe7_io_pipe_phv_out_data_229; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_230 = pipe7_io_pipe_phv_out_data_230; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_231 = pipe7_io_pipe_phv_out_data_231; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_232 = pipe7_io_pipe_phv_out_data_232; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_233 = pipe7_io_pipe_phv_out_data_233; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_234 = pipe7_io_pipe_phv_out_data_234; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_235 = pipe7_io_pipe_phv_out_data_235; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_236 = pipe7_io_pipe_phv_out_data_236; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_237 = pipe7_io_pipe_phv_out_data_237; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_238 = pipe7_io_pipe_phv_out_data_238; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_239 = pipe7_io_pipe_phv_out_data_239; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_240 = pipe7_io_pipe_phv_out_data_240; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_241 = pipe7_io_pipe_phv_out_data_241; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_242 = pipe7_io_pipe_phv_out_data_242; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_243 = pipe7_io_pipe_phv_out_data_243; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_244 = pipe7_io_pipe_phv_out_data_244; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_245 = pipe7_io_pipe_phv_out_data_245; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_246 = pipe7_io_pipe_phv_out_data_246; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_247 = pipe7_io_pipe_phv_out_data_247; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_248 = pipe7_io_pipe_phv_out_data_248; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_249 = pipe7_io_pipe_phv_out_data_249; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_250 = pipe7_io_pipe_phv_out_data_250; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_251 = pipe7_io_pipe_phv_out_data_251; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_252 = pipe7_io_pipe_phv_out_data_252; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_253 = pipe7_io_pipe_phv_out_data_253; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_254 = pipe7_io_pipe_phv_out_data_254; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_255 = pipe7_io_pipe_phv_out_data_255; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_256 = pipe7_io_pipe_phv_out_data_256; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_257 = pipe7_io_pipe_phv_out_data_257; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_258 = pipe7_io_pipe_phv_out_data_258; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_259 = pipe7_io_pipe_phv_out_data_259; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_260 = pipe7_io_pipe_phv_out_data_260; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_261 = pipe7_io_pipe_phv_out_data_261; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_262 = pipe7_io_pipe_phv_out_data_262; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_263 = pipe7_io_pipe_phv_out_data_263; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_264 = pipe7_io_pipe_phv_out_data_264; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_265 = pipe7_io_pipe_phv_out_data_265; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_266 = pipe7_io_pipe_phv_out_data_266; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_267 = pipe7_io_pipe_phv_out_data_267; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_268 = pipe7_io_pipe_phv_out_data_268; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_269 = pipe7_io_pipe_phv_out_data_269; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_270 = pipe7_io_pipe_phv_out_data_270; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_271 = pipe7_io_pipe_phv_out_data_271; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_272 = pipe7_io_pipe_phv_out_data_272; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_273 = pipe7_io_pipe_phv_out_data_273; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_274 = pipe7_io_pipe_phv_out_data_274; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_275 = pipe7_io_pipe_phv_out_data_275; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_276 = pipe7_io_pipe_phv_out_data_276; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_277 = pipe7_io_pipe_phv_out_data_277; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_278 = pipe7_io_pipe_phv_out_data_278; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_279 = pipe7_io_pipe_phv_out_data_279; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_280 = pipe7_io_pipe_phv_out_data_280; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_281 = pipe7_io_pipe_phv_out_data_281; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_282 = pipe7_io_pipe_phv_out_data_282; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_283 = pipe7_io_pipe_phv_out_data_283; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_284 = pipe7_io_pipe_phv_out_data_284; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_285 = pipe7_io_pipe_phv_out_data_285; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_286 = pipe7_io_pipe_phv_out_data_286; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_287 = pipe7_io_pipe_phv_out_data_287; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_288 = pipe7_io_pipe_phv_out_data_288; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_289 = pipe7_io_pipe_phv_out_data_289; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_290 = pipe7_io_pipe_phv_out_data_290; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_291 = pipe7_io_pipe_phv_out_data_291; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_292 = pipe7_io_pipe_phv_out_data_292; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_293 = pipe7_io_pipe_phv_out_data_293; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_294 = pipe7_io_pipe_phv_out_data_294; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_295 = pipe7_io_pipe_phv_out_data_295; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_296 = pipe7_io_pipe_phv_out_data_296; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_297 = pipe7_io_pipe_phv_out_data_297; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_298 = pipe7_io_pipe_phv_out_data_298; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_299 = pipe7_io_pipe_phv_out_data_299; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_300 = pipe7_io_pipe_phv_out_data_300; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_301 = pipe7_io_pipe_phv_out_data_301; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_302 = pipe7_io_pipe_phv_out_data_302; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_303 = pipe7_io_pipe_phv_out_data_303; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_304 = pipe7_io_pipe_phv_out_data_304; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_305 = pipe7_io_pipe_phv_out_data_305; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_306 = pipe7_io_pipe_phv_out_data_306; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_307 = pipe7_io_pipe_phv_out_data_307; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_308 = pipe7_io_pipe_phv_out_data_308; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_309 = pipe7_io_pipe_phv_out_data_309; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_310 = pipe7_io_pipe_phv_out_data_310; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_311 = pipe7_io_pipe_phv_out_data_311; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_312 = pipe7_io_pipe_phv_out_data_312; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_313 = pipe7_io_pipe_phv_out_data_313; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_314 = pipe7_io_pipe_phv_out_data_314; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_315 = pipe7_io_pipe_phv_out_data_315; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_316 = pipe7_io_pipe_phv_out_data_316; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_317 = pipe7_io_pipe_phv_out_data_317; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_318 = pipe7_io_pipe_phv_out_data_318; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_319 = pipe7_io_pipe_phv_out_data_319; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_320 = pipe7_io_pipe_phv_out_data_320; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_321 = pipe7_io_pipe_phv_out_data_321; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_322 = pipe7_io_pipe_phv_out_data_322; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_323 = pipe7_io_pipe_phv_out_data_323; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_324 = pipe7_io_pipe_phv_out_data_324; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_325 = pipe7_io_pipe_phv_out_data_325; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_326 = pipe7_io_pipe_phv_out_data_326; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_327 = pipe7_io_pipe_phv_out_data_327; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_328 = pipe7_io_pipe_phv_out_data_328; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_329 = pipe7_io_pipe_phv_out_data_329; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_330 = pipe7_io_pipe_phv_out_data_330; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_331 = pipe7_io_pipe_phv_out_data_331; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_332 = pipe7_io_pipe_phv_out_data_332; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_333 = pipe7_io_pipe_phv_out_data_333; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_334 = pipe7_io_pipe_phv_out_data_334; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_335 = pipe7_io_pipe_phv_out_data_335; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_336 = pipe7_io_pipe_phv_out_data_336; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_337 = pipe7_io_pipe_phv_out_data_337; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_338 = pipe7_io_pipe_phv_out_data_338; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_339 = pipe7_io_pipe_phv_out_data_339; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_340 = pipe7_io_pipe_phv_out_data_340; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_341 = pipe7_io_pipe_phv_out_data_341; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_342 = pipe7_io_pipe_phv_out_data_342; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_343 = pipe7_io_pipe_phv_out_data_343; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_344 = pipe7_io_pipe_phv_out_data_344; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_345 = pipe7_io_pipe_phv_out_data_345; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_346 = pipe7_io_pipe_phv_out_data_346; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_347 = pipe7_io_pipe_phv_out_data_347; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_348 = pipe7_io_pipe_phv_out_data_348; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_349 = pipe7_io_pipe_phv_out_data_349; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_350 = pipe7_io_pipe_phv_out_data_350; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_351 = pipe7_io_pipe_phv_out_data_351; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_352 = pipe7_io_pipe_phv_out_data_352; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_353 = pipe7_io_pipe_phv_out_data_353; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_354 = pipe7_io_pipe_phv_out_data_354; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_355 = pipe7_io_pipe_phv_out_data_355; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_356 = pipe7_io_pipe_phv_out_data_356; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_357 = pipe7_io_pipe_phv_out_data_357; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_358 = pipe7_io_pipe_phv_out_data_358; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_359 = pipe7_io_pipe_phv_out_data_359; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_360 = pipe7_io_pipe_phv_out_data_360; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_361 = pipe7_io_pipe_phv_out_data_361; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_362 = pipe7_io_pipe_phv_out_data_362; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_363 = pipe7_io_pipe_phv_out_data_363; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_364 = pipe7_io_pipe_phv_out_data_364; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_365 = pipe7_io_pipe_phv_out_data_365; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_366 = pipe7_io_pipe_phv_out_data_366; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_367 = pipe7_io_pipe_phv_out_data_367; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_368 = pipe7_io_pipe_phv_out_data_368; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_369 = pipe7_io_pipe_phv_out_data_369; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_370 = pipe7_io_pipe_phv_out_data_370; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_371 = pipe7_io_pipe_phv_out_data_371; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_372 = pipe7_io_pipe_phv_out_data_372; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_373 = pipe7_io_pipe_phv_out_data_373; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_374 = pipe7_io_pipe_phv_out_data_374; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_375 = pipe7_io_pipe_phv_out_data_375; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_376 = pipe7_io_pipe_phv_out_data_376; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_377 = pipe7_io_pipe_phv_out_data_377; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_378 = pipe7_io_pipe_phv_out_data_378; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_379 = pipe7_io_pipe_phv_out_data_379; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_380 = pipe7_io_pipe_phv_out_data_380; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_381 = pipe7_io_pipe_phv_out_data_381; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_382 = pipe7_io_pipe_phv_out_data_382; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_383 = pipe7_io_pipe_phv_out_data_383; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_384 = pipe7_io_pipe_phv_out_data_384; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_385 = pipe7_io_pipe_phv_out_data_385; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_386 = pipe7_io_pipe_phv_out_data_386; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_387 = pipe7_io_pipe_phv_out_data_387; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_388 = pipe7_io_pipe_phv_out_data_388; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_389 = pipe7_io_pipe_phv_out_data_389; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_390 = pipe7_io_pipe_phv_out_data_390; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_391 = pipe7_io_pipe_phv_out_data_391; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_392 = pipe7_io_pipe_phv_out_data_392; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_393 = pipe7_io_pipe_phv_out_data_393; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_394 = pipe7_io_pipe_phv_out_data_394; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_395 = pipe7_io_pipe_phv_out_data_395; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_396 = pipe7_io_pipe_phv_out_data_396; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_397 = pipe7_io_pipe_phv_out_data_397; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_398 = pipe7_io_pipe_phv_out_data_398; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_399 = pipe7_io_pipe_phv_out_data_399; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_400 = pipe7_io_pipe_phv_out_data_400; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_401 = pipe7_io_pipe_phv_out_data_401; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_402 = pipe7_io_pipe_phv_out_data_402; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_403 = pipe7_io_pipe_phv_out_data_403; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_404 = pipe7_io_pipe_phv_out_data_404; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_405 = pipe7_io_pipe_phv_out_data_405; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_406 = pipe7_io_pipe_phv_out_data_406; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_407 = pipe7_io_pipe_phv_out_data_407; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_408 = pipe7_io_pipe_phv_out_data_408; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_409 = pipe7_io_pipe_phv_out_data_409; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_410 = pipe7_io_pipe_phv_out_data_410; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_411 = pipe7_io_pipe_phv_out_data_411; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_412 = pipe7_io_pipe_phv_out_data_412; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_413 = pipe7_io_pipe_phv_out_data_413; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_414 = pipe7_io_pipe_phv_out_data_414; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_415 = pipe7_io_pipe_phv_out_data_415; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_416 = pipe7_io_pipe_phv_out_data_416; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_417 = pipe7_io_pipe_phv_out_data_417; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_418 = pipe7_io_pipe_phv_out_data_418; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_419 = pipe7_io_pipe_phv_out_data_419; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_420 = pipe7_io_pipe_phv_out_data_420; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_421 = pipe7_io_pipe_phv_out_data_421; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_422 = pipe7_io_pipe_phv_out_data_422; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_423 = pipe7_io_pipe_phv_out_data_423; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_424 = pipe7_io_pipe_phv_out_data_424; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_425 = pipe7_io_pipe_phv_out_data_425; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_426 = pipe7_io_pipe_phv_out_data_426; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_427 = pipe7_io_pipe_phv_out_data_427; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_428 = pipe7_io_pipe_phv_out_data_428; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_429 = pipe7_io_pipe_phv_out_data_429; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_430 = pipe7_io_pipe_phv_out_data_430; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_431 = pipe7_io_pipe_phv_out_data_431; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_432 = pipe7_io_pipe_phv_out_data_432; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_433 = pipe7_io_pipe_phv_out_data_433; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_434 = pipe7_io_pipe_phv_out_data_434; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_435 = pipe7_io_pipe_phv_out_data_435; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_436 = pipe7_io_pipe_phv_out_data_436; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_437 = pipe7_io_pipe_phv_out_data_437; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_438 = pipe7_io_pipe_phv_out_data_438; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_439 = pipe7_io_pipe_phv_out_data_439; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_440 = pipe7_io_pipe_phv_out_data_440; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_441 = pipe7_io_pipe_phv_out_data_441; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_442 = pipe7_io_pipe_phv_out_data_442; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_443 = pipe7_io_pipe_phv_out_data_443; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_444 = pipe7_io_pipe_phv_out_data_444; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_445 = pipe7_io_pipe_phv_out_data_445; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_446 = pipe7_io_pipe_phv_out_data_446; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_447 = pipe7_io_pipe_phv_out_data_447; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_448 = pipe7_io_pipe_phv_out_data_448; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_449 = pipe7_io_pipe_phv_out_data_449; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_450 = pipe7_io_pipe_phv_out_data_450; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_451 = pipe7_io_pipe_phv_out_data_451; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_452 = pipe7_io_pipe_phv_out_data_452; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_453 = pipe7_io_pipe_phv_out_data_453; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_454 = pipe7_io_pipe_phv_out_data_454; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_455 = pipe7_io_pipe_phv_out_data_455; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_456 = pipe7_io_pipe_phv_out_data_456; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_457 = pipe7_io_pipe_phv_out_data_457; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_458 = pipe7_io_pipe_phv_out_data_458; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_459 = pipe7_io_pipe_phv_out_data_459; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_460 = pipe7_io_pipe_phv_out_data_460; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_461 = pipe7_io_pipe_phv_out_data_461; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_462 = pipe7_io_pipe_phv_out_data_462; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_463 = pipe7_io_pipe_phv_out_data_463; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_464 = pipe7_io_pipe_phv_out_data_464; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_465 = pipe7_io_pipe_phv_out_data_465; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_466 = pipe7_io_pipe_phv_out_data_466; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_467 = pipe7_io_pipe_phv_out_data_467; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_468 = pipe7_io_pipe_phv_out_data_468; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_469 = pipe7_io_pipe_phv_out_data_469; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_470 = pipe7_io_pipe_phv_out_data_470; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_471 = pipe7_io_pipe_phv_out_data_471; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_472 = pipe7_io_pipe_phv_out_data_472; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_473 = pipe7_io_pipe_phv_out_data_473; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_474 = pipe7_io_pipe_phv_out_data_474; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_475 = pipe7_io_pipe_phv_out_data_475; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_476 = pipe7_io_pipe_phv_out_data_476; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_477 = pipe7_io_pipe_phv_out_data_477; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_478 = pipe7_io_pipe_phv_out_data_478; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_479 = pipe7_io_pipe_phv_out_data_479; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_480 = pipe7_io_pipe_phv_out_data_480; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_481 = pipe7_io_pipe_phv_out_data_481; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_482 = pipe7_io_pipe_phv_out_data_482; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_483 = pipe7_io_pipe_phv_out_data_483; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_484 = pipe7_io_pipe_phv_out_data_484; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_485 = pipe7_io_pipe_phv_out_data_485; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_486 = pipe7_io_pipe_phv_out_data_486; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_487 = pipe7_io_pipe_phv_out_data_487; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_488 = pipe7_io_pipe_phv_out_data_488; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_489 = pipe7_io_pipe_phv_out_data_489; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_490 = pipe7_io_pipe_phv_out_data_490; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_491 = pipe7_io_pipe_phv_out_data_491; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_492 = pipe7_io_pipe_phv_out_data_492; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_493 = pipe7_io_pipe_phv_out_data_493; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_494 = pipe7_io_pipe_phv_out_data_494; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_495 = pipe7_io_pipe_phv_out_data_495; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_496 = pipe7_io_pipe_phv_out_data_496; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_497 = pipe7_io_pipe_phv_out_data_497; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_498 = pipe7_io_pipe_phv_out_data_498; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_499 = pipe7_io_pipe_phv_out_data_499; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_500 = pipe7_io_pipe_phv_out_data_500; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_501 = pipe7_io_pipe_phv_out_data_501; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_502 = pipe7_io_pipe_phv_out_data_502; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_503 = pipe7_io_pipe_phv_out_data_503; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_504 = pipe7_io_pipe_phv_out_data_504; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_505 = pipe7_io_pipe_phv_out_data_505; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_506 = pipe7_io_pipe_phv_out_data_506; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_507 = pipe7_io_pipe_phv_out_data_507; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_508 = pipe7_io_pipe_phv_out_data_508; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_509 = pipe7_io_pipe_phv_out_data_509; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_510 = pipe7_io_pipe_phv_out_data_510; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_511 = pipe7_io_pipe_phv_out_data_511; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_0 = pipe7_io_pipe_phv_out_header_0; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_1 = pipe7_io_pipe_phv_out_header_1; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_2 = pipe7_io_pipe_phv_out_header_2; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_3 = pipe7_io_pipe_phv_out_header_3; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_4 = pipe7_io_pipe_phv_out_header_4; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_5 = pipe7_io_pipe_phv_out_header_5; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_6 = pipe7_io_pipe_phv_out_header_6; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_7 = pipe7_io_pipe_phv_out_header_7; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_8 = pipe7_io_pipe_phv_out_header_8; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_9 = pipe7_io_pipe_phv_out_header_9; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_10 = pipe7_io_pipe_phv_out_header_10; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_11 = pipe7_io_pipe_phv_out_header_11; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_12 = pipe7_io_pipe_phv_out_header_12; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_13 = pipe7_io_pipe_phv_out_header_13; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_14 = pipe7_io_pipe_phv_out_header_14; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_15 = pipe7_io_pipe_phv_out_header_15; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_current_state = pipe7_io_pipe_phv_out_parse_current_state; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_current_offset = pipe7_io_pipe_phv_out_parse_current_offset; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_transition_field = pipe7_io_pipe_phv_out_parse_transition_field; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_next_processor_id = pipe7_io_pipe_phv_out_next_processor_id; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_next_config_id = pipe7_io_pipe_phv_out_next_config_id; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_is_valid_processor = pipe7_io_pipe_phv_out_is_valid_processor; // @[hash.scala 170:27]
  assign pipe8_io_hash_depth_0 = hash_depth_0; // @[hash.scala 174:27]
  assign pipe8_io_hash_depth_1 = hash_depth_1; // @[hash.scala 174:27]
  assign pipe8_io_key_in = pipe7_io_key_out; // @[hash.scala 171:27]
  assign pipe8_io_sum_in = pipe7_io_sum_out; // @[hash.scala 172:27]
  assign pipe8_io_val_in = pipe7_io_val_out; // @[hash.scala 173:27]
  always @(posedge clock) begin
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (~io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_0 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_1 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hash_depth_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  hash_depth_1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
