module PrimitiveWriteBack(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [31:0] io_vliw_in_4,
  input  [31:0] io_vliw_in_5,
  input  [31:0] io_vliw_in_6,
  input  [31:0] io_vliw_in_7,
  input  [31:0] io_field_in_0,
  input  [31:0] io_field_in_1,
  input  [31:0] io_field_in_2,
  input  [31:0] io_field_in_3,
  input  [31:0] io_field_in_4,
  input  [31:0] io_field_in_5,
  input  [31:0] io_field_in_6,
  input  [31:0] io_field_in_7,
  input  [3:0]  io_mask_in_0,
  input  [3:0]  io_mask_in_1,
  input  [3:0]  io_mask_in_2,
  input  [3:0]  io_mask_in_3,
  input  [3:0]  io_mask_in_4,
  input  [3:0]  io_mask_in_5,
  input  [3:0]  io_mask_in_6,
  input  [3:0]  io_mask_in_7,
  input  [5:0]  io_dst_offset_in_0,
  input  [5:0]  io_dst_offset_in_1,
  input  [5:0]  io_dst_offset_in_2,
  input  [5:0]  io_dst_offset_in_3,
  input  [5:0]  io_dst_offset_in_4,
  input  [5:0]  io_dst_offset_in_5,
  input  [5:0]  io_dst_offset_in_6,
  input  [5:0]  io_dst_offset_in_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 448:22]
  reg [7:0] phv_data_1; // @[executor.scala 448:22]
  reg [7:0] phv_data_2; // @[executor.scala 448:22]
  reg [7:0] phv_data_3; // @[executor.scala 448:22]
  reg [7:0] phv_data_4; // @[executor.scala 448:22]
  reg [7:0] phv_data_5; // @[executor.scala 448:22]
  reg [7:0] phv_data_6; // @[executor.scala 448:22]
  reg [7:0] phv_data_7; // @[executor.scala 448:22]
  reg [7:0] phv_data_8; // @[executor.scala 448:22]
  reg [7:0] phv_data_9; // @[executor.scala 448:22]
  reg [7:0] phv_data_10; // @[executor.scala 448:22]
  reg [7:0] phv_data_11; // @[executor.scala 448:22]
  reg [7:0] phv_data_12; // @[executor.scala 448:22]
  reg [7:0] phv_data_13; // @[executor.scala 448:22]
  reg [7:0] phv_data_14; // @[executor.scala 448:22]
  reg [7:0] phv_data_15; // @[executor.scala 448:22]
  reg [7:0] phv_data_16; // @[executor.scala 448:22]
  reg [7:0] phv_data_17; // @[executor.scala 448:22]
  reg [7:0] phv_data_18; // @[executor.scala 448:22]
  reg [7:0] phv_data_19; // @[executor.scala 448:22]
  reg [7:0] phv_data_20; // @[executor.scala 448:22]
  reg [7:0] phv_data_21; // @[executor.scala 448:22]
  reg [7:0] phv_data_22; // @[executor.scala 448:22]
  reg [7:0] phv_data_23; // @[executor.scala 448:22]
  reg [7:0] phv_data_24; // @[executor.scala 448:22]
  reg [7:0] phv_data_25; // @[executor.scala 448:22]
  reg [7:0] phv_data_26; // @[executor.scala 448:22]
  reg [7:0] phv_data_27; // @[executor.scala 448:22]
  reg [7:0] phv_data_28; // @[executor.scala 448:22]
  reg [7:0] phv_data_29; // @[executor.scala 448:22]
  reg [7:0] phv_data_30; // @[executor.scala 448:22]
  reg [7:0] phv_data_31; // @[executor.scala 448:22]
  reg [7:0] phv_data_32; // @[executor.scala 448:22]
  reg [7:0] phv_data_33; // @[executor.scala 448:22]
  reg [7:0] phv_data_34; // @[executor.scala 448:22]
  reg [7:0] phv_data_35; // @[executor.scala 448:22]
  reg [7:0] phv_data_36; // @[executor.scala 448:22]
  reg [7:0] phv_data_37; // @[executor.scala 448:22]
  reg [7:0] phv_data_38; // @[executor.scala 448:22]
  reg [7:0] phv_data_39; // @[executor.scala 448:22]
  reg [7:0] phv_data_40; // @[executor.scala 448:22]
  reg [7:0] phv_data_41; // @[executor.scala 448:22]
  reg [7:0] phv_data_42; // @[executor.scala 448:22]
  reg [7:0] phv_data_43; // @[executor.scala 448:22]
  reg [7:0] phv_data_44; // @[executor.scala 448:22]
  reg [7:0] phv_data_45; // @[executor.scala 448:22]
  reg [7:0] phv_data_46; // @[executor.scala 448:22]
  reg [7:0] phv_data_47; // @[executor.scala 448:22]
  reg [7:0] phv_data_48; // @[executor.scala 448:22]
  reg [7:0] phv_data_49; // @[executor.scala 448:22]
  reg [7:0] phv_data_50; // @[executor.scala 448:22]
  reg [7:0] phv_data_51; // @[executor.scala 448:22]
  reg [7:0] phv_data_52; // @[executor.scala 448:22]
  reg [7:0] phv_data_53; // @[executor.scala 448:22]
  reg [7:0] phv_data_54; // @[executor.scala 448:22]
  reg [7:0] phv_data_55; // @[executor.scala 448:22]
  reg [7:0] phv_data_56; // @[executor.scala 448:22]
  reg [7:0] phv_data_57; // @[executor.scala 448:22]
  reg [7:0] phv_data_58; // @[executor.scala 448:22]
  reg [7:0] phv_data_59; // @[executor.scala 448:22]
  reg [7:0] phv_data_60; // @[executor.scala 448:22]
  reg [7:0] phv_data_61; // @[executor.scala 448:22]
  reg [7:0] phv_data_62; // @[executor.scala 448:22]
  reg [7:0] phv_data_63; // @[executor.scala 448:22]
  reg [7:0] phv_data_64; // @[executor.scala 448:22]
  reg [7:0] phv_data_65; // @[executor.scala 448:22]
  reg [7:0] phv_data_66; // @[executor.scala 448:22]
  reg [7:0] phv_data_67; // @[executor.scala 448:22]
  reg [7:0] phv_data_68; // @[executor.scala 448:22]
  reg [7:0] phv_data_69; // @[executor.scala 448:22]
  reg [7:0] phv_data_70; // @[executor.scala 448:22]
  reg [7:0] phv_data_71; // @[executor.scala 448:22]
  reg [7:0] phv_data_72; // @[executor.scala 448:22]
  reg [7:0] phv_data_73; // @[executor.scala 448:22]
  reg [7:0] phv_data_74; // @[executor.scala 448:22]
  reg [7:0] phv_data_75; // @[executor.scala 448:22]
  reg [7:0] phv_data_76; // @[executor.scala 448:22]
  reg [7:0] phv_data_77; // @[executor.scala 448:22]
  reg [7:0] phv_data_78; // @[executor.scala 448:22]
  reg [7:0] phv_data_79; // @[executor.scala 448:22]
  reg [7:0] phv_data_80; // @[executor.scala 448:22]
  reg [7:0] phv_data_81; // @[executor.scala 448:22]
  reg [7:0] phv_data_82; // @[executor.scala 448:22]
  reg [7:0] phv_data_83; // @[executor.scala 448:22]
  reg [7:0] phv_data_84; // @[executor.scala 448:22]
  reg [7:0] phv_data_85; // @[executor.scala 448:22]
  reg [7:0] phv_data_86; // @[executor.scala 448:22]
  reg [7:0] phv_data_87; // @[executor.scala 448:22]
  reg [7:0] phv_data_88; // @[executor.scala 448:22]
  reg [7:0] phv_data_89; // @[executor.scala 448:22]
  reg [7:0] phv_data_90; // @[executor.scala 448:22]
  reg [7:0] phv_data_91; // @[executor.scala 448:22]
  reg [7:0] phv_data_92; // @[executor.scala 448:22]
  reg [7:0] phv_data_93; // @[executor.scala 448:22]
  reg [7:0] phv_data_94; // @[executor.scala 448:22]
  reg [7:0] phv_data_95; // @[executor.scala 448:22]
  reg [7:0] phv_data_96; // @[executor.scala 448:22]
  reg [7:0] phv_data_97; // @[executor.scala 448:22]
  reg [7:0] phv_data_98; // @[executor.scala 448:22]
  reg [7:0] phv_data_99; // @[executor.scala 448:22]
  reg [7:0] phv_data_100; // @[executor.scala 448:22]
  reg [7:0] phv_data_101; // @[executor.scala 448:22]
  reg [7:0] phv_data_102; // @[executor.scala 448:22]
  reg [7:0] phv_data_103; // @[executor.scala 448:22]
  reg [7:0] phv_data_104; // @[executor.scala 448:22]
  reg [7:0] phv_data_105; // @[executor.scala 448:22]
  reg [7:0] phv_data_106; // @[executor.scala 448:22]
  reg [7:0] phv_data_107; // @[executor.scala 448:22]
  reg [7:0] phv_data_108; // @[executor.scala 448:22]
  reg [7:0] phv_data_109; // @[executor.scala 448:22]
  reg [7:0] phv_data_110; // @[executor.scala 448:22]
  reg [7:0] phv_data_111; // @[executor.scala 448:22]
  reg [7:0] phv_data_112; // @[executor.scala 448:22]
  reg [7:0] phv_data_113; // @[executor.scala 448:22]
  reg [7:0] phv_data_114; // @[executor.scala 448:22]
  reg [7:0] phv_data_115; // @[executor.scala 448:22]
  reg [7:0] phv_data_116; // @[executor.scala 448:22]
  reg [7:0] phv_data_117; // @[executor.scala 448:22]
  reg [7:0] phv_data_118; // @[executor.scala 448:22]
  reg [7:0] phv_data_119; // @[executor.scala 448:22]
  reg [7:0] phv_data_120; // @[executor.scala 448:22]
  reg [7:0] phv_data_121; // @[executor.scala 448:22]
  reg [7:0] phv_data_122; // @[executor.scala 448:22]
  reg [7:0] phv_data_123; // @[executor.scala 448:22]
  reg [7:0] phv_data_124; // @[executor.scala 448:22]
  reg [7:0] phv_data_125; // @[executor.scala 448:22]
  reg [7:0] phv_data_126; // @[executor.scala 448:22]
  reg [7:0] phv_data_127; // @[executor.scala 448:22]
  reg [7:0] phv_data_128; // @[executor.scala 448:22]
  reg [7:0] phv_data_129; // @[executor.scala 448:22]
  reg [7:0] phv_data_130; // @[executor.scala 448:22]
  reg [7:0] phv_data_131; // @[executor.scala 448:22]
  reg [7:0] phv_data_132; // @[executor.scala 448:22]
  reg [7:0] phv_data_133; // @[executor.scala 448:22]
  reg [7:0] phv_data_134; // @[executor.scala 448:22]
  reg [7:0] phv_data_135; // @[executor.scala 448:22]
  reg [7:0] phv_data_136; // @[executor.scala 448:22]
  reg [7:0] phv_data_137; // @[executor.scala 448:22]
  reg [7:0] phv_data_138; // @[executor.scala 448:22]
  reg [7:0] phv_data_139; // @[executor.scala 448:22]
  reg [7:0] phv_data_140; // @[executor.scala 448:22]
  reg [7:0] phv_data_141; // @[executor.scala 448:22]
  reg [7:0] phv_data_142; // @[executor.scala 448:22]
  reg [7:0] phv_data_143; // @[executor.scala 448:22]
  reg [7:0] phv_data_144; // @[executor.scala 448:22]
  reg [7:0] phv_data_145; // @[executor.scala 448:22]
  reg [7:0] phv_data_146; // @[executor.scala 448:22]
  reg [7:0] phv_data_147; // @[executor.scala 448:22]
  reg [7:0] phv_data_148; // @[executor.scala 448:22]
  reg [7:0] phv_data_149; // @[executor.scala 448:22]
  reg [7:0] phv_data_150; // @[executor.scala 448:22]
  reg [7:0] phv_data_151; // @[executor.scala 448:22]
  reg [7:0] phv_data_152; // @[executor.scala 448:22]
  reg [7:0] phv_data_153; // @[executor.scala 448:22]
  reg [7:0] phv_data_154; // @[executor.scala 448:22]
  reg [7:0] phv_data_155; // @[executor.scala 448:22]
  reg [7:0] phv_data_156; // @[executor.scala 448:22]
  reg [7:0] phv_data_157; // @[executor.scala 448:22]
  reg [7:0] phv_data_158; // @[executor.scala 448:22]
  reg [7:0] phv_data_159; // @[executor.scala 448:22]
  reg [7:0] phv_data_160; // @[executor.scala 448:22]
  reg [7:0] phv_data_161; // @[executor.scala 448:22]
  reg [7:0] phv_data_162; // @[executor.scala 448:22]
  reg [7:0] phv_data_163; // @[executor.scala 448:22]
  reg [7:0] phv_data_164; // @[executor.scala 448:22]
  reg [7:0] phv_data_165; // @[executor.scala 448:22]
  reg [7:0] phv_data_166; // @[executor.scala 448:22]
  reg [7:0] phv_data_167; // @[executor.scala 448:22]
  reg [7:0] phv_data_168; // @[executor.scala 448:22]
  reg [7:0] phv_data_169; // @[executor.scala 448:22]
  reg [7:0] phv_data_170; // @[executor.scala 448:22]
  reg [7:0] phv_data_171; // @[executor.scala 448:22]
  reg [7:0] phv_data_172; // @[executor.scala 448:22]
  reg [7:0] phv_data_173; // @[executor.scala 448:22]
  reg [7:0] phv_data_174; // @[executor.scala 448:22]
  reg [7:0] phv_data_175; // @[executor.scala 448:22]
  reg [7:0] phv_data_176; // @[executor.scala 448:22]
  reg [7:0] phv_data_177; // @[executor.scala 448:22]
  reg [7:0] phv_data_178; // @[executor.scala 448:22]
  reg [7:0] phv_data_179; // @[executor.scala 448:22]
  reg [7:0] phv_data_180; // @[executor.scala 448:22]
  reg [7:0] phv_data_181; // @[executor.scala 448:22]
  reg [7:0] phv_data_182; // @[executor.scala 448:22]
  reg [7:0] phv_data_183; // @[executor.scala 448:22]
  reg [7:0] phv_data_184; // @[executor.scala 448:22]
  reg [7:0] phv_data_185; // @[executor.scala 448:22]
  reg [7:0] phv_data_186; // @[executor.scala 448:22]
  reg [7:0] phv_data_187; // @[executor.scala 448:22]
  reg [7:0] phv_data_188; // @[executor.scala 448:22]
  reg [7:0] phv_data_189; // @[executor.scala 448:22]
  reg [7:0] phv_data_190; // @[executor.scala 448:22]
  reg [7:0] phv_data_191; // @[executor.scala 448:22]
  reg [7:0] phv_data_192; // @[executor.scala 448:22]
  reg [7:0] phv_data_193; // @[executor.scala 448:22]
  reg [7:0] phv_data_194; // @[executor.scala 448:22]
  reg [7:0] phv_data_195; // @[executor.scala 448:22]
  reg [7:0] phv_data_196; // @[executor.scala 448:22]
  reg [7:0] phv_data_197; // @[executor.scala 448:22]
  reg [7:0] phv_data_198; // @[executor.scala 448:22]
  reg [7:0] phv_data_199; // @[executor.scala 448:22]
  reg [7:0] phv_data_200; // @[executor.scala 448:22]
  reg [7:0] phv_data_201; // @[executor.scala 448:22]
  reg [7:0] phv_data_202; // @[executor.scala 448:22]
  reg [7:0] phv_data_203; // @[executor.scala 448:22]
  reg [7:0] phv_data_204; // @[executor.scala 448:22]
  reg [7:0] phv_data_205; // @[executor.scala 448:22]
  reg [7:0] phv_data_206; // @[executor.scala 448:22]
  reg [7:0] phv_data_207; // @[executor.scala 448:22]
  reg [7:0] phv_data_208; // @[executor.scala 448:22]
  reg [7:0] phv_data_209; // @[executor.scala 448:22]
  reg [7:0] phv_data_210; // @[executor.scala 448:22]
  reg [7:0] phv_data_211; // @[executor.scala 448:22]
  reg [7:0] phv_data_212; // @[executor.scala 448:22]
  reg [7:0] phv_data_213; // @[executor.scala 448:22]
  reg [7:0] phv_data_214; // @[executor.scala 448:22]
  reg [7:0] phv_data_215; // @[executor.scala 448:22]
  reg [7:0] phv_data_216; // @[executor.scala 448:22]
  reg [7:0] phv_data_217; // @[executor.scala 448:22]
  reg [7:0] phv_data_218; // @[executor.scala 448:22]
  reg [7:0] phv_data_219; // @[executor.scala 448:22]
  reg [7:0] phv_data_220; // @[executor.scala 448:22]
  reg [7:0] phv_data_221; // @[executor.scala 448:22]
  reg [7:0] phv_data_222; // @[executor.scala 448:22]
  reg [7:0] phv_data_223; // @[executor.scala 448:22]
  reg [7:0] phv_data_224; // @[executor.scala 448:22]
  reg [7:0] phv_data_225; // @[executor.scala 448:22]
  reg [7:0] phv_data_226; // @[executor.scala 448:22]
  reg [7:0] phv_data_227; // @[executor.scala 448:22]
  reg [7:0] phv_data_228; // @[executor.scala 448:22]
  reg [7:0] phv_data_229; // @[executor.scala 448:22]
  reg [7:0] phv_data_230; // @[executor.scala 448:22]
  reg [7:0] phv_data_231; // @[executor.scala 448:22]
  reg [7:0] phv_data_232; // @[executor.scala 448:22]
  reg [7:0] phv_data_233; // @[executor.scala 448:22]
  reg [7:0] phv_data_234; // @[executor.scala 448:22]
  reg [7:0] phv_data_235; // @[executor.scala 448:22]
  reg [7:0] phv_data_236; // @[executor.scala 448:22]
  reg [7:0] phv_data_237; // @[executor.scala 448:22]
  reg [7:0] phv_data_238; // @[executor.scala 448:22]
  reg [7:0] phv_data_239; // @[executor.scala 448:22]
  reg [7:0] phv_data_240; // @[executor.scala 448:22]
  reg [7:0] phv_data_241; // @[executor.scala 448:22]
  reg [7:0] phv_data_242; // @[executor.scala 448:22]
  reg [7:0] phv_data_243; // @[executor.scala 448:22]
  reg [7:0] phv_data_244; // @[executor.scala 448:22]
  reg [7:0] phv_data_245; // @[executor.scala 448:22]
  reg [7:0] phv_data_246; // @[executor.scala 448:22]
  reg [7:0] phv_data_247; // @[executor.scala 448:22]
  reg [7:0] phv_data_248; // @[executor.scala 448:22]
  reg [7:0] phv_data_249; // @[executor.scala 448:22]
  reg [7:0] phv_data_250; // @[executor.scala 448:22]
  reg [7:0] phv_data_251; // @[executor.scala 448:22]
  reg [7:0] phv_data_252; // @[executor.scala 448:22]
  reg [7:0] phv_data_253; // @[executor.scala 448:22]
  reg [7:0] phv_data_254; // @[executor.scala 448:22]
  reg [7:0] phv_data_255; // @[executor.scala 448:22]
  reg [15:0] phv_header_0; // @[executor.scala 448:22]
  reg [15:0] phv_header_1; // @[executor.scala 448:22]
  reg [15:0] phv_header_2; // @[executor.scala 448:22]
  reg [15:0] phv_header_3; // @[executor.scala 448:22]
  reg [15:0] phv_header_4; // @[executor.scala 448:22]
  reg [15:0] phv_header_5; // @[executor.scala 448:22]
  reg [15:0] phv_header_6; // @[executor.scala 448:22]
  reg [15:0] phv_header_7; // @[executor.scala 448:22]
  reg [15:0] phv_header_8; // @[executor.scala 448:22]
  reg [15:0] phv_header_9; // @[executor.scala 448:22]
  reg [15:0] phv_header_10; // @[executor.scala 448:22]
  reg [15:0] phv_header_11; // @[executor.scala 448:22]
  reg [15:0] phv_header_12; // @[executor.scala 448:22]
  reg [15:0] phv_header_13; // @[executor.scala 448:22]
  reg [15:0] phv_header_14; // @[executor.scala 448:22]
  reg [15:0] phv_header_15; // @[executor.scala 448:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 448:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 448:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 448:22]
  reg [3:0] phv_next_processor_id; // @[executor.scala 448:22]
  reg  phv_next_config_id; // @[executor.scala 448:22]
  reg  phv_is_valid_processor; // @[executor.scala 448:22]
  reg [31:0] vliw_0; // @[executor.scala 452:23]
  reg [31:0] vliw_1; // @[executor.scala 452:23]
  reg [31:0] vliw_2; // @[executor.scala 452:23]
  reg [31:0] vliw_3; // @[executor.scala 452:23]
  reg [31:0] vliw_4; // @[executor.scala 452:23]
  reg [31:0] vliw_5; // @[executor.scala 452:23]
  reg [31:0] vliw_6; // @[executor.scala 452:23]
  reg [31:0] vliw_7; // @[executor.scala 452:23]
  reg [31:0] field_0; // @[executor.scala 454:24]
  reg [31:0] field_1; // @[executor.scala 454:24]
  reg [31:0] field_2; // @[executor.scala 454:24]
  reg [31:0] field_3; // @[executor.scala 454:24]
  reg [31:0] field_4; // @[executor.scala 454:24]
  reg [31:0] field_5; // @[executor.scala 454:24]
  reg [31:0] field_6; // @[executor.scala 454:24]
  reg [31:0] field_7; // @[executor.scala 454:24]
  reg [3:0] mask_0; // @[executor.scala 456:23]
  reg [3:0] mask_1; // @[executor.scala 456:23]
  reg [3:0] mask_2; // @[executor.scala 456:23]
  reg [3:0] mask_3; // @[executor.scala 456:23]
  reg [3:0] mask_4; // @[executor.scala 456:23]
  reg [3:0] mask_5; // @[executor.scala 456:23]
  reg [3:0] mask_6; // @[executor.scala 456:23]
  reg [3:0] mask_7; // @[executor.scala 456:23]
  reg [5:0] dst_offset_0; // @[executor.scala 458:29]
  reg [5:0] dst_offset_1; // @[executor.scala 458:29]
  reg [5:0] dst_offset_2; // @[executor.scala 458:29]
  reg [5:0] dst_offset_3; // @[executor.scala 458:29]
  reg [5:0] dst_offset_4; // @[executor.scala 458:29]
  reg [5:0] dst_offset_5; // @[executor.scala 458:29]
  reg [5:0] dst_offset_6; // @[executor.scala 458:29]
  reg [5:0] dst_offset_7; // @[executor.scala 458:29]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2 = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8466 = {{2'd0}, dst_offset_0}; // @[executor.scala 473:49]
  wire [7:0] byte_ = field_0[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_0 = mask_0[0] ? byte_ : phv_data_3; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_1 = field_0[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1 = mask_0[1] ? byte_1 : phv_data_2; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_2 = field_0[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2 = mask_0[2] ? byte_2 : phv_data_1; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_3 = field_0[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3 = mask_0[3] ? byte_3 : phv_data_0; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_4 = _GEN_8466 == 8'h0 ? _GEN_0 : phv_data_3; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_5 = _GEN_8466 == 8'h0 ? _GEN_1 : phv_data_2; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_6 = _GEN_8466 == 8'h0 ? _GEN_2 : phv_data_1; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_7 = _GEN_8466 == 8'h0 ? _GEN_3 : phv_data_0; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_8 = mask_0[0] ? byte_ : phv_data_7; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_9 = mask_0[1] ? byte_1 : phv_data_6; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_10 = mask_0[2] ? byte_2 : phv_data_5; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_11 = mask_0[3] ? byte_3 : phv_data_4; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_12 = _GEN_8466 == 8'h1 ? _GEN_8 : phv_data_7; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_13 = _GEN_8466 == 8'h1 ? _GEN_9 : phv_data_6; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_14 = _GEN_8466 == 8'h1 ? _GEN_10 : phv_data_5; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_15 = _GEN_8466 == 8'h1 ? _GEN_11 : phv_data_4; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_16 = mask_0[0] ? byte_ : phv_data_11; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_17 = mask_0[1] ? byte_1 : phv_data_10; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_18 = mask_0[2] ? byte_2 : phv_data_9; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_19 = mask_0[3] ? byte_3 : phv_data_8; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_20 = _GEN_8466 == 8'h2 ? _GEN_16 : phv_data_11; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_21 = _GEN_8466 == 8'h2 ? _GEN_17 : phv_data_10; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_22 = _GEN_8466 == 8'h2 ? _GEN_18 : phv_data_9; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_23 = _GEN_8466 == 8'h2 ? _GEN_19 : phv_data_8; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_24 = mask_0[0] ? byte_ : phv_data_15; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_25 = mask_0[1] ? byte_1 : phv_data_14; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_26 = mask_0[2] ? byte_2 : phv_data_13; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_27 = mask_0[3] ? byte_3 : phv_data_12; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_28 = _GEN_8466 == 8'h3 ? _GEN_24 : phv_data_15; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_29 = _GEN_8466 == 8'h3 ? _GEN_25 : phv_data_14; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_30 = _GEN_8466 == 8'h3 ? _GEN_26 : phv_data_13; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_31 = _GEN_8466 == 8'h3 ? _GEN_27 : phv_data_12; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_32 = mask_0[0] ? byte_ : phv_data_19; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_33 = mask_0[1] ? byte_1 : phv_data_18; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_34 = mask_0[2] ? byte_2 : phv_data_17; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_35 = mask_0[3] ? byte_3 : phv_data_16; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_36 = _GEN_8466 == 8'h4 ? _GEN_32 : phv_data_19; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_37 = _GEN_8466 == 8'h4 ? _GEN_33 : phv_data_18; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_38 = _GEN_8466 == 8'h4 ? _GEN_34 : phv_data_17; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_39 = _GEN_8466 == 8'h4 ? _GEN_35 : phv_data_16; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_40 = mask_0[0] ? byte_ : phv_data_23; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_41 = mask_0[1] ? byte_1 : phv_data_22; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_42 = mask_0[2] ? byte_2 : phv_data_21; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_43 = mask_0[3] ? byte_3 : phv_data_20; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_44 = _GEN_8466 == 8'h5 ? _GEN_40 : phv_data_23; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_45 = _GEN_8466 == 8'h5 ? _GEN_41 : phv_data_22; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_46 = _GEN_8466 == 8'h5 ? _GEN_42 : phv_data_21; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_47 = _GEN_8466 == 8'h5 ? _GEN_43 : phv_data_20; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_48 = mask_0[0] ? byte_ : phv_data_27; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_49 = mask_0[1] ? byte_1 : phv_data_26; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_50 = mask_0[2] ? byte_2 : phv_data_25; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_51 = mask_0[3] ? byte_3 : phv_data_24; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_52 = _GEN_8466 == 8'h6 ? _GEN_48 : phv_data_27; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_53 = _GEN_8466 == 8'h6 ? _GEN_49 : phv_data_26; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_54 = _GEN_8466 == 8'h6 ? _GEN_50 : phv_data_25; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_55 = _GEN_8466 == 8'h6 ? _GEN_51 : phv_data_24; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_56 = mask_0[0] ? byte_ : phv_data_31; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_57 = mask_0[1] ? byte_1 : phv_data_30; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_58 = mask_0[2] ? byte_2 : phv_data_29; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_59 = mask_0[3] ? byte_3 : phv_data_28; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_60 = _GEN_8466 == 8'h7 ? _GEN_56 : phv_data_31; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_61 = _GEN_8466 == 8'h7 ? _GEN_57 : phv_data_30; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_62 = _GEN_8466 == 8'h7 ? _GEN_58 : phv_data_29; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_63 = _GEN_8466 == 8'h7 ? _GEN_59 : phv_data_28; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_64 = mask_0[0] ? byte_ : phv_data_35; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_65 = mask_0[1] ? byte_1 : phv_data_34; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_66 = mask_0[2] ? byte_2 : phv_data_33; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_67 = mask_0[3] ? byte_3 : phv_data_32; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_68 = _GEN_8466 == 8'h8 ? _GEN_64 : phv_data_35; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_69 = _GEN_8466 == 8'h8 ? _GEN_65 : phv_data_34; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_70 = _GEN_8466 == 8'h8 ? _GEN_66 : phv_data_33; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_71 = _GEN_8466 == 8'h8 ? _GEN_67 : phv_data_32; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_72 = mask_0[0] ? byte_ : phv_data_39; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_73 = mask_0[1] ? byte_1 : phv_data_38; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_74 = mask_0[2] ? byte_2 : phv_data_37; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_75 = mask_0[3] ? byte_3 : phv_data_36; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_76 = _GEN_8466 == 8'h9 ? _GEN_72 : phv_data_39; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_77 = _GEN_8466 == 8'h9 ? _GEN_73 : phv_data_38; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_78 = _GEN_8466 == 8'h9 ? _GEN_74 : phv_data_37; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_79 = _GEN_8466 == 8'h9 ? _GEN_75 : phv_data_36; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_80 = mask_0[0] ? byte_ : phv_data_43; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_81 = mask_0[1] ? byte_1 : phv_data_42; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_82 = mask_0[2] ? byte_2 : phv_data_41; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_83 = mask_0[3] ? byte_3 : phv_data_40; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_84 = _GEN_8466 == 8'ha ? _GEN_80 : phv_data_43; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_85 = _GEN_8466 == 8'ha ? _GEN_81 : phv_data_42; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_86 = _GEN_8466 == 8'ha ? _GEN_82 : phv_data_41; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_87 = _GEN_8466 == 8'ha ? _GEN_83 : phv_data_40; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_88 = mask_0[0] ? byte_ : phv_data_47; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_89 = mask_0[1] ? byte_1 : phv_data_46; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_90 = mask_0[2] ? byte_2 : phv_data_45; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_91 = mask_0[3] ? byte_3 : phv_data_44; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_92 = _GEN_8466 == 8'hb ? _GEN_88 : phv_data_47; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_93 = _GEN_8466 == 8'hb ? _GEN_89 : phv_data_46; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_94 = _GEN_8466 == 8'hb ? _GEN_90 : phv_data_45; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_95 = _GEN_8466 == 8'hb ? _GEN_91 : phv_data_44; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_96 = mask_0[0] ? byte_ : phv_data_51; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_97 = mask_0[1] ? byte_1 : phv_data_50; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_98 = mask_0[2] ? byte_2 : phv_data_49; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_99 = mask_0[3] ? byte_3 : phv_data_48; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_100 = _GEN_8466 == 8'hc ? _GEN_96 : phv_data_51; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_101 = _GEN_8466 == 8'hc ? _GEN_97 : phv_data_50; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_102 = _GEN_8466 == 8'hc ? _GEN_98 : phv_data_49; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_103 = _GEN_8466 == 8'hc ? _GEN_99 : phv_data_48; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_104 = mask_0[0] ? byte_ : phv_data_55; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_105 = mask_0[1] ? byte_1 : phv_data_54; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_106 = mask_0[2] ? byte_2 : phv_data_53; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_107 = mask_0[3] ? byte_3 : phv_data_52; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_108 = _GEN_8466 == 8'hd ? _GEN_104 : phv_data_55; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_109 = _GEN_8466 == 8'hd ? _GEN_105 : phv_data_54; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_110 = _GEN_8466 == 8'hd ? _GEN_106 : phv_data_53; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_111 = _GEN_8466 == 8'hd ? _GEN_107 : phv_data_52; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_112 = mask_0[0] ? byte_ : phv_data_59; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_113 = mask_0[1] ? byte_1 : phv_data_58; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_114 = mask_0[2] ? byte_2 : phv_data_57; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_115 = mask_0[3] ? byte_3 : phv_data_56; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_116 = _GEN_8466 == 8'he ? _GEN_112 : phv_data_59; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_117 = _GEN_8466 == 8'he ? _GEN_113 : phv_data_58; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_118 = _GEN_8466 == 8'he ? _GEN_114 : phv_data_57; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_119 = _GEN_8466 == 8'he ? _GEN_115 : phv_data_56; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_120 = mask_0[0] ? byte_ : phv_data_63; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_121 = mask_0[1] ? byte_1 : phv_data_62; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_122 = mask_0[2] ? byte_2 : phv_data_61; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_123 = mask_0[3] ? byte_3 : phv_data_60; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_124 = _GEN_8466 == 8'hf ? _GEN_120 : phv_data_63; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_125 = _GEN_8466 == 8'hf ? _GEN_121 : phv_data_62; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_126 = _GEN_8466 == 8'hf ? _GEN_122 : phv_data_61; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_127 = _GEN_8466 == 8'hf ? _GEN_123 : phv_data_60; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_128 = mask_0[0] ? byte_ : phv_data_67; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_129 = mask_0[1] ? byte_1 : phv_data_66; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_130 = mask_0[2] ? byte_2 : phv_data_65; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_131 = mask_0[3] ? byte_3 : phv_data_64; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_132 = _GEN_8466 == 8'h10 ? _GEN_128 : phv_data_67; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_133 = _GEN_8466 == 8'h10 ? _GEN_129 : phv_data_66; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_134 = _GEN_8466 == 8'h10 ? _GEN_130 : phv_data_65; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_135 = _GEN_8466 == 8'h10 ? _GEN_131 : phv_data_64; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_136 = mask_0[0] ? byte_ : phv_data_71; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_137 = mask_0[1] ? byte_1 : phv_data_70; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_138 = mask_0[2] ? byte_2 : phv_data_69; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_139 = mask_0[3] ? byte_3 : phv_data_68; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_140 = _GEN_8466 == 8'h11 ? _GEN_136 : phv_data_71; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_141 = _GEN_8466 == 8'h11 ? _GEN_137 : phv_data_70; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_142 = _GEN_8466 == 8'h11 ? _GEN_138 : phv_data_69; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_143 = _GEN_8466 == 8'h11 ? _GEN_139 : phv_data_68; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_144 = mask_0[0] ? byte_ : phv_data_75; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_145 = mask_0[1] ? byte_1 : phv_data_74; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_146 = mask_0[2] ? byte_2 : phv_data_73; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_147 = mask_0[3] ? byte_3 : phv_data_72; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_148 = _GEN_8466 == 8'h12 ? _GEN_144 : phv_data_75; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_149 = _GEN_8466 == 8'h12 ? _GEN_145 : phv_data_74; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_150 = _GEN_8466 == 8'h12 ? _GEN_146 : phv_data_73; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_151 = _GEN_8466 == 8'h12 ? _GEN_147 : phv_data_72; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_152 = mask_0[0] ? byte_ : phv_data_79; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_153 = mask_0[1] ? byte_1 : phv_data_78; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_154 = mask_0[2] ? byte_2 : phv_data_77; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_155 = mask_0[3] ? byte_3 : phv_data_76; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_156 = _GEN_8466 == 8'h13 ? _GEN_152 : phv_data_79; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_157 = _GEN_8466 == 8'h13 ? _GEN_153 : phv_data_78; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_158 = _GEN_8466 == 8'h13 ? _GEN_154 : phv_data_77; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_159 = _GEN_8466 == 8'h13 ? _GEN_155 : phv_data_76; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_160 = mask_0[0] ? byte_ : phv_data_83; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_161 = mask_0[1] ? byte_1 : phv_data_82; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_162 = mask_0[2] ? byte_2 : phv_data_81; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_163 = mask_0[3] ? byte_3 : phv_data_80; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_164 = _GEN_8466 == 8'h14 ? _GEN_160 : phv_data_83; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_165 = _GEN_8466 == 8'h14 ? _GEN_161 : phv_data_82; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_166 = _GEN_8466 == 8'h14 ? _GEN_162 : phv_data_81; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_167 = _GEN_8466 == 8'h14 ? _GEN_163 : phv_data_80; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_168 = mask_0[0] ? byte_ : phv_data_87; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_169 = mask_0[1] ? byte_1 : phv_data_86; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_170 = mask_0[2] ? byte_2 : phv_data_85; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_171 = mask_0[3] ? byte_3 : phv_data_84; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_172 = _GEN_8466 == 8'h15 ? _GEN_168 : phv_data_87; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_173 = _GEN_8466 == 8'h15 ? _GEN_169 : phv_data_86; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_174 = _GEN_8466 == 8'h15 ? _GEN_170 : phv_data_85; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_175 = _GEN_8466 == 8'h15 ? _GEN_171 : phv_data_84; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_176 = mask_0[0] ? byte_ : phv_data_91; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_177 = mask_0[1] ? byte_1 : phv_data_90; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_178 = mask_0[2] ? byte_2 : phv_data_89; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_179 = mask_0[3] ? byte_3 : phv_data_88; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_180 = _GEN_8466 == 8'h16 ? _GEN_176 : phv_data_91; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_181 = _GEN_8466 == 8'h16 ? _GEN_177 : phv_data_90; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_182 = _GEN_8466 == 8'h16 ? _GEN_178 : phv_data_89; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_183 = _GEN_8466 == 8'h16 ? _GEN_179 : phv_data_88; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_184 = mask_0[0] ? byte_ : phv_data_95; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_185 = mask_0[1] ? byte_1 : phv_data_94; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_186 = mask_0[2] ? byte_2 : phv_data_93; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_187 = mask_0[3] ? byte_3 : phv_data_92; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_188 = _GEN_8466 == 8'h17 ? _GEN_184 : phv_data_95; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_189 = _GEN_8466 == 8'h17 ? _GEN_185 : phv_data_94; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_190 = _GEN_8466 == 8'h17 ? _GEN_186 : phv_data_93; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_191 = _GEN_8466 == 8'h17 ? _GEN_187 : phv_data_92; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_192 = mask_0[0] ? byte_ : phv_data_99; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_193 = mask_0[1] ? byte_1 : phv_data_98; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_194 = mask_0[2] ? byte_2 : phv_data_97; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_195 = mask_0[3] ? byte_3 : phv_data_96; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_196 = _GEN_8466 == 8'h18 ? _GEN_192 : phv_data_99; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_197 = _GEN_8466 == 8'h18 ? _GEN_193 : phv_data_98; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_198 = _GEN_8466 == 8'h18 ? _GEN_194 : phv_data_97; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_199 = _GEN_8466 == 8'h18 ? _GEN_195 : phv_data_96; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_200 = mask_0[0] ? byte_ : phv_data_103; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_201 = mask_0[1] ? byte_1 : phv_data_102; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_202 = mask_0[2] ? byte_2 : phv_data_101; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_203 = mask_0[3] ? byte_3 : phv_data_100; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_204 = _GEN_8466 == 8'h19 ? _GEN_200 : phv_data_103; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_205 = _GEN_8466 == 8'h19 ? _GEN_201 : phv_data_102; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_206 = _GEN_8466 == 8'h19 ? _GEN_202 : phv_data_101; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_207 = _GEN_8466 == 8'h19 ? _GEN_203 : phv_data_100; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_208 = mask_0[0] ? byte_ : phv_data_107; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_209 = mask_0[1] ? byte_1 : phv_data_106; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_210 = mask_0[2] ? byte_2 : phv_data_105; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_211 = mask_0[3] ? byte_3 : phv_data_104; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_212 = _GEN_8466 == 8'h1a ? _GEN_208 : phv_data_107; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_213 = _GEN_8466 == 8'h1a ? _GEN_209 : phv_data_106; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_214 = _GEN_8466 == 8'h1a ? _GEN_210 : phv_data_105; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_215 = _GEN_8466 == 8'h1a ? _GEN_211 : phv_data_104; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_216 = mask_0[0] ? byte_ : phv_data_111; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_217 = mask_0[1] ? byte_1 : phv_data_110; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_218 = mask_0[2] ? byte_2 : phv_data_109; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_219 = mask_0[3] ? byte_3 : phv_data_108; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_220 = _GEN_8466 == 8'h1b ? _GEN_216 : phv_data_111; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_221 = _GEN_8466 == 8'h1b ? _GEN_217 : phv_data_110; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_222 = _GEN_8466 == 8'h1b ? _GEN_218 : phv_data_109; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_223 = _GEN_8466 == 8'h1b ? _GEN_219 : phv_data_108; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_224 = mask_0[0] ? byte_ : phv_data_115; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_225 = mask_0[1] ? byte_1 : phv_data_114; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_226 = mask_0[2] ? byte_2 : phv_data_113; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_227 = mask_0[3] ? byte_3 : phv_data_112; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_228 = _GEN_8466 == 8'h1c ? _GEN_224 : phv_data_115; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_229 = _GEN_8466 == 8'h1c ? _GEN_225 : phv_data_114; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_230 = _GEN_8466 == 8'h1c ? _GEN_226 : phv_data_113; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_231 = _GEN_8466 == 8'h1c ? _GEN_227 : phv_data_112; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_232 = mask_0[0] ? byte_ : phv_data_119; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_233 = mask_0[1] ? byte_1 : phv_data_118; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_234 = mask_0[2] ? byte_2 : phv_data_117; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_235 = mask_0[3] ? byte_3 : phv_data_116; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_236 = _GEN_8466 == 8'h1d ? _GEN_232 : phv_data_119; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_237 = _GEN_8466 == 8'h1d ? _GEN_233 : phv_data_118; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_238 = _GEN_8466 == 8'h1d ? _GEN_234 : phv_data_117; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_239 = _GEN_8466 == 8'h1d ? _GEN_235 : phv_data_116; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_240 = mask_0[0] ? byte_ : phv_data_123; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_241 = mask_0[1] ? byte_1 : phv_data_122; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_242 = mask_0[2] ? byte_2 : phv_data_121; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_243 = mask_0[3] ? byte_3 : phv_data_120; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_244 = _GEN_8466 == 8'h1e ? _GEN_240 : phv_data_123; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_245 = _GEN_8466 == 8'h1e ? _GEN_241 : phv_data_122; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_246 = _GEN_8466 == 8'h1e ? _GEN_242 : phv_data_121; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_247 = _GEN_8466 == 8'h1e ? _GEN_243 : phv_data_120; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_248 = mask_0[0] ? byte_ : phv_data_127; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_249 = mask_0[1] ? byte_1 : phv_data_126; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_250 = mask_0[2] ? byte_2 : phv_data_125; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_251 = mask_0[3] ? byte_3 : phv_data_124; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_252 = _GEN_8466 == 8'h1f ? _GEN_248 : phv_data_127; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_253 = _GEN_8466 == 8'h1f ? _GEN_249 : phv_data_126; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_254 = _GEN_8466 == 8'h1f ? _GEN_250 : phv_data_125; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_255 = _GEN_8466 == 8'h1f ? _GEN_251 : phv_data_124; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_256 = mask_0[0] ? byte_ : phv_data_131; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_257 = mask_0[1] ? byte_1 : phv_data_130; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_258 = mask_0[2] ? byte_2 : phv_data_129; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_259 = mask_0[3] ? byte_3 : phv_data_128; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_260 = _GEN_8466 == 8'h20 ? _GEN_256 : phv_data_131; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_261 = _GEN_8466 == 8'h20 ? _GEN_257 : phv_data_130; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_262 = _GEN_8466 == 8'h20 ? _GEN_258 : phv_data_129; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_263 = _GEN_8466 == 8'h20 ? _GEN_259 : phv_data_128; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_264 = mask_0[0] ? byte_ : phv_data_135; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_265 = mask_0[1] ? byte_1 : phv_data_134; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_266 = mask_0[2] ? byte_2 : phv_data_133; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_267 = mask_0[3] ? byte_3 : phv_data_132; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_268 = _GEN_8466 == 8'h21 ? _GEN_264 : phv_data_135; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_269 = _GEN_8466 == 8'h21 ? _GEN_265 : phv_data_134; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_270 = _GEN_8466 == 8'h21 ? _GEN_266 : phv_data_133; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_271 = _GEN_8466 == 8'h21 ? _GEN_267 : phv_data_132; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_272 = mask_0[0] ? byte_ : phv_data_139; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_273 = mask_0[1] ? byte_1 : phv_data_138; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_274 = mask_0[2] ? byte_2 : phv_data_137; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_275 = mask_0[3] ? byte_3 : phv_data_136; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_276 = _GEN_8466 == 8'h22 ? _GEN_272 : phv_data_139; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_277 = _GEN_8466 == 8'h22 ? _GEN_273 : phv_data_138; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_278 = _GEN_8466 == 8'h22 ? _GEN_274 : phv_data_137; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_279 = _GEN_8466 == 8'h22 ? _GEN_275 : phv_data_136; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_280 = mask_0[0] ? byte_ : phv_data_143; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_281 = mask_0[1] ? byte_1 : phv_data_142; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_282 = mask_0[2] ? byte_2 : phv_data_141; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_283 = mask_0[3] ? byte_3 : phv_data_140; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_284 = _GEN_8466 == 8'h23 ? _GEN_280 : phv_data_143; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_285 = _GEN_8466 == 8'h23 ? _GEN_281 : phv_data_142; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_286 = _GEN_8466 == 8'h23 ? _GEN_282 : phv_data_141; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_287 = _GEN_8466 == 8'h23 ? _GEN_283 : phv_data_140; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_288 = mask_0[0] ? byte_ : phv_data_147; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_289 = mask_0[1] ? byte_1 : phv_data_146; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_290 = mask_0[2] ? byte_2 : phv_data_145; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_291 = mask_0[3] ? byte_3 : phv_data_144; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_292 = _GEN_8466 == 8'h24 ? _GEN_288 : phv_data_147; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_293 = _GEN_8466 == 8'h24 ? _GEN_289 : phv_data_146; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_294 = _GEN_8466 == 8'h24 ? _GEN_290 : phv_data_145; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_295 = _GEN_8466 == 8'h24 ? _GEN_291 : phv_data_144; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_296 = mask_0[0] ? byte_ : phv_data_151; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_297 = mask_0[1] ? byte_1 : phv_data_150; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_298 = mask_0[2] ? byte_2 : phv_data_149; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_299 = mask_0[3] ? byte_3 : phv_data_148; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_300 = _GEN_8466 == 8'h25 ? _GEN_296 : phv_data_151; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_301 = _GEN_8466 == 8'h25 ? _GEN_297 : phv_data_150; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_302 = _GEN_8466 == 8'h25 ? _GEN_298 : phv_data_149; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_303 = _GEN_8466 == 8'h25 ? _GEN_299 : phv_data_148; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_304 = mask_0[0] ? byte_ : phv_data_155; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_305 = mask_0[1] ? byte_1 : phv_data_154; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_306 = mask_0[2] ? byte_2 : phv_data_153; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_307 = mask_0[3] ? byte_3 : phv_data_152; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_308 = _GEN_8466 == 8'h26 ? _GEN_304 : phv_data_155; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_309 = _GEN_8466 == 8'h26 ? _GEN_305 : phv_data_154; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_310 = _GEN_8466 == 8'h26 ? _GEN_306 : phv_data_153; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_311 = _GEN_8466 == 8'h26 ? _GEN_307 : phv_data_152; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_312 = mask_0[0] ? byte_ : phv_data_159; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_313 = mask_0[1] ? byte_1 : phv_data_158; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_314 = mask_0[2] ? byte_2 : phv_data_157; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_315 = mask_0[3] ? byte_3 : phv_data_156; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_316 = _GEN_8466 == 8'h27 ? _GEN_312 : phv_data_159; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_317 = _GEN_8466 == 8'h27 ? _GEN_313 : phv_data_158; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_318 = _GEN_8466 == 8'h27 ? _GEN_314 : phv_data_157; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_319 = _GEN_8466 == 8'h27 ? _GEN_315 : phv_data_156; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_320 = mask_0[0] ? byte_ : phv_data_163; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_321 = mask_0[1] ? byte_1 : phv_data_162; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_322 = mask_0[2] ? byte_2 : phv_data_161; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_323 = mask_0[3] ? byte_3 : phv_data_160; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_324 = _GEN_8466 == 8'h28 ? _GEN_320 : phv_data_163; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_325 = _GEN_8466 == 8'h28 ? _GEN_321 : phv_data_162; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_326 = _GEN_8466 == 8'h28 ? _GEN_322 : phv_data_161; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_327 = _GEN_8466 == 8'h28 ? _GEN_323 : phv_data_160; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_328 = mask_0[0] ? byte_ : phv_data_167; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_329 = mask_0[1] ? byte_1 : phv_data_166; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_330 = mask_0[2] ? byte_2 : phv_data_165; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_331 = mask_0[3] ? byte_3 : phv_data_164; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_332 = _GEN_8466 == 8'h29 ? _GEN_328 : phv_data_167; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_333 = _GEN_8466 == 8'h29 ? _GEN_329 : phv_data_166; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_334 = _GEN_8466 == 8'h29 ? _GEN_330 : phv_data_165; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_335 = _GEN_8466 == 8'h29 ? _GEN_331 : phv_data_164; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_336 = mask_0[0] ? byte_ : phv_data_171; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_337 = mask_0[1] ? byte_1 : phv_data_170; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_338 = mask_0[2] ? byte_2 : phv_data_169; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_339 = mask_0[3] ? byte_3 : phv_data_168; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_340 = _GEN_8466 == 8'h2a ? _GEN_336 : phv_data_171; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_341 = _GEN_8466 == 8'h2a ? _GEN_337 : phv_data_170; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_342 = _GEN_8466 == 8'h2a ? _GEN_338 : phv_data_169; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_343 = _GEN_8466 == 8'h2a ? _GEN_339 : phv_data_168; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_344 = mask_0[0] ? byte_ : phv_data_175; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_345 = mask_0[1] ? byte_1 : phv_data_174; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_346 = mask_0[2] ? byte_2 : phv_data_173; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_347 = mask_0[3] ? byte_3 : phv_data_172; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_348 = _GEN_8466 == 8'h2b ? _GEN_344 : phv_data_175; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_349 = _GEN_8466 == 8'h2b ? _GEN_345 : phv_data_174; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_350 = _GEN_8466 == 8'h2b ? _GEN_346 : phv_data_173; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_351 = _GEN_8466 == 8'h2b ? _GEN_347 : phv_data_172; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_352 = mask_0[0] ? byte_ : phv_data_179; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_353 = mask_0[1] ? byte_1 : phv_data_178; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_354 = mask_0[2] ? byte_2 : phv_data_177; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_355 = mask_0[3] ? byte_3 : phv_data_176; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_356 = _GEN_8466 == 8'h2c ? _GEN_352 : phv_data_179; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_357 = _GEN_8466 == 8'h2c ? _GEN_353 : phv_data_178; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_358 = _GEN_8466 == 8'h2c ? _GEN_354 : phv_data_177; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_359 = _GEN_8466 == 8'h2c ? _GEN_355 : phv_data_176; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_360 = mask_0[0] ? byte_ : phv_data_183; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_361 = mask_0[1] ? byte_1 : phv_data_182; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_362 = mask_0[2] ? byte_2 : phv_data_181; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_363 = mask_0[3] ? byte_3 : phv_data_180; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_364 = _GEN_8466 == 8'h2d ? _GEN_360 : phv_data_183; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_365 = _GEN_8466 == 8'h2d ? _GEN_361 : phv_data_182; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_366 = _GEN_8466 == 8'h2d ? _GEN_362 : phv_data_181; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_367 = _GEN_8466 == 8'h2d ? _GEN_363 : phv_data_180; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_368 = mask_0[0] ? byte_ : phv_data_187; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_369 = mask_0[1] ? byte_1 : phv_data_186; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_370 = mask_0[2] ? byte_2 : phv_data_185; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_371 = mask_0[3] ? byte_3 : phv_data_184; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_372 = _GEN_8466 == 8'h2e ? _GEN_368 : phv_data_187; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_373 = _GEN_8466 == 8'h2e ? _GEN_369 : phv_data_186; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_374 = _GEN_8466 == 8'h2e ? _GEN_370 : phv_data_185; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_375 = _GEN_8466 == 8'h2e ? _GEN_371 : phv_data_184; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_376 = mask_0[0] ? byte_ : phv_data_191; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_377 = mask_0[1] ? byte_1 : phv_data_190; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_378 = mask_0[2] ? byte_2 : phv_data_189; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_379 = mask_0[3] ? byte_3 : phv_data_188; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_380 = _GEN_8466 == 8'h2f ? _GEN_376 : phv_data_191; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_381 = _GEN_8466 == 8'h2f ? _GEN_377 : phv_data_190; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_382 = _GEN_8466 == 8'h2f ? _GEN_378 : phv_data_189; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_383 = _GEN_8466 == 8'h2f ? _GEN_379 : phv_data_188; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_384 = mask_0[0] ? byte_ : phv_data_195; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_385 = mask_0[1] ? byte_1 : phv_data_194; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_386 = mask_0[2] ? byte_2 : phv_data_193; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_387 = mask_0[3] ? byte_3 : phv_data_192; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_388 = _GEN_8466 == 8'h30 ? _GEN_384 : phv_data_195; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_389 = _GEN_8466 == 8'h30 ? _GEN_385 : phv_data_194; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_390 = _GEN_8466 == 8'h30 ? _GEN_386 : phv_data_193; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_391 = _GEN_8466 == 8'h30 ? _GEN_387 : phv_data_192; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_392 = mask_0[0] ? byte_ : phv_data_199; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_393 = mask_0[1] ? byte_1 : phv_data_198; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_394 = mask_0[2] ? byte_2 : phv_data_197; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_395 = mask_0[3] ? byte_3 : phv_data_196; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_396 = _GEN_8466 == 8'h31 ? _GEN_392 : phv_data_199; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_397 = _GEN_8466 == 8'h31 ? _GEN_393 : phv_data_198; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_398 = _GEN_8466 == 8'h31 ? _GEN_394 : phv_data_197; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_399 = _GEN_8466 == 8'h31 ? _GEN_395 : phv_data_196; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_400 = mask_0[0] ? byte_ : phv_data_203; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_401 = mask_0[1] ? byte_1 : phv_data_202; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_402 = mask_0[2] ? byte_2 : phv_data_201; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_403 = mask_0[3] ? byte_3 : phv_data_200; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_404 = _GEN_8466 == 8'h32 ? _GEN_400 : phv_data_203; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_405 = _GEN_8466 == 8'h32 ? _GEN_401 : phv_data_202; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_406 = _GEN_8466 == 8'h32 ? _GEN_402 : phv_data_201; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_407 = _GEN_8466 == 8'h32 ? _GEN_403 : phv_data_200; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_408 = mask_0[0] ? byte_ : phv_data_207; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_409 = mask_0[1] ? byte_1 : phv_data_206; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_410 = mask_0[2] ? byte_2 : phv_data_205; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_411 = mask_0[3] ? byte_3 : phv_data_204; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_412 = _GEN_8466 == 8'h33 ? _GEN_408 : phv_data_207; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_413 = _GEN_8466 == 8'h33 ? _GEN_409 : phv_data_206; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_414 = _GEN_8466 == 8'h33 ? _GEN_410 : phv_data_205; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_415 = _GEN_8466 == 8'h33 ? _GEN_411 : phv_data_204; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_416 = mask_0[0] ? byte_ : phv_data_211; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_417 = mask_0[1] ? byte_1 : phv_data_210; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_418 = mask_0[2] ? byte_2 : phv_data_209; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_419 = mask_0[3] ? byte_3 : phv_data_208; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_420 = _GEN_8466 == 8'h34 ? _GEN_416 : phv_data_211; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_421 = _GEN_8466 == 8'h34 ? _GEN_417 : phv_data_210; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_422 = _GEN_8466 == 8'h34 ? _GEN_418 : phv_data_209; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_423 = _GEN_8466 == 8'h34 ? _GEN_419 : phv_data_208; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_424 = mask_0[0] ? byte_ : phv_data_215; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_425 = mask_0[1] ? byte_1 : phv_data_214; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_426 = mask_0[2] ? byte_2 : phv_data_213; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_427 = mask_0[3] ? byte_3 : phv_data_212; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_428 = _GEN_8466 == 8'h35 ? _GEN_424 : phv_data_215; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_429 = _GEN_8466 == 8'h35 ? _GEN_425 : phv_data_214; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_430 = _GEN_8466 == 8'h35 ? _GEN_426 : phv_data_213; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_431 = _GEN_8466 == 8'h35 ? _GEN_427 : phv_data_212; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_432 = mask_0[0] ? byte_ : phv_data_219; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_433 = mask_0[1] ? byte_1 : phv_data_218; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_434 = mask_0[2] ? byte_2 : phv_data_217; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_435 = mask_0[3] ? byte_3 : phv_data_216; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_436 = _GEN_8466 == 8'h36 ? _GEN_432 : phv_data_219; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_437 = _GEN_8466 == 8'h36 ? _GEN_433 : phv_data_218; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_438 = _GEN_8466 == 8'h36 ? _GEN_434 : phv_data_217; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_439 = _GEN_8466 == 8'h36 ? _GEN_435 : phv_data_216; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_440 = mask_0[0] ? byte_ : phv_data_223; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_441 = mask_0[1] ? byte_1 : phv_data_222; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_442 = mask_0[2] ? byte_2 : phv_data_221; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_443 = mask_0[3] ? byte_3 : phv_data_220; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_444 = _GEN_8466 == 8'h37 ? _GEN_440 : phv_data_223; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_445 = _GEN_8466 == 8'h37 ? _GEN_441 : phv_data_222; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_446 = _GEN_8466 == 8'h37 ? _GEN_442 : phv_data_221; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_447 = _GEN_8466 == 8'h37 ? _GEN_443 : phv_data_220; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_448 = mask_0[0] ? byte_ : phv_data_227; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_449 = mask_0[1] ? byte_1 : phv_data_226; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_450 = mask_0[2] ? byte_2 : phv_data_225; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_451 = mask_0[3] ? byte_3 : phv_data_224; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_452 = _GEN_8466 == 8'h38 ? _GEN_448 : phv_data_227; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_453 = _GEN_8466 == 8'h38 ? _GEN_449 : phv_data_226; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_454 = _GEN_8466 == 8'h38 ? _GEN_450 : phv_data_225; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_455 = _GEN_8466 == 8'h38 ? _GEN_451 : phv_data_224; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_456 = mask_0[0] ? byte_ : phv_data_231; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_457 = mask_0[1] ? byte_1 : phv_data_230; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_458 = mask_0[2] ? byte_2 : phv_data_229; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_459 = mask_0[3] ? byte_3 : phv_data_228; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_460 = _GEN_8466 == 8'h39 ? _GEN_456 : phv_data_231; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_461 = _GEN_8466 == 8'h39 ? _GEN_457 : phv_data_230; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_462 = _GEN_8466 == 8'h39 ? _GEN_458 : phv_data_229; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_463 = _GEN_8466 == 8'h39 ? _GEN_459 : phv_data_228; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_464 = mask_0[0] ? byte_ : phv_data_235; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_465 = mask_0[1] ? byte_1 : phv_data_234; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_466 = mask_0[2] ? byte_2 : phv_data_233; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_467 = mask_0[3] ? byte_3 : phv_data_232; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_468 = _GEN_8466 == 8'h3a ? _GEN_464 : phv_data_235; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_469 = _GEN_8466 == 8'h3a ? _GEN_465 : phv_data_234; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_470 = _GEN_8466 == 8'h3a ? _GEN_466 : phv_data_233; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_471 = _GEN_8466 == 8'h3a ? _GEN_467 : phv_data_232; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_472 = mask_0[0] ? byte_ : phv_data_239; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_473 = mask_0[1] ? byte_1 : phv_data_238; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_474 = mask_0[2] ? byte_2 : phv_data_237; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_475 = mask_0[3] ? byte_3 : phv_data_236; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_476 = _GEN_8466 == 8'h3b ? _GEN_472 : phv_data_239; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_477 = _GEN_8466 == 8'h3b ? _GEN_473 : phv_data_238; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_478 = _GEN_8466 == 8'h3b ? _GEN_474 : phv_data_237; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_479 = _GEN_8466 == 8'h3b ? _GEN_475 : phv_data_236; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_480 = mask_0[0] ? byte_ : phv_data_243; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_481 = mask_0[1] ? byte_1 : phv_data_242; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_482 = mask_0[2] ? byte_2 : phv_data_241; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_483 = mask_0[3] ? byte_3 : phv_data_240; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_484 = _GEN_8466 == 8'h3c ? _GEN_480 : phv_data_243; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_485 = _GEN_8466 == 8'h3c ? _GEN_481 : phv_data_242; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_486 = _GEN_8466 == 8'h3c ? _GEN_482 : phv_data_241; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_487 = _GEN_8466 == 8'h3c ? _GEN_483 : phv_data_240; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_488 = mask_0[0] ? byte_ : phv_data_247; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_489 = mask_0[1] ? byte_1 : phv_data_246; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_490 = mask_0[2] ? byte_2 : phv_data_245; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_491 = mask_0[3] ? byte_3 : phv_data_244; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_492 = _GEN_8466 == 8'h3d ? _GEN_488 : phv_data_247; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_493 = _GEN_8466 == 8'h3d ? _GEN_489 : phv_data_246; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_494 = _GEN_8466 == 8'h3d ? _GEN_490 : phv_data_245; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_495 = _GEN_8466 == 8'h3d ? _GEN_491 : phv_data_244; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_496 = mask_0[0] ? byte_ : phv_data_251; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_497 = mask_0[1] ? byte_1 : phv_data_250; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_498 = mask_0[2] ? byte_2 : phv_data_249; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_499 = mask_0[3] ? byte_3 : phv_data_248; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_500 = _GEN_8466 == 8'h3e ? _GEN_496 : phv_data_251; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_501 = _GEN_8466 == 8'h3e ? _GEN_497 : phv_data_250; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_502 = _GEN_8466 == 8'h3e ? _GEN_498 : phv_data_249; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_503 = _GEN_8466 == 8'h3e ? _GEN_499 : phv_data_248; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_504 = mask_0[0] ? byte_ : phv_data_255; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_505 = mask_0[1] ? byte_1 : phv_data_254; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_506 = mask_0[2] ? byte_2 : phv_data_253; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_507 = mask_0[3] ? byte_3 : phv_data_252; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_508 = _GEN_8466 == 8'h3f ? _GEN_504 : phv_data_255; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_509 = _GEN_8466 == 8'h3f ? _GEN_505 : phv_data_254; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_510 = _GEN_8466 == 8'h3f ? _GEN_506 : phv_data_253; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_511 = _GEN_8466 == 8'h3f ? _GEN_507 : phv_data_252; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_512 = opcode != 4'h0 ? _GEN_4 : phv_data_3; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_513 = opcode != 4'h0 ? _GEN_5 : phv_data_2; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_514 = opcode != 4'h0 ? _GEN_6 : phv_data_1; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_515 = opcode != 4'h0 ? _GEN_7 : phv_data_0; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_516 = opcode != 4'h0 ? _GEN_12 : phv_data_7; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_517 = opcode != 4'h0 ? _GEN_13 : phv_data_6; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_518 = opcode != 4'h0 ? _GEN_14 : phv_data_5; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_519 = opcode != 4'h0 ? _GEN_15 : phv_data_4; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_520 = opcode != 4'h0 ? _GEN_20 : phv_data_11; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_521 = opcode != 4'h0 ? _GEN_21 : phv_data_10; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_522 = opcode != 4'h0 ? _GEN_22 : phv_data_9; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_523 = opcode != 4'h0 ? _GEN_23 : phv_data_8; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_524 = opcode != 4'h0 ? _GEN_28 : phv_data_15; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_525 = opcode != 4'h0 ? _GEN_29 : phv_data_14; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_526 = opcode != 4'h0 ? _GEN_30 : phv_data_13; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_527 = opcode != 4'h0 ? _GEN_31 : phv_data_12; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_528 = opcode != 4'h0 ? _GEN_36 : phv_data_19; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_529 = opcode != 4'h0 ? _GEN_37 : phv_data_18; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_530 = opcode != 4'h0 ? _GEN_38 : phv_data_17; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_531 = opcode != 4'h0 ? _GEN_39 : phv_data_16; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_532 = opcode != 4'h0 ? _GEN_44 : phv_data_23; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_533 = opcode != 4'h0 ? _GEN_45 : phv_data_22; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_534 = opcode != 4'h0 ? _GEN_46 : phv_data_21; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_535 = opcode != 4'h0 ? _GEN_47 : phv_data_20; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_536 = opcode != 4'h0 ? _GEN_52 : phv_data_27; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_537 = opcode != 4'h0 ? _GEN_53 : phv_data_26; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_538 = opcode != 4'h0 ? _GEN_54 : phv_data_25; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_539 = opcode != 4'h0 ? _GEN_55 : phv_data_24; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_540 = opcode != 4'h0 ? _GEN_60 : phv_data_31; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_541 = opcode != 4'h0 ? _GEN_61 : phv_data_30; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_542 = opcode != 4'h0 ? _GEN_62 : phv_data_29; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_543 = opcode != 4'h0 ? _GEN_63 : phv_data_28; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_544 = opcode != 4'h0 ? _GEN_68 : phv_data_35; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_545 = opcode != 4'h0 ? _GEN_69 : phv_data_34; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_546 = opcode != 4'h0 ? _GEN_70 : phv_data_33; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_547 = opcode != 4'h0 ? _GEN_71 : phv_data_32; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_548 = opcode != 4'h0 ? _GEN_76 : phv_data_39; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_549 = opcode != 4'h0 ? _GEN_77 : phv_data_38; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_550 = opcode != 4'h0 ? _GEN_78 : phv_data_37; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_551 = opcode != 4'h0 ? _GEN_79 : phv_data_36; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_552 = opcode != 4'h0 ? _GEN_84 : phv_data_43; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_553 = opcode != 4'h0 ? _GEN_85 : phv_data_42; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_554 = opcode != 4'h0 ? _GEN_86 : phv_data_41; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_555 = opcode != 4'h0 ? _GEN_87 : phv_data_40; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_556 = opcode != 4'h0 ? _GEN_92 : phv_data_47; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_557 = opcode != 4'h0 ? _GEN_93 : phv_data_46; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_558 = opcode != 4'h0 ? _GEN_94 : phv_data_45; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_559 = opcode != 4'h0 ? _GEN_95 : phv_data_44; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_560 = opcode != 4'h0 ? _GEN_100 : phv_data_51; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_561 = opcode != 4'h0 ? _GEN_101 : phv_data_50; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_562 = opcode != 4'h0 ? _GEN_102 : phv_data_49; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_563 = opcode != 4'h0 ? _GEN_103 : phv_data_48; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_564 = opcode != 4'h0 ? _GEN_108 : phv_data_55; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_565 = opcode != 4'h0 ? _GEN_109 : phv_data_54; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_566 = opcode != 4'h0 ? _GEN_110 : phv_data_53; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_567 = opcode != 4'h0 ? _GEN_111 : phv_data_52; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_568 = opcode != 4'h0 ? _GEN_116 : phv_data_59; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_569 = opcode != 4'h0 ? _GEN_117 : phv_data_58; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_570 = opcode != 4'h0 ? _GEN_118 : phv_data_57; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_571 = opcode != 4'h0 ? _GEN_119 : phv_data_56; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_572 = opcode != 4'h0 ? _GEN_124 : phv_data_63; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_573 = opcode != 4'h0 ? _GEN_125 : phv_data_62; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_574 = opcode != 4'h0 ? _GEN_126 : phv_data_61; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_575 = opcode != 4'h0 ? _GEN_127 : phv_data_60; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_576 = opcode != 4'h0 ? _GEN_132 : phv_data_67; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_577 = opcode != 4'h0 ? _GEN_133 : phv_data_66; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_578 = opcode != 4'h0 ? _GEN_134 : phv_data_65; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_579 = opcode != 4'h0 ? _GEN_135 : phv_data_64; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_580 = opcode != 4'h0 ? _GEN_140 : phv_data_71; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_581 = opcode != 4'h0 ? _GEN_141 : phv_data_70; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_582 = opcode != 4'h0 ? _GEN_142 : phv_data_69; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_583 = opcode != 4'h0 ? _GEN_143 : phv_data_68; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_584 = opcode != 4'h0 ? _GEN_148 : phv_data_75; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_585 = opcode != 4'h0 ? _GEN_149 : phv_data_74; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_586 = opcode != 4'h0 ? _GEN_150 : phv_data_73; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_587 = opcode != 4'h0 ? _GEN_151 : phv_data_72; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_588 = opcode != 4'h0 ? _GEN_156 : phv_data_79; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_589 = opcode != 4'h0 ? _GEN_157 : phv_data_78; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_590 = opcode != 4'h0 ? _GEN_158 : phv_data_77; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_591 = opcode != 4'h0 ? _GEN_159 : phv_data_76; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_592 = opcode != 4'h0 ? _GEN_164 : phv_data_83; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_593 = opcode != 4'h0 ? _GEN_165 : phv_data_82; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_594 = opcode != 4'h0 ? _GEN_166 : phv_data_81; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_595 = opcode != 4'h0 ? _GEN_167 : phv_data_80; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_596 = opcode != 4'h0 ? _GEN_172 : phv_data_87; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_597 = opcode != 4'h0 ? _GEN_173 : phv_data_86; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_598 = opcode != 4'h0 ? _GEN_174 : phv_data_85; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_599 = opcode != 4'h0 ? _GEN_175 : phv_data_84; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_600 = opcode != 4'h0 ? _GEN_180 : phv_data_91; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_601 = opcode != 4'h0 ? _GEN_181 : phv_data_90; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_602 = opcode != 4'h0 ? _GEN_182 : phv_data_89; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_603 = opcode != 4'h0 ? _GEN_183 : phv_data_88; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_604 = opcode != 4'h0 ? _GEN_188 : phv_data_95; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_605 = opcode != 4'h0 ? _GEN_189 : phv_data_94; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_606 = opcode != 4'h0 ? _GEN_190 : phv_data_93; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_607 = opcode != 4'h0 ? _GEN_191 : phv_data_92; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_608 = opcode != 4'h0 ? _GEN_196 : phv_data_99; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_609 = opcode != 4'h0 ? _GEN_197 : phv_data_98; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_610 = opcode != 4'h0 ? _GEN_198 : phv_data_97; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_611 = opcode != 4'h0 ? _GEN_199 : phv_data_96; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_612 = opcode != 4'h0 ? _GEN_204 : phv_data_103; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_613 = opcode != 4'h0 ? _GEN_205 : phv_data_102; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_614 = opcode != 4'h0 ? _GEN_206 : phv_data_101; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_615 = opcode != 4'h0 ? _GEN_207 : phv_data_100; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_616 = opcode != 4'h0 ? _GEN_212 : phv_data_107; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_617 = opcode != 4'h0 ? _GEN_213 : phv_data_106; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_618 = opcode != 4'h0 ? _GEN_214 : phv_data_105; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_619 = opcode != 4'h0 ? _GEN_215 : phv_data_104; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_620 = opcode != 4'h0 ? _GEN_220 : phv_data_111; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_621 = opcode != 4'h0 ? _GEN_221 : phv_data_110; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_622 = opcode != 4'h0 ? _GEN_222 : phv_data_109; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_623 = opcode != 4'h0 ? _GEN_223 : phv_data_108; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_624 = opcode != 4'h0 ? _GEN_228 : phv_data_115; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_625 = opcode != 4'h0 ? _GEN_229 : phv_data_114; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_626 = opcode != 4'h0 ? _GEN_230 : phv_data_113; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_627 = opcode != 4'h0 ? _GEN_231 : phv_data_112; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_628 = opcode != 4'h0 ? _GEN_236 : phv_data_119; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_629 = opcode != 4'h0 ? _GEN_237 : phv_data_118; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_630 = opcode != 4'h0 ? _GEN_238 : phv_data_117; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_631 = opcode != 4'h0 ? _GEN_239 : phv_data_116; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_632 = opcode != 4'h0 ? _GEN_244 : phv_data_123; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_633 = opcode != 4'h0 ? _GEN_245 : phv_data_122; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_634 = opcode != 4'h0 ? _GEN_246 : phv_data_121; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_635 = opcode != 4'h0 ? _GEN_247 : phv_data_120; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_636 = opcode != 4'h0 ? _GEN_252 : phv_data_127; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_637 = opcode != 4'h0 ? _GEN_253 : phv_data_126; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_638 = opcode != 4'h0 ? _GEN_254 : phv_data_125; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_639 = opcode != 4'h0 ? _GEN_255 : phv_data_124; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_640 = opcode != 4'h0 ? _GEN_260 : phv_data_131; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_641 = opcode != 4'h0 ? _GEN_261 : phv_data_130; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_642 = opcode != 4'h0 ? _GEN_262 : phv_data_129; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_643 = opcode != 4'h0 ? _GEN_263 : phv_data_128; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_644 = opcode != 4'h0 ? _GEN_268 : phv_data_135; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_645 = opcode != 4'h0 ? _GEN_269 : phv_data_134; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_646 = opcode != 4'h0 ? _GEN_270 : phv_data_133; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_647 = opcode != 4'h0 ? _GEN_271 : phv_data_132; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_648 = opcode != 4'h0 ? _GEN_276 : phv_data_139; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_649 = opcode != 4'h0 ? _GEN_277 : phv_data_138; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_650 = opcode != 4'h0 ? _GEN_278 : phv_data_137; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_651 = opcode != 4'h0 ? _GEN_279 : phv_data_136; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_652 = opcode != 4'h0 ? _GEN_284 : phv_data_143; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_653 = opcode != 4'h0 ? _GEN_285 : phv_data_142; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_654 = opcode != 4'h0 ? _GEN_286 : phv_data_141; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_655 = opcode != 4'h0 ? _GEN_287 : phv_data_140; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_656 = opcode != 4'h0 ? _GEN_292 : phv_data_147; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_657 = opcode != 4'h0 ? _GEN_293 : phv_data_146; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_658 = opcode != 4'h0 ? _GEN_294 : phv_data_145; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_659 = opcode != 4'h0 ? _GEN_295 : phv_data_144; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_660 = opcode != 4'h0 ? _GEN_300 : phv_data_151; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_661 = opcode != 4'h0 ? _GEN_301 : phv_data_150; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_662 = opcode != 4'h0 ? _GEN_302 : phv_data_149; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_663 = opcode != 4'h0 ? _GEN_303 : phv_data_148; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_664 = opcode != 4'h0 ? _GEN_308 : phv_data_155; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_665 = opcode != 4'h0 ? _GEN_309 : phv_data_154; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_666 = opcode != 4'h0 ? _GEN_310 : phv_data_153; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_667 = opcode != 4'h0 ? _GEN_311 : phv_data_152; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_668 = opcode != 4'h0 ? _GEN_316 : phv_data_159; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_669 = opcode != 4'h0 ? _GEN_317 : phv_data_158; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_670 = opcode != 4'h0 ? _GEN_318 : phv_data_157; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_671 = opcode != 4'h0 ? _GEN_319 : phv_data_156; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_672 = opcode != 4'h0 ? _GEN_324 : phv_data_163; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_673 = opcode != 4'h0 ? _GEN_325 : phv_data_162; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_674 = opcode != 4'h0 ? _GEN_326 : phv_data_161; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_675 = opcode != 4'h0 ? _GEN_327 : phv_data_160; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_676 = opcode != 4'h0 ? _GEN_332 : phv_data_167; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_677 = opcode != 4'h0 ? _GEN_333 : phv_data_166; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_678 = opcode != 4'h0 ? _GEN_334 : phv_data_165; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_679 = opcode != 4'h0 ? _GEN_335 : phv_data_164; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_680 = opcode != 4'h0 ? _GEN_340 : phv_data_171; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_681 = opcode != 4'h0 ? _GEN_341 : phv_data_170; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_682 = opcode != 4'h0 ? _GEN_342 : phv_data_169; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_683 = opcode != 4'h0 ? _GEN_343 : phv_data_168; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_684 = opcode != 4'h0 ? _GEN_348 : phv_data_175; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_685 = opcode != 4'h0 ? _GEN_349 : phv_data_174; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_686 = opcode != 4'h0 ? _GEN_350 : phv_data_173; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_687 = opcode != 4'h0 ? _GEN_351 : phv_data_172; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_688 = opcode != 4'h0 ? _GEN_356 : phv_data_179; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_689 = opcode != 4'h0 ? _GEN_357 : phv_data_178; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_690 = opcode != 4'h0 ? _GEN_358 : phv_data_177; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_691 = opcode != 4'h0 ? _GEN_359 : phv_data_176; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_692 = opcode != 4'h0 ? _GEN_364 : phv_data_183; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_693 = opcode != 4'h0 ? _GEN_365 : phv_data_182; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_694 = opcode != 4'h0 ? _GEN_366 : phv_data_181; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_695 = opcode != 4'h0 ? _GEN_367 : phv_data_180; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_696 = opcode != 4'h0 ? _GEN_372 : phv_data_187; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_697 = opcode != 4'h0 ? _GEN_373 : phv_data_186; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_698 = opcode != 4'h0 ? _GEN_374 : phv_data_185; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_699 = opcode != 4'h0 ? _GEN_375 : phv_data_184; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_700 = opcode != 4'h0 ? _GEN_380 : phv_data_191; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_701 = opcode != 4'h0 ? _GEN_381 : phv_data_190; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_702 = opcode != 4'h0 ? _GEN_382 : phv_data_189; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_703 = opcode != 4'h0 ? _GEN_383 : phv_data_188; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_704 = opcode != 4'h0 ? _GEN_388 : phv_data_195; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_705 = opcode != 4'h0 ? _GEN_389 : phv_data_194; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_706 = opcode != 4'h0 ? _GEN_390 : phv_data_193; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_707 = opcode != 4'h0 ? _GEN_391 : phv_data_192; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_708 = opcode != 4'h0 ? _GEN_396 : phv_data_199; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_709 = opcode != 4'h0 ? _GEN_397 : phv_data_198; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_710 = opcode != 4'h0 ? _GEN_398 : phv_data_197; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_711 = opcode != 4'h0 ? _GEN_399 : phv_data_196; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_712 = opcode != 4'h0 ? _GEN_404 : phv_data_203; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_713 = opcode != 4'h0 ? _GEN_405 : phv_data_202; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_714 = opcode != 4'h0 ? _GEN_406 : phv_data_201; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_715 = opcode != 4'h0 ? _GEN_407 : phv_data_200; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_716 = opcode != 4'h0 ? _GEN_412 : phv_data_207; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_717 = opcode != 4'h0 ? _GEN_413 : phv_data_206; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_718 = opcode != 4'h0 ? _GEN_414 : phv_data_205; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_719 = opcode != 4'h0 ? _GEN_415 : phv_data_204; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_720 = opcode != 4'h0 ? _GEN_420 : phv_data_211; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_721 = opcode != 4'h0 ? _GEN_421 : phv_data_210; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_722 = opcode != 4'h0 ? _GEN_422 : phv_data_209; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_723 = opcode != 4'h0 ? _GEN_423 : phv_data_208; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_724 = opcode != 4'h0 ? _GEN_428 : phv_data_215; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_725 = opcode != 4'h0 ? _GEN_429 : phv_data_214; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_726 = opcode != 4'h0 ? _GEN_430 : phv_data_213; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_727 = opcode != 4'h0 ? _GEN_431 : phv_data_212; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_728 = opcode != 4'h0 ? _GEN_436 : phv_data_219; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_729 = opcode != 4'h0 ? _GEN_437 : phv_data_218; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_730 = opcode != 4'h0 ? _GEN_438 : phv_data_217; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_731 = opcode != 4'h0 ? _GEN_439 : phv_data_216; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_732 = opcode != 4'h0 ? _GEN_444 : phv_data_223; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_733 = opcode != 4'h0 ? _GEN_445 : phv_data_222; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_734 = opcode != 4'h0 ? _GEN_446 : phv_data_221; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_735 = opcode != 4'h0 ? _GEN_447 : phv_data_220; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_736 = opcode != 4'h0 ? _GEN_452 : phv_data_227; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_737 = opcode != 4'h0 ? _GEN_453 : phv_data_226; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_738 = opcode != 4'h0 ? _GEN_454 : phv_data_225; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_739 = opcode != 4'h0 ? _GEN_455 : phv_data_224; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_740 = opcode != 4'h0 ? _GEN_460 : phv_data_231; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_741 = opcode != 4'h0 ? _GEN_461 : phv_data_230; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_742 = opcode != 4'h0 ? _GEN_462 : phv_data_229; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_743 = opcode != 4'h0 ? _GEN_463 : phv_data_228; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_744 = opcode != 4'h0 ? _GEN_468 : phv_data_235; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_745 = opcode != 4'h0 ? _GEN_469 : phv_data_234; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_746 = opcode != 4'h0 ? _GEN_470 : phv_data_233; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_747 = opcode != 4'h0 ? _GEN_471 : phv_data_232; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_748 = opcode != 4'h0 ? _GEN_476 : phv_data_239; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_749 = opcode != 4'h0 ? _GEN_477 : phv_data_238; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_750 = opcode != 4'h0 ? _GEN_478 : phv_data_237; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_751 = opcode != 4'h0 ? _GEN_479 : phv_data_236; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_752 = opcode != 4'h0 ? _GEN_484 : phv_data_243; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_753 = opcode != 4'h0 ? _GEN_485 : phv_data_242; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_754 = opcode != 4'h0 ? _GEN_486 : phv_data_241; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_755 = opcode != 4'h0 ? _GEN_487 : phv_data_240; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_756 = opcode != 4'h0 ? _GEN_492 : phv_data_247; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_757 = opcode != 4'h0 ? _GEN_493 : phv_data_246; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_758 = opcode != 4'h0 ? _GEN_494 : phv_data_245; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_759 = opcode != 4'h0 ? _GEN_495 : phv_data_244; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_760 = opcode != 4'h0 ? _GEN_500 : phv_data_251; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_761 = opcode != 4'h0 ? _GEN_501 : phv_data_250; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_762 = opcode != 4'h0 ? _GEN_502 : phv_data_249; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_763 = opcode != 4'h0 ? _GEN_503 : phv_data_248; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_764 = opcode != 4'h0 ? _GEN_508 : phv_data_255; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_765 = opcode != 4'h0 ? _GEN_509 : phv_data_254; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_766 = opcode != 4'h0 ? _GEN_510 : phv_data_253; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_767 = opcode != 4'h0 ? _GEN_511 : phv_data_252; // @[executor.scala 470:55 executor.scala 450:25]
  wire [3:0] _GEN_768 = opcode == 4'hf ? parameter_2[13:10] : phv_next_processor_id; // @[executor.scala 466:52 executor.scala 467:55 executor.scala 450:25]
  wire  _GEN_769 = opcode == 4'hf ? parameter_2[0] : phv_next_config_id; // @[executor.scala 466:52 executor.scala 468:55 executor.scala 450:25]
  wire [7:0] _GEN_770 = opcode == 4'hf ? phv_data_3 : _GEN_512; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_771 = opcode == 4'hf ? phv_data_2 : _GEN_513; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_772 = opcode == 4'hf ? phv_data_1 : _GEN_514; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_773 = opcode == 4'hf ? phv_data_0 : _GEN_515; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_774 = opcode == 4'hf ? phv_data_7 : _GEN_516; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_775 = opcode == 4'hf ? phv_data_6 : _GEN_517; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_776 = opcode == 4'hf ? phv_data_5 : _GEN_518; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_777 = opcode == 4'hf ? phv_data_4 : _GEN_519; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_778 = opcode == 4'hf ? phv_data_11 : _GEN_520; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_779 = opcode == 4'hf ? phv_data_10 : _GEN_521; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_780 = opcode == 4'hf ? phv_data_9 : _GEN_522; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_781 = opcode == 4'hf ? phv_data_8 : _GEN_523; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_782 = opcode == 4'hf ? phv_data_15 : _GEN_524; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_783 = opcode == 4'hf ? phv_data_14 : _GEN_525; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_784 = opcode == 4'hf ? phv_data_13 : _GEN_526; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_785 = opcode == 4'hf ? phv_data_12 : _GEN_527; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_786 = opcode == 4'hf ? phv_data_19 : _GEN_528; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_787 = opcode == 4'hf ? phv_data_18 : _GEN_529; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_788 = opcode == 4'hf ? phv_data_17 : _GEN_530; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_789 = opcode == 4'hf ? phv_data_16 : _GEN_531; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_790 = opcode == 4'hf ? phv_data_23 : _GEN_532; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_791 = opcode == 4'hf ? phv_data_22 : _GEN_533; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_792 = opcode == 4'hf ? phv_data_21 : _GEN_534; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_793 = opcode == 4'hf ? phv_data_20 : _GEN_535; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_794 = opcode == 4'hf ? phv_data_27 : _GEN_536; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_795 = opcode == 4'hf ? phv_data_26 : _GEN_537; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_796 = opcode == 4'hf ? phv_data_25 : _GEN_538; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_797 = opcode == 4'hf ? phv_data_24 : _GEN_539; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_798 = opcode == 4'hf ? phv_data_31 : _GEN_540; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_799 = opcode == 4'hf ? phv_data_30 : _GEN_541; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_800 = opcode == 4'hf ? phv_data_29 : _GEN_542; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_801 = opcode == 4'hf ? phv_data_28 : _GEN_543; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_802 = opcode == 4'hf ? phv_data_35 : _GEN_544; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_803 = opcode == 4'hf ? phv_data_34 : _GEN_545; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_804 = opcode == 4'hf ? phv_data_33 : _GEN_546; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_805 = opcode == 4'hf ? phv_data_32 : _GEN_547; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_806 = opcode == 4'hf ? phv_data_39 : _GEN_548; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_807 = opcode == 4'hf ? phv_data_38 : _GEN_549; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_808 = opcode == 4'hf ? phv_data_37 : _GEN_550; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_809 = opcode == 4'hf ? phv_data_36 : _GEN_551; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_810 = opcode == 4'hf ? phv_data_43 : _GEN_552; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_811 = opcode == 4'hf ? phv_data_42 : _GEN_553; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_812 = opcode == 4'hf ? phv_data_41 : _GEN_554; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_813 = opcode == 4'hf ? phv_data_40 : _GEN_555; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_814 = opcode == 4'hf ? phv_data_47 : _GEN_556; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_815 = opcode == 4'hf ? phv_data_46 : _GEN_557; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_816 = opcode == 4'hf ? phv_data_45 : _GEN_558; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_817 = opcode == 4'hf ? phv_data_44 : _GEN_559; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_818 = opcode == 4'hf ? phv_data_51 : _GEN_560; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_819 = opcode == 4'hf ? phv_data_50 : _GEN_561; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_820 = opcode == 4'hf ? phv_data_49 : _GEN_562; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_821 = opcode == 4'hf ? phv_data_48 : _GEN_563; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_822 = opcode == 4'hf ? phv_data_55 : _GEN_564; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_823 = opcode == 4'hf ? phv_data_54 : _GEN_565; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_824 = opcode == 4'hf ? phv_data_53 : _GEN_566; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_825 = opcode == 4'hf ? phv_data_52 : _GEN_567; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_826 = opcode == 4'hf ? phv_data_59 : _GEN_568; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_827 = opcode == 4'hf ? phv_data_58 : _GEN_569; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_828 = opcode == 4'hf ? phv_data_57 : _GEN_570; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_829 = opcode == 4'hf ? phv_data_56 : _GEN_571; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_830 = opcode == 4'hf ? phv_data_63 : _GEN_572; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_831 = opcode == 4'hf ? phv_data_62 : _GEN_573; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_832 = opcode == 4'hf ? phv_data_61 : _GEN_574; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_833 = opcode == 4'hf ? phv_data_60 : _GEN_575; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_834 = opcode == 4'hf ? phv_data_67 : _GEN_576; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_835 = opcode == 4'hf ? phv_data_66 : _GEN_577; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_836 = opcode == 4'hf ? phv_data_65 : _GEN_578; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_837 = opcode == 4'hf ? phv_data_64 : _GEN_579; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_838 = opcode == 4'hf ? phv_data_71 : _GEN_580; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_839 = opcode == 4'hf ? phv_data_70 : _GEN_581; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_840 = opcode == 4'hf ? phv_data_69 : _GEN_582; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_841 = opcode == 4'hf ? phv_data_68 : _GEN_583; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_842 = opcode == 4'hf ? phv_data_75 : _GEN_584; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_843 = opcode == 4'hf ? phv_data_74 : _GEN_585; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_844 = opcode == 4'hf ? phv_data_73 : _GEN_586; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_845 = opcode == 4'hf ? phv_data_72 : _GEN_587; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_846 = opcode == 4'hf ? phv_data_79 : _GEN_588; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_847 = opcode == 4'hf ? phv_data_78 : _GEN_589; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_848 = opcode == 4'hf ? phv_data_77 : _GEN_590; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_849 = opcode == 4'hf ? phv_data_76 : _GEN_591; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_850 = opcode == 4'hf ? phv_data_83 : _GEN_592; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_851 = opcode == 4'hf ? phv_data_82 : _GEN_593; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_852 = opcode == 4'hf ? phv_data_81 : _GEN_594; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_853 = opcode == 4'hf ? phv_data_80 : _GEN_595; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_854 = opcode == 4'hf ? phv_data_87 : _GEN_596; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_855 = opcode == 4'hf ? phv_data_86 : _GEN_597; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_856 = opcode == 4'hf ? phv_data_85 : _GEN_598; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_857 = opcode == 4'hf ? phv_data_84 : _GEN_599; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_858 = opcode == 4'hf ? phv_data_91 : _GEN_600; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_859 = opcode == 4'hf ? phv_data_90 : _GEN_601; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_860 = opcode == 4'hf ? phv_data_89 : _GEN_602; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_861 = opcode == 4'hf ? phv_data_88 : _GEN_603; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_862 = opcode == 4'hf ? phv_data_95 : _GEN_604; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_863 = opcode == 4'hf ? phv_data_94 : _GEN_605; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_864 = opcode == 4'hf ? phv_data_93 : _GEN_606; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_865 = opcode == 4'hf ? phv_data_92 : _GEN_607; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_866 = opcode == 4'hf ? phv_data_99 : _GEN_608; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_867 = opcode == 4'hf ? phv_data_98 : _GEN_609; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_868 = opcode == 4'hf ? phv_data_97 : _GEN_610; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_869 = opcode == 4'hf ? phv_data_96 : _GEN_611; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_870 = opcode == 4'hf ? phv_data_103 : _GEN_612; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_871 = opcode == 4'hf ? phv_data_102 : _GEN_613; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_872 = opcode == 4'hf ? phv_data_101 : _GEN_614; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_873 = opcode == 4'hf ? phv_data_100 : _GEN_615; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_874 = opcode == 4'hf ? phv_data_107 : _GEN_616; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_875 = opcode == 4'hf ? phv_data_106 : _GEN_617; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_876 = opcode == 4'hf ? phv_data_105 : _GEN_618; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_877 = opcode == 4'hf ? phv_data_104 : _GEN_619; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_878 = opcode == 4'hf ? phv_data_111 : _GEN_620; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_879 = opcode == 4'hf ? phv_data_110 : _GEN_621; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_880 = opcode == 4'hf ? phv_data_109 : _GEN_622; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_881 = opcode == 4'hf ? phv_data_108 : _GEN_623; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_882 = opcode == 4'hf ? phv_data_115 : _GEN_624; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_883 = opcode == 4'hf ? phv_data_114 : _GEN_625; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_884 = opcode == 4'hf ? phv_data_113 : _GEN_626; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_885 = opcode == 4'hf ? phv_data_112 : _GEN_627; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_886 = opcode == 4'hf ? phv_data_119 : _GEN_628; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_887 = opcode == 4'hf ? phv_data_118 : _GEN_629; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_888 = opcode == 4'hf ? phv_data_117 : _GEN_630; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_889 = opcode == 4'hf ? phv_data_116 : _GEN_631; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_890 = opcode == 4'hf ? phv_data_123 : _GEN_632; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_891 = opcode == 4'hf ? phv_data_122 : _GEN_633; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_892 = opcode == 4'hf ? phv_data_121 : _GEN_634; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_893 = opcode == 4'hf ? phv_data_120 : _GEN_635; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_894 = opcode == 4'hf ? phv_data_127 : _GEN_636; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_895 = opcode == 4'hf ? phv_data_126 : _GEN_637; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_896 = opcode == 4'hf ? phv_data_125 : _GEN_638; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_897 = opcode == 4'hf ? phv_data_124 : _GEN_639; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_898 = opcode == 4'hf ? phv_data_131 : _GEN_640; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_899 = opcode == 4'hf ? phv_data_130 : _GEN_641; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_900 = opcode == 4'hf ? phv_data_129 : _GEN_642; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_901 = opcode == 4'hf ? phv_data_128 : _GEN_643; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_902 = opcode == 4'hf ? phv_data_135 : _GEN_644; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_903 = opcode == 4'hf ? phv_data_134 : _GEN_645; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_904 = opcode == 4'hf ? phv_data_133 : _GEN_646; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_905 = opcode == 4'hf ? phv_data_132 : _GEN_647; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_906 = opcode == 4'hf ? phv_data_139 : _GEN_648; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_907 = opcode == 4'hf ? phv_data_138 : _GEN_649; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_908 = opcode == 4'hf ? phv_data_137 : _GEN_650; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_909 = opcode == 4'hf ? phv_data_136 : _GEN_651; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_910 = opcode == 4'hf ? phv_data_143 : _GEN_652; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_911 = opcode == 4'hf ? phv_data_142 : _GEN_653; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_912 = opcode == 4'hf ? phv_data_141 : _GEN_654; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_913 = opcode == 4'hf ? phv_data_140 : _GEN_655; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_914 = opcode == 4'hf ? phv_data_147 : _GEN_656; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_915 = opcode == 4'hf ? phv_data_146 : _GEN_657; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_916 = opcode == 4'hf ? phv_data_145 : _GEN_658; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_917 = opcode == 4'hf ? phv_data_144 : _GEN_659; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_918 = opcode == 4'hf ? phv_data_151 : _GEN_660; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_919 = opcode == 4'hf ? phv_data_150 : _GEN_661; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_920 = opcode == 4'hf ? phv_data_149 : _GEN_662; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_921 = opcode == 4'hf ? phv_data_148 : _GEN_663; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_922 = opcode == 4'hf ? phv_data_155 : _GEN_664; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_923 = opcode == 4'hf ? phv_data_154 : _GEN_665; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_924 = opcode == 4'hf ? phv_data_153 : _GEN_666; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_925 = opcode == 4'hf ? phv_data_152 : _GEN_667; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_926 = opcode == 4'hf ? phv_data_159 : _GEN_668; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_927 = opcode == 4'hf ? phv_data_158 : _GEN_669; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_928 = opcode == 4'hf ? phv_data_157 : _GEN_670; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_929 = opcode == 4'hf ? phv_data_156 : _GEN_671; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_930 = opcode == 4'hf ? phv_data_163 : _GEN_672; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_931 = opcode == 4'hf ? phv_data_162 : _GEN_673; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_932 = opcode == 4'hf ? phv_data_161 : _GEN_674; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_933 = opcode == 4'hf ? phv_data_160 : _GEN_675; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_934 = opcode == 4'hf ? phv_data_167 : _GEN_676; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_935 = opcode == 4'hf ? phv_data_166 : _GEN_677; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_936 = opcode == 4'hf ? phv_data_165 : _GEN_678; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_937 = opcode == 4'hf ? phv_data_164 : _GEN_679; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_938 = opcode == 4'hf ? phv_data_171 : _GEN_680; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_939 = opcode == 4'hf ? phv_data_170 : _GEN_681; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_940 = opcode == 4'hf ? phv_data_169 : _GEN_682; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_941 = opcode == 4'hf ? phv_data_168 : _GEN_683; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_942 = opcode == 4'hf ? phv_data_175 : _GEN_684; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_943 = opcode == 4'hf ? phv_data_174 : _GEN_685; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_944 = opcode == 4'hf ? phv_data_173 : _GEN_686; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_945 = opcode == 4'hf ? phv_data_172 : _GEN_687; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_946 = opcode == 4'hf ? phv_data_179 : _GEN_688; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_947 = opcode == 4'hf ? phv_data_178 : _GEN_689; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_948 = opcode == 4'hf ? phv_data_177 : _GEN_690; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_949 = opcode == 4'hf ? phv_data_176 : _GEN_691; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_950 = opcode == 4'hf ? phv_data_183 : _GEN_692; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_951 = opcode == 4'hf ? phv_data_182 : _GEN_693; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_952 = opcode == 4'hf ? phv_data_181 : _GEN_694; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_953 = opcode == 4'hf ? phv_data_180 : _GEN_695; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_954 = opcode == 4'hf ? phv_data_187 : _GEN_696; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_955 = opcode == 4'hf ? phv_data_186 : _GEN_697; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_956 = opcode == 4'hf ? phv_data_185 : _GEN_698; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_957 = opcode == 4'hf ? phv_data_184 : _GEN_699; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_958 = opcode == 4'hf ? phv_data_191 : _GEN_700; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_959 = opcode == 4'hf ? phv_data_190 : _GEN_701; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_960 = opcode == 4'hf ? phv_data_189 : _GEN_702; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_961 = opcode == 4'hf ? phv_data_188 : _GEN_703; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_962 = opcode == 4'hf ? phv_data_195 : _GEN_704; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_963 = opcode == 4'hf ? phv_data_194 : _GEN_705; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_964 = opcode == 4'hf ? phv_data_193 : _GEN_706; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_965 = opcode == 4'hf ? phv_data_192 : _GEN_707; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_966 = opcode == 4'hf ? phv_data_199 : _GEN_708; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_967 = opcode == 4'hf ? phv_data_198 : _GEN_709; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_968 = opcode == 4'hf ? phv_data_197 : _GEN_710; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_969 = opcode == 4'hf ? phv_data_196 : _GEN_711; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_970 = opcode == 4'hf ? phv_data_203 : _GEN_712; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_971 = opcode == 4'hf ? phv_data_202 : _GEN_713; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_972 = opcode == 4'hf ? phv_data_201 : _GEN_714; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_973 = opcode == 4'hf ? phv_data_200 : _GEN_715; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_974 = opcode == 4'hf ? phv_data_207 : _GEN_716; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_975 = opcode == 4'hf ? phv_data_206 : _GEN_717; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_976 = opcode == 4'hf ? phv_data_205 : _GEN_718; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_977 = opcode == 4'hf ? phv_data_204 : _GEN_719; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_978 = opcode == 4'hf ? phv_data_211 : _GEN_720; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_979 = opcode == 4'hf ? phv_data_210 : _GEN_721; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_980 = opcode == 4'hf ? phv_data_209 : _GEN_722; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_981 = opcode == 4'hf ? phv_data_208 : _GEN_723; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_982 = opcode == 4'hf ? phv_data_215 : _GEN_724; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_983 = opcode == 4'hf ? phv_data_214 : _GEN_725; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_984 = opcode == 4'hf ? phv_data_213 : _GEN_726; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_985 = opcode == 4'hf ? phv_data_212 : _GEN_727; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_986 = opcode == 4'hf ? phv_data_219 : _GEN_728; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_987 = opcode == 4'hf ? phv_data_218 : _GEN_729; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_988 = opcode == 4'hf ? phv_data_217 : _GEN_730; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_989 = opcode == 4'hf ? phv_data_216 : _GEN_731; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_990 = opcode == 4'hf ? phv_data_223 : _GEN_732; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_991 = opcode == 4'hf ? phv_data_222 : _GEN_733; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_992 = opcode == 4'hf ? phv_data_221 : _GEN_734; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_993 = opcode == 4'hf ? phv_data_220 : _GEN_735; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_994 = opcode == 4'hf ? phv_data_227 : _GEN_736; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_995 = opcode == 4'hf ? phv_data_226 : _GEN_737; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_996 = opcode == 4'hf ? phv_data_225 : _GEN_738; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_997 = opcode == 4'hf ? phv_data_224 : _GEN_739; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_998 = opcode == 4'hf ? phv_data_231 : _GEN_740; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_999 = opcode == 4'hf ? phv_data_230 : _GEN_741; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1000 = opcode == 4'hf ? phv_data_229 : _GEN_742; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1001 = opcode == 4'hf ? phv_data_228 : _GEN_743; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1002 = opcode == 4'hf ? phv_data_235 : _GEN_744; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1003 = opcode == 4'hf ? phv_data_234 : _GEN_745; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1004 = opcode == 4'hf ? phv_data_233 : _GEN_746; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1005 = opcode == 4'hf ? phv_data_232 : _GEN_747; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1006 = opcode == 4'hf ? phv_data_239 : _GEN_748; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1007 = opcode == 4'hf ? phv_data_238 : _GEN_749; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1008 = opcode == 4'hf ? phv_data_237 : _GEN_750; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1009 = opcode == 4'hf ? phv_data_236 : _GEN_751; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1010 = opcode == 4'hf ? phv_data_243 : _GEN_752; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1011 = opcode == 4'hf ? phv_data_242 : _GEN_753; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1012 = opcode == 4'hf ? phv_data_241 : _GEN_754; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1013 = opcode == 4'hf ? phv_data_240 : _GEN_755; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1014 = opcode == 4'hf ? phv_data_247 : _GEN_756; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1015 = opcode == 4'hf ? phv_data_246 : _GEN_757; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1016 = opcode == 4'hf ? phv_data_245 : _GEN_758; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1017 = opcode == 4'hf ? phv_data_244 : _GEN_759; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1018 = opcode == 4'hf ? phv_data_251 : _GEN_760; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1019 = opcode == 4'hf ? phv_data_250 : _GEN_761; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1020 = opcode == 4'hf ? phv_data_249 : _GEN_762; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1021 = opcode == 4'hf ? phv_data_248 : _GEN_763; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1022 = opcode == 4'hf ? phv_data_255 : _GEN_764; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1023 = opcode == 4'hf ? phv_data_254 : _GEN_765; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1024 = opcode == 4'hf ? phv_data_253 : _GEN_766; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1025 = opcode == 4'hf ? phv_data_252 : _GEN_767; // @[executor.scala 466:52 executor.scala 450:25]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_1 = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8530 = {{2'd0}, dst_offset_1}; // @[executor.scala 473:49]
  wire [7:0] byte_256 = field_1[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1026 = mask_1[0] ? byte_256 : _GEN_770; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_257 = field_1[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1027 = mask_1[1] ? byte_257 : _GEN_771; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_258 = field_1[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1028 = mask_1[2] ? byte_258 : _GEN_772; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_259 = field_1[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1029 = mask_1[3] ? byte_259 : _GEN_773; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1030 = _GEN_8530 == 8'h0 ? _GEN_1026 : _GEN_770; // @[executor.scala 473:84]
  wire [7:0] _GEN_1031 = _GEN_8530 == 8'h0 ? _GEN_1027 : _GEN_771; // @[executor.scala 473:84]
  wire [7:0] _GEN_1032 = _GEN_8530 == 8'h0 ? _GEN_1028 : _GEN_772; // @[executor.scala 473:84]
  wire [7:0] _GEN_1033 = _GEN_8530 == 8'h0 ? _GEN_1029 : _GEN_773; // @[executor.scala 473:84]
  wire [7:0] _GEN_1034 = mask_1[0] ? byte_256 : _GEN_774; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1035 = mask_1[1] ? byte_257 : _GEN_775; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1036 = mask_1[2] ? byte_258 : _GEN_776; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1037 = mask_1[3] ? byte_259 : _GEN_777; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1038 = _GEN_8530 == 8'h1 ? _GEN_1034 : _GEN_774; // @[executor.scala 473:84]
  wire [7:0] _GEN_1039 = _GEN_8530 == 8'h1 ? _GEN_1035 : _GEN_775; // @[executor.scala 473:84]
  wire [7:0] _GEN_1040 = _GEN_8530 == 8'h1 ? _GEN_1036 : _GEN_776; // @[executor.scala 473:84]
  wire [7:0] _GEN_1041 = _GEN_8530 == 8'h1 ? _GEN_1037 : _GEN_777; // @[executor.scala 473:84]
  wire [7:0] _GEN_1042 = mask_1[0] ? byte_256 : _GEN_778; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1043 = mask_1[1] ? byte_257 : _GEN_779; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1044 = mask_1[2] ? byte_258 : _GEN_780; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1045 = mask_1[3] ? byte_259 : _GEN_781; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1046 = _GEN_8530 == 8'h2 ? _GEN_1042 : _GEN_778; // @[executor.scala 473:84]
  wire [7:0] _GEN_1047 = _GEN_8530 == 8'h2 ? _GEN_1043 : _GEN_779; // @[executor.scala 473:84]
  wire [7:0] _GEN_1048 = _GEN_8530 == 8'h2 ? _GEN_1044 : _GEN_780; // @[executor.scala 473:84]
  wire [7:0] _GEN_1049 = _GEN_8530 == 8'h2 ? _GEN_1045 : _GEN_781; // @[executor.scala 473:84]
  wire [7:0] _GEN_1050 = mask_1[0] ? byte_256 : _GEN_782; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1051 = mask_1[1] ? byte_257 : _GEN_783; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1052 = mask_1[2] ? byte_258 : _GEN_784; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1053 = mask_1[3] ? byte_259 : _GEN_785; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1054 = _GEN_8530 == 8'h3 ? _GEN_1050 : _GEN_782; // @[executor.scala 473:84]
  wire [7:0] _GEN_1055 = _GEN_8530 == 8'h3 ? _GEN_1051 : _GEN_783; // @[executor.scala 473:84]
  wire [7:0] _GEN_1056 = _GEN_8530 == 8'h3 ? _GEN_1052 : _GEN_784; // @[executor.scala 473:84]
  wire [7:0] _GEN_1057 = _GEN_8530 == 8'h3 ? _GEN_1053 : _GEN_785; // @[executor.scala 473:84]
  wire [7:0] _GEN_1058 = mask_1[0] ? byte_256 : _GEN_786; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1059 = mask_1[1] ? byte_257 : _GEN_787; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1060 = mask_1[2] ? byte_258 : _GEN_788; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1061 = mask_1[3] ? byte_259 : _GEN_789; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1062 = _GEN_8530 == 8'h4 ? _GEN_1058 : _GEN_786; // @[executor.scala 473:84]
  wire [7:0] _GEN_1063 = _GEN_8530 == 8'h4 ? _GEN_1059 : _GEN_787; // @[executor.scala 473:84]
  wire [7:0] _GEN_1064 = _GEN_8530 == 8'h4 ? _GEN_1060 : _GEN_788; // @[executor.scala 473:84]
  wire [7:0] _GEN_1065 = _GEN_8530 == 8'h4 ? _GEN_1061 : _GEN_789; // @[executor.scala 473:84]
  wire [7:0] _GEN_1066 = mask_1[0] ? byte_256 : _GEN_790; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1067 = mask_1[1] ? byte_257 : _GEN_791; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1068 = mask_1[2] ? byte_258 : _GEN_792; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1069 = mask_1[3] ? byte_259 : _GEN_793; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1070 = _GEN_8530 == 8'h5 ? _GEN_1066 : _GEN_790; // @[executor.scala 473:84]
  wire [7:0] _GEN_1071 = _GEN_8530 == 8'h5 ? _GEN_1067 : _GEN_791; // @[executor.scala 473:84]
  wire [7:0] _GEN_1072 = _GEN_8530 == 8'h5 ? _GEN_1068 : _GEN_792; // @[executor.scala 473:84]
  wire [7:0] _GEN_1073 = _GEN_8530 == 8'h5 ? _GEN_1069 : _GEN_793; // @[executor.scala 473:84]
  wire [7:0] _GEN_1074 = mask_1[0] ? byte_256 : _GEN_794; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1075 = mask_1[1] ? byte_257 : _GEN_795; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1076 = mask_1[2] ? byte_258 : _GEN_796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1077 = mask_1[3] ? byte_259 : _GEN_797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1078 = _GEN_8530 == 8'h6 ? _GEN_1074 : _GEN_794; // @[executor.scala 473:84]
  wire [7:0] _GEN_1079 = _GEN_8530 == 8'h6 ? _GEN_1075 : _GEN_795; // @[executor.scala 473:84]
  wire [7:0] _GEN_1080 = _GEN_8530 == 8'h6 ? _GEN_1076 : _GEN_796; // @[executor.scala 473:84]
  wire [7:0] _GEN_1081 = _GEN_8530 == 8'h6 ? _GEN_1077 : _GEN_797; // @[executor.scala 473:84]
  wire [7:0] _GEN_1082 = mask_1[0] ? byte_256 : _GEN_798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1083 = mask_1[1] ? byte_257 : _GEN_799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1084 = mask_1[2] ? byte_258 : _GEN_800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1085 = mask_1[3] ? byte_259 : _GEN_801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1086 = _GEN_8530 == 8'h7 ? _GEN_1082 : _GEN_798; // @[executor.scala 473:84]
  wire [7:0] _GEN_1087 = _GEN_8530 == 8'h7 ? _GEN_1083 : _GEN_799; // @[executor.scala 473:84]
  wire [7:0] _GEN_1088 = _GEN_8530 == 8'h7 ? _GEN_1084 : _GEN_800; // @[executor.scala 473:84]
  wire [7:0] _GEN_1089 = _GEN_8530 == 8'h7 ? _GEN_1085 : _GEN_801; // @[executor.scala 473:84]
  wire [7:0] _GEN_1090 = mask_1[0] ? byte_256 : _GEN_802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1091 = mask_1[1] ? byte_257 : _GEN_803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1092 = mask_1[2] ? byte_258 : _GEN_804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1093 = mask_1[3] ? byte_259 : _GEN_805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1094 = _GEN_8530 == 8'h8 ? _GEN_1090 : _GEN_802; // @[executor.scala 473:84]
  wire [7:0] _GEN_1095 = _GEN_8530 == 8'h8 ? _GEN_1091 : _GEN_803; // @[executor.scala 473:84]
  wire [7:0] _GEN_1096 = _GEN_8530 == 8'h8 ? _GEN_1092 : _GEN_804; // @[executor.scala 473:84]
  wire [7:0] _GEN_1097 = _GEN_8530 == 8'h8 ? _GEN_1093 : _GEN_805; // @[executor.scala 473:84]
  wire [7:0] _GEN_1098 = mask_1[0] ? byte_256 : _GEN_806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1099 = mask_1[1] ? byte_257 : _GEN_807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1100 = mask_1[2] ? byte_258 : _GEN_808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1101 = mask_1[3] ? byte_259 : _GEN_809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1102 = _GEN_8530 == 8'h9 ? _GEN_1098 : _GEN_806; // @[executor.scala 473:84]
  wire [7:0] _GEN_1103 = _GEN_8530 == 8'h9 ? _GEN_1099 : _GEN_807; // @[executor.scala 473:84]
  wire [7:0] _GEN_1104 = _GEN_8530 == 8'h9 ? _GEN_1100 : _GEN_808; // @[executor.scala 473:84]
  wire [7:0] _GEN_1105 = _GEN_8530 == 8'h9 ? _GEN_1101 : _GEN_809; // @[executor.scala 473:84]
  wire [7:0] _GEN_1106 = mask_1[0] ? byte_256 : _GEN_810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1107 = mask_1[1] ? byte_257 : _GEN_811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1108 = mask_1[2] ? byte_258 : _GEN_812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1109 = mask_1[3] ? byte_259 : _GEN_813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1110 = _GEN_8530 == 8'ha ? _GEN_1106 : _GEN_810; // @[executor.scala 473:84]
  wire [7:0] _GEN_1111 = _GEN_8530 == 8'ha ? _GEN_1107 : _GEN_811; // @[executor.scala 473:84]
  wire [7:0] _GEN_1112 = _GEN_8530 == 8'ha ? _GEN_1108 : _GEN_812; // @[executor.scala 473:84]
  wire [7:0] _GEN_1113 = _GEN_8530 == 8'ha ? _GEN_1109 : _GEN_813; // @[executor.scala 473:84]
  wire [7:0] _GEN_1114 = mask_1[0] ? byte_256 : _GEN_814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1115 = mask_1[1] ? byte_257 : _GEN_815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1116 = mask_1[2] ? byte_258 : _GEN_816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1117 = mask_1[3] ? byte_259 : _GEN_817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1118 = _GEN_8530 == 8'hb ? _GEN_1114 : _GEN_814; // @[executor.scala 473:84]
  wire [7:0] _GEN_1119 = _GEN_8530 == 8'hb ? _GEN_1115 : _GEN_815; // @[executor.scala 473:84]
  wire [7:0] _GEN_1120 = _GEN_8530 == 8'hb ? _GEN_1116 : _GEN_816; // @[executor.scala 473:84]
  wire [7:0] _GEN_1121 = _GEN_8530 == 8'hb ? _GEN_1117 : _GEN_817; // @[executor.scala 473:84]
  wire [7:0] _GEN_1122 = mask_1[0] ? byte_256 : _GEN_818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1123 = mask_1[1] ? byte_257 : _GEN_819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1124 = mask_1[2] ? byte_258 : _GEN_820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1125 = mask_1[3] ? byte_259 : _GEN_821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1126 = _GEN_8530 == 8'hc ? _GEN_1122 : _GEN_818; // @[executor.scala 473:84]
  wire [7:0] _GEN_1127 = _GEN_8530 == 8'hc ? _GEN_1123 : _GEN_819; // @[executor.scala 473:84]
  wire [7:0] _GEN_1128 = _GEN_8530 == 8'hc ? _GEN_1124 : _GEN_820; // @[executor.scala 473:84]
  wire [7:0] _GEN_1129 = _GEN_8530 == 8'hc ? _GEN_1125 : _GEN_821; // @[executor.scala 473:84]
  wire [7:0] _GEN_1130 = mask_1[0] ? byte_256 : _GEN_822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1131 = mask_1[1] ? byte_257 : _GEN_823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1132 = mask_1[2] ? byte_258 : _GEN_824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1133 = mask_1[3] ? byte_259 : _GEN_825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1134 = _GEN_8530 == 8'hd ? _GEN_1130 : _GEN_822; // @[executor.scala 473:84]
  wire [7:0] _GEN_1135 = _GEN_8530 == 8'hd ? _GEN_1131 : _GEN_823; // @[executor.scala 473:84]
  wire [7:0] _GEN_1136 = _GEN_8530 == 8'hd ? _GEN_1132 : _GEN_824; // @[executor.scala 473:84]
  wire [7:0] _GEN_1137 = _GEN_8530 == 8'hd ? _GEN_1133 : _GEN_825; // @[executor.scala 473:84]
  wire [7:0] _GEN_1138 = mask_1[0] ? byte_256 : _GEN_826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1139 = mask_1[1] ? byte_257 : _GEN_827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1140 = mask_1[2] ? byte_258 : _GEN_828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1141 = mask_1[3] ? byte_259 : _GEN_829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1142 = _GEN_8530 == 8'he ? _GEN_1138 : _GEN_826; // @[executor.scala 473:84]
  wire [7:0] _GEN_1143 = _GEN_8530 == 8'he ? _GEN_1139 : _GEN_827; // @[executor.scala 473:84]
  wire [7:0] _GEN_1144 = _GEN_8530 == 8'he ? _GEN_1140 : _GEN_828; // @[executor.scala 473:84]
  wire [7:0] _GEN_1145 = _GEN_8530 == 8'he ? _GEN_1141 : _GEN_829; // @[executor.scala 473:84]
  wire [7:0] _GEN_1146 = mask_1[0] ? byte_256 : _GEN_830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1147 = mask_1[1] ? byte_257 : _GEN_831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1148 = mask_1[2] ? byte_258 : _GEN_832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1149 = mask_1[3] ? byte_259 : _GEN_833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1150 = _GEN_8530 == 8'hf ? _GEN_1146 : _GEN_830; // @[executor.scala 473:84]
  wire [7:0] _GEN_1151 = _GEN_8530 == 8'hf ? _GEN_1147 : _GEN_831; // @[executor.scala 473:84]
  wire [7:0] _GEN_1152 = _GEN_8530 == 8'hf ? _GEN_1148 : _GEN_832; // @[executor.scala 473:84]
  wire [7:0] _GEN_1153 = _GEN_8530 == 8'hf ? _GEN_1149 : _GEN_833; // @[executor.scala 473:84]
  wire [7:0] _GEN_1154 = mask_1[0] ? byte_256 : _GEN_834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1155 = mask_1[1] ? byte_257 : _GEN_835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1156 = mask_1[2] ? byte_258 : _GEN_836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1157 = mask_1[3] ? byte_259 : _GEN_837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1158 = _GEN_8530 == 8'h10 ? _GEN_1154 : _GEN_834; // @[executor.scala 473:84]
  wire [7:0] _GEN_1159 = _GEN_8530 == 8'h10 ? _GEN_1155 : _GEN_835; // @[executor.scala 473:84]
  wire [7:0] _GEN_1160 = _GEN_8530 == 8'h10 ? _GEN_1156 : _GEN_836; // @[executor.scala 473:84]
  wire [7:0] _GEN_1161 = _GEN_8530 == 8'h10 ? _GEN_1157 : _GEN_837; // @[executor.scala 473:84]
  wire [7:0] _GEN_1162 = mask_1[0] ? byte_256 : _GEN_838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1163 = mask_1[1] ? byte_257 : _GEN_839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1164 = mask_1[2] ? byte_258 : _GEN_840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1165 = mask_1[3] ? byte_259 : _GEN_841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1166 = _GEN_8530 == 8'h11 ? _GEN_1162 : _GEN_838; // @[executor.scala 473:84]
  wire [7:0] _GEN_1167 = _GEN_8530 == 8'h11 ? _GEN_1163 : _GEN_839; // @[executor.scala 473:84]
  wire [7:0] _GEN_1168 = _GEN_8530 == 8'h11 ? _GEN_1164 : _GEN_840; // @[executor.scala 473:84]
  wire [7:0] _GEN_1169 = _GEN_8530 == 8'h11 ? _GEN_1165 : _GEN_841; // @[executor.scala 473:84]
  wire [7:0] _GEN_1170 = mask_1[0] ? byte_256 : _GEN_842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1171 = mask_1[1] ? byte_257 : _GEN_843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1172 = mask_1[2] ? byte_258 : _GEN_844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1173 = mask_1[3] ? byte_259 : _GEN_845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1174 = _GEN_8530 == 8'h12 ? _GEN_1170 : _GEN_842; // @[executor.scala 473:84]
  wire [7:0] _GEN_1175 = _GEN_8530 == 8'h12 ? _GEN_1171 : _GEN_843; // @[executor.scala 473:84]
  wire [7:0] _GEN_1176 = _GEN_8530 == 8'h12 ? _GEN_1172 : _GEN_844; // @[executor.scala 473:84]
  wire [7:0] _GEN_1177 = _GEN_8530 == 8'h12 ? _GEN_1173 : _GEN_845; // @[executor.scala 473:84]
  wire [7:0] _GEN_1178 = mask_1[0] ? byte_256 : _GEN_846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1179 = mask_1[1] ? byte_257 : _GEN_847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1180 = mask_1[2] ? byte_258 : _GEN_848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1181 = mask_1[3] ? byte_259 : _GEN_849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1182 = _GEN_8530 == 8'h13 ? _GEN_1178 : _GEN_846; // @[executor.scala 473:84]
  wire [7:0] _GEN_1183 = _GEN_8530 == 8'h13 ? _GEN_1179 : _GEN_847; // @[executor.scala 473:84]
  wire [7:0] _GEN_1184 = _GEN_8530 == 8'h13 ? _GEN_1180 : _GEN_848; // @[executor.scala 473:84]
  wire [7:0] _GEN_1185 = _GEN_8530 == 8'h13 ? _GEN_1181 : _GEN_849; // @[executor.scala 473:84]
  wire [7:0] _GEN_1186 = mask_1[0] ? byte_256 : _GEN_850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1187 = mask_1[1] ? byte_257 : _GEN_851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1188 = mask_1[2] ? byte_258 : _GEN_852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1189 = mask_1[3] ? byte_259 : _GEN_853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1190 = _GEN_8530 == 8'h14 ? _GEN_1186 : _GEN_850; // @[executor.scala 473:84]
  wire [7:0] _GEN_1191 = _GEN_8530 == 8'h14 ? _GEN_1187 : _GEN_851; // @[executor.scala 473:84]
  wire [7:0] _GEN_1192 = _GEN_8530 == 8'h14 ? _GEN_1188 : _GEN_852; // @[executor.scala 473:84]
  wire [7:0] _GEN_1193 = _GEN_8530 == 8'h14 ? _GEN_1189 : _GEN_853; // @[executor.scala 473:84]
  wire [7:0] _GEN_1194 = mask_1[0] ? byte_256 : _GEN_854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1195 = mask_1[1] ? byte_257 : _GEN_855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1196 = mask_1[2] ? byte_258 : _GEN_856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1197 = mask_1[3] ? byte_259 : _GEN_857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1198 = _GEN_8530 == 8'h15 ? _GEN_1194 : _GEN_854; // @[executor.scala 473:84]
  wire [7:0] _GEN_1199 = _GEN_8530 == 8'h15 ? _GEN_1195 : _GEN_855; // @[executor.scala 473:84]
  wire [7:0] _GEN_1200 = _GEN_8530 == 8'h15 ? _GEN_1196 : _GEN_856; // @[executor.scala 473:84]
  wire [7:0] _GEN_1201 = _GEN_8530 == 8'h15 ? _GEN_1197 : _GEN_857; // @[executor.scala 473:84]
  wire [7:0] _GEN_1202 = mask_1[0] ? byte_256 : _GEN_858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1203 = mask_1[1] ? byte_257 : _GEN_859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1204 = mask_1[2] ? byte_258 : _GEN_860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1205 = mask_1[3] ? byte_259 : _GEN_861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1206 = _GEN_8530 == 8'h16 ? _GEN_1202 : _GEN_858; // @[executor.scala 473:84]
  wire [7:0] _GEN_1207 = _GEN_8530 == 8'h16 ? _GEN_1203 : _GEN_859; // @[executor.scala 473:84]
  wire [7:0] _GEN_1208 = _GEN_8530 == 8'h16 ? _GEN_1204 : _GEN_860; // @[executor.scala 473:84]
  wire [7:0] _GEN_1209 = _GEN_8530 == 8'h16 ? _GEN_1205 : _GEN_861; // @[executor.scala 473:84]
  wire [7:0] _GEN_1210 = mask_1[0] ? byte_256 : _GEN_862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1211 = mask_1[1] ? byte_257 : _GEN_863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1212 = mask_1[2] ? byte_258 : _GEN_864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1213 = mask_1[3] ? byte_259 : _GEN_865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1214 = _GEN_8530 == 8'h17 ? _GEN_1210 : _GEN_862; // @[executor.scala 473:84]
  wire [7:0] _GEN_1215 = _GEN_8530 == 8'h17 ? _GEN_1211 : _GEN_863; // @[executor.scala 473:84]
  wire [7:0] _GEN_1216 = _GEN_8530 == 8'h17 ? _GEN_1212 : _GEN_864; // @[executor.scala 473:84]
  wire [7:0] _GEN_1217 = _GEN_8530 == 8'h17 ? _GEN_1213 : _GEN_865; // @[executor.scala 473:84]
  wire [7:0] _GEN_1218 = mask_1[0] ? byte_256 : _GEN_866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1219 = mask_1[1] ? byte_257 : _GEN_867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1220 = mask_1[2] ? byte_258 : _GEN_868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1221 = mask_1[3] ? byte_259 : _GEN_869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1222 = _GEN_8530 == 8'h18 ? _GEN_1218 : _GEN_866; // @[executor.scala 473:84]
  wire [7:0] _GEN_1223 = _GEN_8530 == 8'h18 ? _GEN_1219 : _GEN_867; // @[executor.scala 473:84]
  wire [7:0] _GEN_1224 = _GEN_8530 == 8'h18 ? _GEN_1220 : _GEN_868; // @[executor.scala 473:84]
  wire [7:0] _GEN_1225 = _GEN_8530 == 8'h18 ? _GEN_1221 : _GEN_869; // @[executor.scala 473:84]
  wire [7:0] _GEN_1226 = mask_1[0] ? byte_256 : _GEN_870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1227 = mask_1[1] ? byte_257 : _GEN_871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1228 = mask_1[2] ? byte_258 : _GEN_872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1229 = mask_1[3] ? byte_259 : _GEN_873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1230 = _GEN_8530 == 8'h19 ? _GEN_1226 : _GEN_870; // @[executor.scala 473:84]
  wire [7:0] _GEN_1231 = _GEN_8530 == 8'h19 ? _GEN_1227 : _GEN_871; // @[executor.scala 473:84]
  wire [7:0] _GEN_1232 = _GEN_8530 == 8'h19 ? _GEN_1228 : _GEN_872; // @[executor.scala 473:84]
  wire [7:0] _GEN_1233 = _GEN_8530 == 8'h19 ? _GEN_1229 : _GEN_873; // @[executor.scala 473:84]
  wire [7:0] _GEN_1234 = mask_1[0] ? byte_256 : _GEN_874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1235 = mask_1[1] ? byte_257 : _GEN_875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1236 = mask_1[2] ? byte_258 : _GEN_876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1237 = mask_1[3] ? byte_259 : _GEN_877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1238 = _GEN_8530 == 8'h1a ? _GEN_1234 : _GEN_874; // @[executor.scala 473:84]
  wire [7:0] _GEN_1239 = _GEN_8530 == 8'h1a ? _GEN_1235 : _GEN_875; // @[executor.scala 473:84]
  wire [7:0] _GEN_1240 = _GEN_8530 == 8'h1a ? _GEN_1236 : _GEN_876; // @[executor.scala 473:84]
  wire [7:0] _GEN_1241 = _GEN_8530 == 8'h1a ? _GEN_1237 : _GEN_877; // @[executor.scala 473:84]
  wire [7:0] _GEN_1242 = mask_1[0] ? byte_256 : _GEN_878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1243 = mask_1[1] ? byte_257 : _GEN_879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1244 = mask_1[2] ? byte_258 : _GEN_880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1245 = mask_1[3] ? byte_259 : _GEN_881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1246 = _GEN_8530 == 8'h1b ? _GEN_1242 : _GEN_878; // @[executor.scala 473:84]
  wire [7:0] _GEN_1247 = _GEN_8530 == 8'h1b ? _GEN_1243 : _GEN_879; // @[executor.scala 473:84]
  wire [7:0] _GEN_1248 = _GEN_8530 == 8'h1b ? _GEN_1244 : _GEN_880; // @[executor.scala 473:84]
  wire [7:0] _GEN_1249 = _GEN_8530 == 8'h1b ? _GEN_1245 : _GEN_881; // @[executor.scala 473:84]
  wire [7:0] _GEN_1250 = mask_1[0] ? byte_256 : _GEN_882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1251 = mask_1[1] ? byte_257 : _GEN_883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1252 = mask_1[2] ? byte_258 : _GEN_884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1253 = mask_1[3] ? byte_259 : _GEN_885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1254 = _GEN_8530 == 8'h1c ? _GEN_1250 : _GEN_882; // @[executor.scala 473:84]
  wire [7:0] _GEN_1255 = _GEN_8530 == 8'h1c ? _GEN_1251 : _GEN_883; // @[executor.scala 473:84]
  wire [7:0] _GEN_1256 = _GEN_8530 == 8'h1c ? _GEN_1252 : _GEN_884; // @[executor.scala 473:84]
  wire [7:0] _GEN_1257 = _GEN_8530 == 8'h1c ? _GEN_1253 : _GEN_885; // @[executor.scala 473:84]
  wire [7:0] _GEN_1258 = mask_1[0] ? byte_256 : _GEN_886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1259 = mask_1[1] ? byte_257 : _GEN_887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1260 = mask_1[2] ? byte_258 : _GEN_888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1261 = mask_1[3] ? byte_259 : _GEN_889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1262 = _GEN_8530 == 8'h1d ? _GEN_1258 : _GEN_886; // @[executor.scala 473:84]
  wire [7:0] _GEN_1263 = _GEN_8530 == 8'h1d ? _GEN_1259 : _GEN_887; // @[executor.scala 473:84]
  wire [7:0] _GEN_1264 = _GEN_8530 == 8'h1d ? _GEN_1260 : _GEN_888; // @[executor.scala 473:84]
  wire [7:0] _GEN_1265 = _GEN_8530 == 8'h1d ? _GEN_1261 : _GEN_889; // @[executor.scala 473:84]
  wire [7:0] _GEN_1266 = mask_1[0] ? byte_256 : _GEN_890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1267 = mask_1[1] ? byte_257 : _GEN_891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1268 = mask_1[2] ? byte_258 : _GEN_892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1269 = mask_1[3] ? byte_259 : _GEN_893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1270 = _GEN_8530 == 8'h1e ? _GEN_1266 : _GEN_890; // @[executor.scala 473:84]
  wire [7:0] _GEN_1271 = _GEN_8530 == 8'h1e ? _GEN_1267 : _GEN_891; // @[executor.scala 473:84]
  wire [7:0] _GEN_1272 = _GEN_8530 == 8'h1e ? _GEN_1268 : _GEN_892; // @[executor.scala 473:84]
  wire [7:0] _GEN_1273 = _GEN_8530 == 8'h1e ? _GEN_1269 : _GEN_893; // @[executor.scala 473:84]
  wire [7:0] _GEN_1274 = mask_1[0] ? byte_256 : _GEN_894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1275 = mask_1[1] ? byte_257 : _GEN_895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1276 = mask_1[2] ? byte_258 : _GEN_896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1277 = mask_1[3] ? byte_259 : _GEN_897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1278 = _GEN_8530 == 8'h1f ? _GEN_1274 : _GEN_894; // @[executor.scala 473:84]
  wire [7:0] _GEN_1279 = _GEN_8530 == 8'h1f ? _GEN_1275 : _GEN_895; // @[executor.scala 473:84]
  wire [7:0] _GEN_1280 = _GEN_8530 == 8'h1f ? _GEN_1276 : _GEN_896; // @[executor.scala 473:84]
  wire [7:0] _GEN_1281 = _GEN_8530 == 8'h1f ? _GEN_1277 : _GEN_897; // @[executor.scala 473:84]
  wire [7:0] _GEN_1282 = mask_1[0] ? byte_256 : _GEN_898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1283 = mask_1[1] ? byte_257 : _GEN_899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1284 = mask_1[2] ? byte_258 : _GEN_900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1285 = mask_1[3] ? byte_259 : _GEN_901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1286 = _GEN_8530 == 8'h20 ? _GEN_1282 : _GEN_898; // @[executor.scala 473:84]
  wire [7:0] _GEN_1287 = _GEN_8530 == 8'h20 ? _GEN_1283 : _GEN_899; // @[executor.scala 473:84]
  wire [7:0] _GEN_1288 = _GEN_8530 == 8'h20 ? _GEN_1284 : _GEN_900; // @[executor.scala 473:84]
  wire [7:0] _GEN_1289 = _GEN_8530 == 8'h20 ? _GEN_1285 : _GEN_901; // @[executor.scala 473:84]
  wire [7:0] _GEN_1290 = mask_1[0] ? byte_256 : _GEN_902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1291 = mask_1[1] ? byte_257 : _GEN_903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1292 = mask_1[2] ? byte_258 : _GEN_904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1293 = mask_1[3] ? byte_259 : _GEN_905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1294 = _GEN_8530 == 8'h21 ? _GEN_1290 : _GEN_902; // @[executor.scala 473:84]
  wire [7:0] _GEN_1295 = _GEN_8530 == 8'h21 ? _GEN_1291 : _GEN_903; // @[executor.scala 473:84]
  wire [7:0] _GEN_1296 = _GEN_8530 == 8'h21 ? _GEN_1292 : _GEN_904; // @[executor.scala 473:84]
  wire [7:0] _GEN_1297 = _GEN_8530 == 8'h21 ? _GEN_1293 : _GEN_905; // @[executor.scala 473:84]
  wire [7:0] _GEN_1298 = mask_1[0] ? byte_256 : _GEN_906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1299 = mask_1[1] ? byte_257 : _GEN_907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1300 = mask_1[2] ? byte_258 : _GEN_908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1301 = mask_1[3] ? byte_259 : _GEN_909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1302 = _GEN_8530 == 8'h22 ? _GEN_1298 : _GEN_906; // @[executor.scala 473:84]
  wire [7:0] _GEN_1303 = _GEN_8530 == 8'h22 ? _GEN_1299 : _GEN_907; // @[executor.scala 473:84]
  wire [7:0] _GEN_1304 = _GEN_8530 == 8'h22 ? _GEN_1300 : _GEN_908; // @[executor.scala 473:84]
  wire [7:0] _GEN_1305 = _GEN_8530 == 8'h22 ? _GEN_1301 : _GEN_909; // @[executor.scala 473:84]
  wire [7:0] _GEN_1306 = mask_1[0] ? byte_256 : _GEN_910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1307 = mask_1[1] ? byte_257 : _GEN_911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1308 = mask_1[2] ? byte_258 : _GEN_912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1309 = mask_1[3] ? byte_259 : _GEN_913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1310 = _GEN_8530 == 8'h23 ? _GEN_1306 : _GEN_910; // @[executor.scala 473:84]
  wire [7:0] _GEN_1311 = _GEN_8530 == 8'h23 ? _GEN_1307 : _GEN_911; // @[executor.scala 473:84]
  wire [7:0] _GEN_1312 = _GEN_8530 == 8'h23 ? _GEN_1308 : _GEN_912; // @[executor.scala 473:84]
  wire [7:0] _GEN_1313 = _GEN_8530 == 8'h23 ? _GEN_1309 : _GEN_913; // @[executor.scala 473:84]
  wire [7:0] _GEN_1314 = mask_1[0] ? byte_256 : _GEN_914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1315 = mask_1[1] ? byte_257 : _GEN_915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1316 = mask_1[2] ? byte_258 : _GEN_916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1317 = mask_1[3] ? byte_259 : _GEN_917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1318 = _GEN_8530 == 8'h24 ? _GEN_1314 : _GEN_914; // @[executor.scala 473:84]
  wire [7:0] _GEN_1319 = _GEN_8530 == 8'h24 ? _GEN_1315 : _GEN_915; // @[executor.scala 473:84]
  wire [7:0] _GEN_1320 = _GEN_8530 == 8'h24 ? _GEN_1316 : _GEN_916; // @[executor.scala 473:84]
  wire [7:0] _GEN_1321 = _GEN_8530 == 8'h24 ? _GEN_1317 : _GEN_917; // @[executor.scala 473:84]
  wire [7:0] _GEN_1322 = mask_1[0] ? byte_256 : _GEN_918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1323 = mask_1[1] ? byte_257 : _GEN_919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1324 = mask_1[2] ? byte_258 : _GEN_920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1325 = mask_1[3] ? byte_259 : _GEN_921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1326 = _GEN_8530 == 8'h25 ? _GEN_1322 : _GEN_918; // @[executor.scala 473:84]
  wire [7:0] _GEN_1327 = _GEN_8530 == 8'h25 ? _GEN_1323 : _GEN_919; // @[executor.scala 473:84]
  wire [7:0] _GEN_1328 = _GEN_8530 == 8'h25 ? _GEN_1324 : _GEN_920; // @[executor.scala 473:84]
  wire [7:0] _GEN_1329 = _GEN_8530 == 8'h25 ? _GEN_1325 : _GEN_921; // @[executor.scala 473:84]
  wire [7:0] _GEN_1330 = mask_1[0] ? byte_256 : _GEN_922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1331 = mask_1[1] ? byte_257 : _GEN_923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1332 = mask_1[2] ? byte_258 : _GEN_924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1333 = mask_1[3] ? byte_259 : _GEN_925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1334 = _GEN_8530 == 8'h26 ? _GEN_1330 : _GEN_922; // @[executor.scala 473:84]
  wire [7:0] _GEN_1335 = _GEN_8530 == 8'h26 ? _GEN_1331 : _GEN_923; // @[executor.scala 473:84]
  wire [7:0] _GEN_1336 = _GEN_8530 == 8'h26 ? _GEN_1332 : _GEN_924; // @[executor.scala 473:84]
  wire [7:0] _GEN_1337 = _GEN_8530 == 8'h26 ? _GEN_1333 : _GEN_925; // @[executor.scala 473:84]
  wire [7:0] _GEN_1338 = mask_1[0] ? byte_256 : _GEN_926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1339 = mask_1[1] ? byte_257 : _GEN_927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1340 = mask_1[2] ? byte_258 : _GEN_928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1341 = mask_1[3] ? byte_259 : _GEN_929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1342 = _GEN_8530 == 8'h27 ? _GEN_1338 : _GEN_926; // @[executor.scala 473:84]
  wire [7:0] _GEN_1343 = _GEN_8530 == 8'h27 ? _GEN_1339 : _GEN_927; // @[executor.scala 473:84]
  wire [7:0] _GEN_1344 = _GEN_8530 == 8'h27 ? _GEN_1340 : _GEN_928; // @[executor.scala 473:84]
  wire [7:0] _GEN_1345 = _GEN_8530 == 8'h27 ? _GEN_1341 : _GEN_929; // @[executor.scala 473:84]
  wire [7:0] _GEN_1346 = mask_1[0] ? byte_256 : _GEN_930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1347 = mask_1[1] ? byte_257 : _GEN_931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1348 = mask_1[2] ? byte_258 : _GEN_932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1349 = mask_1[3] ? byte_259 : _GEN_933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1350 = _GEN_8530 == 8'h28 ? _GEN_1346 : _GEN_930; // @[executor.scala 473:84]
  wire [7:0] _GEN_1351 = _GEN_8530 == 8'h28 ? _GEN_1347 : _GEN_931; // @[executor.scala 473:84]
  wire [7:0] _GEN_1352 = _GEN_8530 == 8'h28 ? _GEN_1348 : _GEN_932; // @[executor.scala 473:84]
  wire [7:0] _GEN_1353 = _GEN_8530 == 8'h28 ? _GEN_1349 : _GEN_933; // @[executor.scala 473:84]
  wire [7:0] _GEN_1354 = mask_1[0] ? byte_256 : _GEN_934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1355 = mask_1[1] ? byte_257 : _GEN_935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1356 = mask_1[2] ? byte_258 : _GEN_936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1357 = mask_1[3] ? byte_259 : _GEN_937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1358 = _GEN_8530 == 8'h29 ? _GEN_1354 : _GEN_934; // @[executor.scala 473:84]
  wire [7:0] _GEN_1359 = _GEN_8530 == 8'h29 ? _GEN_1355 : _GEN_935; // @[executor.scala 473:84]
  wire [7:0] _GEN_1360 = _GEN_8530 == 8'h29 ? _GEN_1356 : _GEN_936; // @[executor.scala 473:84]
  wire [7:0] _GEN_1361 = _GEN_8530 == 8'h29 ? _GEN_1357 : _GEN_937; // @[executor.scala 473:84]
  wire [7:0] _GEN_1362 = mask_1[0] ? byte_256 : _GEN_938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1363 = mask_1[1] ? byte_257 : _GEN_939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1364 = mask_1[2] ? byte_258 : _GEN_940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1365 = mask_1[3] ? byte_259 : _GEN_941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1366 = _GEN_8530 == 8'h2a ? _GEN_1362 : _GEN_938; // @[executor.scala 473:84]
  wire [7:0] _GEN_1367 = _GEN_8530 == 8'h2a ? _GEN_1363 : _GEN_939; // @[executor.scala 473:84]
  wire [7:0] _GEN_1368 = _GEN_8530 == 8'h2a ? _GEN_1364 : _GEN_940; // @[executor.scala 473:84]
  wire [7:0] _GEN_1369 = _GEN_8530 == 8'h2a ? _GEN_1365 : _GEN_941; // @[executor.scala 473:84]
  wire [7:0] _GEN_1370 = mask_1[0] ? byte_256 : _GEN_942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1371 = mask_1[1] ? byte_257 : _GEN_943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1372 = mask_1[2] ? byte_258 : _GEN_944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1373 = mask_1[3] ? byte_259 : _GEN_945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1374 = _GEN_8530 == 8'h2b ? _GEN_1370 : _GEN_942; // @[executor.scala 473:84]
  wire [7:0] _GEN_1375 = _GEN_8530 == 8'h2b ? _GEN_1371 : _GEN_943; // @[executor.scala 473:84]
  wire [7:0] _GEN_1376 = _GEN_8530 == 8'h2b ? _GEN_1372 : _GEN_944; // @[executor.scala 473:84]
  wire [7:0] _GEN_1377 = _GEN_8530 == 8'h2b ? _GEN_1373 : _GEN_945; // @[executor.scala 473:84]
  wire [7:0] _GEN_1378 = mask_1[0] ? byte_256 : _GEN_946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1379 = mask_1[1] ? byte_257 : _GEN_947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1380 = mask_1[2] ? byte_258 : _GEN_948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1381 = mask_1[3] ? byte_259 : _GEN_949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1382 = _GEN_8530 == 8'h2c ? _GEN_1378 : _GEN_946; // @[executor.scala 473:84]
  wire [7:0] _GEN_1383 = _GEN_8530 == 8'h2c ? _GEN_1379 : _GEN_947; // @[executor.scala 473:84]
  wire [7:0] _GEN_1384 = _GEN_8530 == 8'h2c ? _GEN_1380 : _GEN_948; // @[executor.scala 473:84]
  wire [7:0] _GEN_1385 = _GEN_8530 == 8'h2c ? _GEN_1381 : _GEN_949; // @[executor.scala 473:84]
  wire [7:0] _GEN_1386 = mask_1[0] ? byte_256 : _GEN_950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1387 = mask_1[1] ? byte_257 : _GEN_951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1388 = mask_1[2] ? byte_258 : _GEN_952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1389 = mask_1[3] ? byte_259 : _GEN_953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1390 = _GEN_8530 == 8'h2d ? _GEN_1386 : _GEN_950; // @[executor.scala 473:84]
  wire [7:0] _GEN_1391 = _GEN_8530 == 8'h2d ? _GEN_1387 : _GEN_951; // @[executor.scala 473:84]
  wire [7:0] _GEN_1392 = _GEN_8530 == 8'h2d ? _GEN_1388 : _GEN_952; // @[executor.scala 473:84]
  wire [7:0] _GEN_1393 = _GEN_8530 == 8'h2d ? _GEN_1389 : _GEN_953; // @[executor.scala 473:84]
  wire [7:0] _GEN_1394 = mask_1[0] ? byte_256 : _GEN_954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1395 = mask_1[1] ? byte_257 : _GEN_955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1396 = mask_1[2] ? byte_258 : _GEN_956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1397 = mask_1[3] ? byte_259 : _GEN_957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1398 = _GEN_8530 == 8'h2e ? _GEN_1394 : _GEN_954; // @[executor.scala 473:84]
  wire [7:0] _GEN_1399 = _GEN_8530 == 8'h2e ? _GEN_1395 : _GEN_955; // @[executor.scala 473:84]
  wire [7:0] _GEN_1400 = _GEN_8530 == 8'h2e ? _GEN_1396 : _GEN_956; // @[executor.scala 473:84]
  wire [7:0] _GEN_1401 = _GEN_8530 == 8'h2e ? _GEN_1397 : _GEN_957; // @[executor.scala 473:84]
  wire [7:0] _GEN_1402 = mask_1[0] ? byte_256 : _GEN_958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1403 = mask_1[1] ? byte_257 : _GEN_959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1404 = mask_1[2] ? byte_258 : _GEN_960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1405 = mask_1[3] ? byte_259 : _GEN_961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1406 = _GEN_8530 == 8'h2f ? _GEN_1402 : _GEN_958; // @[executor.scala 473:84]
  wire [7:0] _GEN_1407 = _GEN_8530 == 8'h2f ? _GEN_1403 : _GEN_959; // @[executor.scala 473:84]
  wire [7:0] _GEN_1408 = _GEN_8530 == 8'h2f ? _GEN_1404 : _GEN_960; // @[executor.scala 473:84]
  wire [7:0] _GEN_1409 = _GEN_8530 == 8'h2f ? _GEN_1405 : _GEN_961; // @[executor.scala 473:84]
  wire [7:0] _GEN_1410 = mask_1[0] ? byte_256 : _GEN_962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1411 = mask_1[1] ? byte_257 : _GEN_963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1412 = mask_1[2] ? byte_258 : _GEN_964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1413 = mask_1[3] ? byte_259 : _GEN_965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1414 = _GEN_8530 == 8'h30 ? _GEN_1410 : _GEN_962; // @[executor.scala 473:84]
  wire [7:0] _GEN_1415 = _GEN_8530 == 8'h30 ? _GEN_1411 : _GEN_963; // @[executor.scala 473:84]
  wire [7:0] _GEN_1416 = _GEN_8530 == 8'h30 ? _GEN_1412 : _GEN_964; // @[executor.scala 473:84]
  wire [7:0] _GEN_1417 = _GEN_8530 == 8'h30 ? _GEN_1413 : _GEN_965; // @[executor.scala 473:84]
  wire [7:0] _GEN_1418 = mask_1[0] ? byte_256 : _GEN_966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1419 = mask_1[1] ? byte_257 : _GEN_967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1420 = mask_1[2] ? byte_258 : _GEN_968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1421 = mask_1[3] ? byte_259 : _GEN_969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1422 = _GEN_8530 == 8'h31 ? _GEN_1418 : _GEN_966; // @[executor.scala 473:84]
  wire [7:0] _GEN_1423 = _GEN_8530 == 8'h31 ? _GEN_1419 : _GEN_967; // @[executor.scala 473:84]
  wire [7:0] _GEN_1424 = _GEN_8530 == 8'h31 ? _GEN_1420 : _GEN_968; // @[executor.scala 473:84]
  wire [7:0] _GEN_1425 = _GEN_8530 == 8'h31 ? _GEN_1421 : _GEN_969; // @[executor.scala 473:84]
  wire [7:0] _GEN_1426 = mask_1[0] ? byte_256 : _GEN_970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1427 = mask_1[1] ? byte_257 : _GEN_971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1428 = mask_1[2] ? byte_258 : _GEN_972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1429 = mask_1[3] ? byte_259 : _GEN_973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1430 = _GEN_8530 == 8'h32 ? _GEN_1426 : _GEN_970; // @[executor.scala 473:84]
  wire [7:0] _GEN_1431 = _GEN_8530 == 8'h32 ? _GEN_1427 : _GEN_971; // @[executor.scala 473:84]
  wire [7:0] _GEN_1432 = _GEN_8530 == 8'h32 ? _GEN_1428 : _GEN_972; // @[executor.scala 473:84]
  wire [7:0] _GEN_1433 = _GEN_8530 == 8'h32 ? _GEN_1429 : _GEN_973; // @[executor.scala 473:84]
  wire [7:0] _GEN_1434 = mask_1[0] ? byte_256 : _GEN_974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1435 = mask_1[1] ? byte_257 : _GEN_975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1436 = mask_1[2] ? byte_258 : _GEN_976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1437 = mask_1[3] ? byte_259 : _GEN_977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1438 = _GEN_8530 == 8'h33 ? _GEN_1434 : _GEN_974; // @[executor.scala 473:84]
  wire [7:0] _GEN_1439 = _GEN_8530 == 8'h33 ? _GEN_1435 : _GEN_975; // @[executor.scala 473:84]
  wire [7:0] _GEN_1440 = _GEN_8530 == 8'h33 ? _GEN_1436 : _GEN_976; // @[executor.scala 473:84]
  wire [7:0] _GEN_1441 = _GEN_8530 == 8'h33 ? _GEN_1437 : _GEN_977; // @[executor.scala 473:84]
  wire [7:0] _GEN_1442 = mask_1[0] ? byte_256 : _GEN_978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1443 = mask_1[1] ? byte_257 : _GEN_979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1444 = mask_1[2] ? byte_258 : _GEN_980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1445 = mask_1[3] ? byte_259 : _GEN_981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1446 = _GEN_8530 == 8'h34 ? _GEN_1442 : _GEN_978; // @[executor.scala 473:84]
  wire [7:0] _GEN_1447 = _GEN_8530 == 8'h34 ? _GEN_1443 : _GEN_979; // @[executor.scala 473:84]
  wire [7:0] _GEN_1448 = _GEN_8530 == 8'h34 ? _GEN_1444 : _GEN_980; // @[executor.scala 473:84]
  wire [7:0] _GEN_1449 = _GEN_8530 == 8'h34 ? _GEN_1445 : _GEN_981; // @[executor.scala 473:84]
  wire [7:0] _GEN_1450 = mask_1[0] ? byte_256 : _GEN_982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1451 = mask_1[1] ? byte_257 : _GEN_983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1452 = mask_1[2] ? byte_258 : _GEN_984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1453 = mask_1[3] ? byte_259 : _GEN_985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1454 = _GEN_8530 == 8'h35 ? _GEN_1450 : _GEN_982; // @[executor.scala 473:84]
  wire [7:0] _GEN_1455 = _GEN_8530 == 8'h35 ? _GEN_1451 : _GEN_983; // @[executor.scala 473:84]
  wire [7:0] _GEN_1456 = _GEN_8530 == 8'h35 ? _GEN_1452 : _GEN_984; // @[executor.scala 473:84]
  wire [7:0] _GEN_1457 = _GEN_8530 == 8'h35 ? _GEN_1453 : _GEN_985; // @[executor.scala 473:84]
  wire [7:0] _GEN_1458 = mask_1[0] ? byte_256 : _GEN_986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1459 = mask_1[1] ? byte_257 : _GEN_987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1460 = mask_1[2] ? byte_258 : _GEN_988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1461 = mask_1[3] ? byte_259 : _GEN_989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1462 = _GEN_8530 == 8'h36 ? _GEN_1458 : _GEN_986; // @[executor.scala 473:84]
  wire [7:0] _GEN_1463 = _GEN_8530 == 8'h36 ? _GEN_1459 : _GEN_987; // @[executor.scala 473:84]
  wire [7:0] _GEN_1464 = _GEN_8530 == 8'h36 ? _GEN_1460 : _GEN_988; // @[executor.scala 473:84]
  wire [7:0] _GEN_1465 = _GEN_8530 == 8'h36 ? _GEN_1461 : _GEN_989; // @[executor.scala 473:84]
  wire [7:0] _GEN_1466 = mask_1[0] ? byte_256 : _GEN_990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1467 = mask_1[1] ? byte_257 : _GEN_991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1468 = mask_1[2] ? byte_258 : _GEN_992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1469 = mask_1[3] ? byte_259 : _GEN_993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1470 = _GEN_8530 == 8'h37 ? _GEN_1466 : _GEN_990; // @[executor.scala 473:84]
  wire [7:0] _GEN_1471 = _GEN_8530 == 8'h37 ? _GEN_1467 : _GEN_991; // @[executor.scala 473:84]
  wire [7:0] _GEN_1472 = _GEN_8530 == 8'h37 ? _GEN_1468 : _GEN_992; // @[executor.scala 473:84]
  wire [7:0] _GEN_1473 = _GEN_8530 == 8'h37 ? _GEN_1469 : _GEN_993; // @[executor.scala 473:84]
  wire [7:0] _GEN_1474 = mask_1[0] ? byte_256 : _GEN_994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1475 = mask_1[1] ? byte_257 : _GEN_995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1476 = mask_1[2] ? byte_258 : _GEN_996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1477 = mask_1[3] ? byte_259 : _GEN_997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1478 = _GEN_8530 == 8'h38 ? _GEN_1474 : _GEN_994; // @[executor.scala 473:84]
  wire [7:0] _GEN_1479 = _GEN_8530 == 8'h38 ? _GEN_1475 : _GEN_995; // @[executor.scala 473:84]
  wire [7:0] _GEN_1480 = _GEN_8530 == 8'h38 ? _GEN_1476 : _GEN_996; // @[executor.scala 473:84]
  wire [7:0] _GEN_1481 = _GEN_8530 == 8'h38 ? _GEN_1477 : _GEN_997; // @[executor.scala 473:84]
  wire [7:0] _GEN_1482 = mask_1[0] ? byte_256 : _GEN_998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1483 = mask_1[1] ? byte_257 : _GEN_999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1484 = mask_1[2] ? byte_258 : _GEN_1000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1485 = mask_1[3] ? byte_259 : _GEN_1001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1486 = _GEN_8530 == 8'h39 ? _GEN_1482 : _GEN_998; // @[executor.scala 473:84]
  wire [7:0] _GEN_1487 = _GEN_8530 == 8'h39 ? _GEN_1483 : _GEN_999; // @[executor.scala 473:84]
  wire [7:0] _GEN_1488 = _GEN_8530 == 8'h39 ? _GEN_1484 : _GEN_1000; // @[executor.scala 473:84]
  wire [7:0] _GEN_1489 = _GEN_8530 == 8'h39 ? _GEN_1485 : _GEN_1001; // @[executor.scala 473:84]
  wire [7:0] _GEN_1490 = mask_1[0] ? byte_256 : _GEN_1002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1491 = mask_1[1] ? byte_257 : _GEN_1003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1492 = mask_1[2] ? byte_258 : _GEN_1004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1493 = mask_1[3] ? byte_259 : _GEN_1005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1494 = _GEN_8530 == 8'h3a ? _GEN_1490 : _GEN_1002; // @[executor.scala 473:84]
  wire [7:0] _GEN_1495 = _GEN_8530 == 8'h3a ? _GEN_1491 : _GEN_1003; // @[executor.scala 473:84]
  wire [7:0] _GEN_1496 = _GEN_8530 == 8'h3a ? _GEN_1492 : _GEN_1004; // @[executor.scala 473:84]
  wire [7:0] _GEN_1497 = _GEN_8530 == 8'h3a ? _GEN_1493 : _GEN_1005; // @[executor.scala 473:84]
  wire [7:0] _GEN_1498 = mask_1[0] ? byte_256 : _GEN_1006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1499 = mask_1[1] ? byte_257 : _GEN_1007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1500 = mask_1[2] ? byte_258 : _GEN_1008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1501 = mask_1[3] ? byte_259 : _GEN_1009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1502 = _GEN_8530 == 8'h3b ? _GEN_1498 : _GEN_1006; // @[executor.scala 473:84]
  wire [7:0] _GEN_1503 = _GEN_8530 == 8'h3b ? _GEN_1499 : _GEN_1007; // @[executor.scala 473:84]
  wire [7:0] _GEN_1504 = _GEN_8530 == 8'h3b ? _GEN_1500 : _GEN_1008; // @[executor.scala 473:84]
  wire [7:0] _GEN_1505 = _GEN_8530 == 8'h3b ? _GEN_1501 : _GEN_1009; // @[executor.scala 473:84]
  wire [7:0] _GEN_1506 = mask_1[0] ? byte_256 : _GEN_1010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1507 = mask_1[1] ? byte_257 : _GEN_1011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1508 = mask_1[2] ? byte_258 : _GEN_1012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1509 = mask_1[3] ? byte_259 : _GEN_1013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1510 = _GEN_8530 == 8'h3c ? _GEN_1506 : _GEN_1010; // @[executor.scala 473:84]
  wire [7:0] _GEN_1511 = _GEN_8530 == 8'h3c ? _GEN_1507 : _GEN_1011; // @[executor.scala 473:84]
  wire [7:0] _GEN_1512 = _GEN_8530 == 8'h3c ? _GEN_1508 : _GEN_1012; // @[executor.scala 473:84]
  wire [7:0] _GEN_1513 = _GEN_8530 == 8'h3c ? _GEN_1509 : _GEN_1013; // @[executor.scala 473:84]
  wire [7:0] _GEN_1514 = mask_1[0] ? byte_256 : _GEN_1014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1515 = mask_1[1] ? byte_257 : _GEN_1015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1516 = mask_1[2] ? byte_258 : _GEN_1016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1517 = mask_1[3] ? byte_259 : _GEN_1017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1518 = _GEN_8530 == 8'h3d ? _GEN_1514 : _GEN_1014; // @[executor.scala 473:84]
  wire [7:0] _GEN_1519 = _GEN_8530 == 8'h3d ? _GEN_1515 : _GEN_1015; // @[executor.scala 473:84]
  wire [7:0] _GEN_1520 = _GEN_8530 == 8'h3d ? _GEN_1516 : _GEN_1016; // @[executor.scala 473:84]
  wire [7:0] _GEN_1521 = _GEN_8530 == 8'h3d ? _GEN_1517 : _GEN_1017; // @[executor.scala 473:84]
  wire [7:0] _GEN_1522 = mask_1[0] ? byte_256 : _GEN_1018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1523 = mask_1[1] ? byte_257 : _GEN_1019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1524 = mask_1[2] ? byte_258 : _GEN_1020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1525 = mask_1[3] ? byte_259 : _GEN_1021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1526 = _GEN_8530 == 8'h3e ? _GEN_1522 : _GEN_1018; // @[executor.scala 473:84]
  wire [7:0] _GEN_1527 = _GEN_8530 == 8'h3e ? _GEN_1523 : _GEN_1019; // @[executor.scala 473:84]
  wire [7:0] _GEN_1528 = _GEN_8530 == 8'h3e ? _GEN_1524 : _GEN_1020; // @[executor.scala 473:84]
  wire [7:0] _GEN_1529 = _GEN_8530 == 8'h3e ? _GEN_1525 : _GEN_1021; // @[executor.scala 473:84]
  wire [7:0] _GEN_1530 = mask_1[0] ? byte_256 : _GEN_1022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1531 = mask_1[1] ? byte_257 : _GEN_1023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1532 = mask_1[2] ? byte_258 : _GEN_1024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1533 = mask_1[3] ? byte_259 : _GEN_1025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_1534 = _GEN_8530 == 8'h3f ? _GEN_1530 : _GEN_1022; // @[executor.scala 473:84]
  wire [7:0] _GEN_1535 = _GEN_8530 == 8'h3f ? _GEN_1531 : _GEN_1023; // @[executor.scala 473:84]
  wire [7:0] _GEN_1536 = _GEN_8530 == 8'h3f ? _GEN_1532 : _GEN_1024; // @[executor.scala 473:84]
  wire [7:0] _GEN_1537 = _GEN_8530 == 8'h3f ? _GEN_1533 : _GEN_1025; // @[executor.scala 473:84]
  wire [7:0] _GEN_1538 = opcode_1 != 4'h0 ? _GEN_1030 : _GEN_770; // @[executor.scala 470:55]
  wire [7:0] _GEN_1539 = opcode_1 != 4'h0 ? _GEN_1031 : _GEN_771; // @[executor.scala 470:55]
  wire [7:0] _GEN_1540 = opcode_1 != 4'h0 ? _GEN_1032 : _GEN_772; // @[executor.scala 470:55]
  wire [7:0] _GEN_1541 = opcode_1 != 4'h0 ? _GEN_1033 : _GEN_773; // @[executor.scala 470:55]
  wire [7:0] _GEN_1542 = opcode_1 != 4'h0 ? _GEN_1038 : _GEN_774; // @[executor.scala 470:55]
  wire [7:0] _GEN_1543 = opcode_1 != 4'h0 ? _GEN_1039 : _GEN_775; // @[executor.scala 470:55]
  wire [7:0] _GEN_1544 = opcode_1 != 4'h0 ? _GEN_1040 : _GEN_776; // @[executor.scala 470:55]
  wire [7:0] _GEN_1545 = opcode_1 != 4'h0 ? _GEN_1041 : _GEN_777; // @[executor.scala 470:55]
  wire [7:0] _GEN_1546 = opcode_1 != 4'h0 ? _GEN_1046 : _GEN_778; // @[executor.scala 470:55]
  wire [7:0] _GEN_1547 = opcode_1 != 4'h0 ? _GEN_1047 : _GEN_779; // @[executor.scala 470:55]
  wire [7:0] _GEN_1548 = opcode_1 != 4'h0 ? _GEN_1048 : _GEN_780; // @[executor.scala 470:55]
  wire [7:0] _GEN_1549 = opcode_1 != 4'h0 ? _GEN_1049 : _GEN_781; // @[executor.scala 470:55]
  wire [7:0] _GEN_1550 = opcode_1 != 4'h0 ? _GEN_1054 : _GEN_782; // @[executor.scala 470:55]
  wire [7:0] _GEN_1551 = opcode_1 != 4'h0 ? _GEN_1055 : _GEN_783; // @[executor.scala 470:55]
  wire [7:0] _GEN_1552 = opcode_1 != 4'h0 ? _GEN_1056 : _GEN_784; // @[executor.scala 470:55]
  wire [7:0] _GEN_1553 = opcode_1 != 4'h0 ? _GEN_1057 : _GEN_785; // @[executor.scala 470:55]
  wire [7:0] _GEN_1554 = opcode_1 != 4'h0 ? _GEN_1062 : _GEN_786; // @[executor.scala 470:55]
  wire [7:0] _GEN_1555 = opcode_1 != 4'h0 ? _GEN_1063 : _GEN_787; // @[executor.scala 470:55]
  wire [7:0] _GEN_1556 = opcode_1 != 4'h0 ? _GEN_1064 : _GEN_788; // @[executor.scala 470:55]
  wire [7:0] _GEN_1557 = opcode_1 != 4'h0 ? _GEN_1065 : _GEN_789; // @[executor.scala 470:55]
  wire [7:0] _GEN_1558 = opcode_1 != 4'h0 ? _GEN_1070 : _GEN_790; // @[executor.scala 470:55]
  wire [7:0] _GEN_1559 = opcode_1 != 4'h0 ? _GEN_1071 : _GEN_791; // @[executor.scala 470:55]
  wire [7:0] _GEN_1560 = opcode_1 != 4'h0 ? _GEN_1072 : _GEN_792; // @[executor.scala 470:55]
  wire [7:0] _GEN_1561 = opcode_1 != 4'h0 ? _GEN_1073 : _GEN_793; // @[executor.scala 470:55]
  wire [7:0] _GEN_1562 = opcode_1 != 4'h0 ? _GEN_1078 : _GEN_794; // @[executor.scala 470:55]
  wire [7:0] _GEN_1563 = opcode_1 != 4'h0 ? _GEN_1079 : _GEN_795; // @[executor.scala 470:55]
  wire [7:0] _GEN_1564 = opcode_1 != 4'h0 ? _GEN_1080 : _GEN_796; // @[executor.scala 470:55]
  wire [7:0] _GEN_1565 = opcode_1 != 4'h0 ? _GEN_1081 : _GEN_797; // @[executor.scala 470:55]
  wire [7:0] _GEN_1566 = opcode_1 != 4'h0 ? _GEN_1086 : _GEN_798; // @[executor.scala 470:55]
  wire [7:0] _GEN_1567 = opcode_1 != 4'h0 ? _GEN_1087 : _GEN_799; // @[executor.scala 470:55]
  wire [7:0] _GEN_1568 = opcode_1 != 4'h0 ? _GEN_1088 : _GEN_800; // @[executor.scala 470:55]
  wire [7:0] _GEN_1569 = opcode_1 != 4'h0 ? _GEN_1089 : _GEN_801; // @[executor.scala 470:55]
  wire [7:0] _GEN_1570 = opcode_1 != 4'h0 ? _GEN_1094 : _GEN_802; // @[executor.scala 470:55]
  wire [7:0] _GEN_1571 = opcode_1 != 4'h0 ? _GEN_1095 : _GEN_803; // @[executor.scala 470:55]
  wire [7:0] _GEN_1572 = opcode_1 != 4'h0 ? _GEN_1096 : _GEN_804; // @[executor.scala 470:55]
  wire [7:0] _GEN_1573 = opcode_1 != 4'h0 ? _GEN_1097 : _GEN_805; // @[executor.scala 470:55]
  wire [7:0] _GEN_1574 = opcode_1 != 4'h0 ? _GEN_1102 : _GEN_806; // @[executor.scala 470:55]
  wire [7:0] _GEN_1575 = opcode_1 != 4'h0 ? _GEN_1103 : _GEN_807; // @[executor.scala 470:55]
  wire [7:0] _GEN_1576 = opcode_1 != 4'h0 ? _GEN_1104 : _GEN_808; // @[executor.scala 470:55]
  wire [7:0] _GEN_1577 = opcode_1 != 4'h0 ? _GEN_1105 : _GEN_809; // @[executor.scala 470:55]
  wire [7:0] _GEN_1578 = opcode_1 != 4'h0 ? _GEN_1110 : _GEN_810; // @[executor.scala 470:55]
  wire [7:0] _GEN_1579 = opcode_1 != 4'h0 ? _GEN_1111 : _GEN_811; // @[executor.scala 470:55]
  wire [7:0] _GEN_1580 = opcode_1 != 4'h0 ? _GEN_1112 : _GEN_812; // @[executor.scala 470:55]
  wire [7:0] _GEN_1581 = opcode_1 != 4'h0 ? _GEN_1113 : _GEN_813; // @[executor.scala 470:55]
  wire [7:0] _GEN_1582 = opcode_1 != 4'h0 ? _GEN_1118 : _GEN_814; // @[executor.scala 470:55]
  wire [7:0] _GEN_1583 = opcode_1 != 4'h0 ? _GEN_1119 : _GEN_815; // @[executor.scala 470:55]
  wire [7:0] _GEN_1584 = opcode_1 != 4'h0 ? _GEN_1120 : _GEN_816; // @[executor.scala 470:55]
  wire [7:0] _GEN_1585 = opcode_1 != 4'h0 ? _GEN_1121 : _GEN_817; // @[executor.scala 470:55]
  wire [7:0] _GEN_1586 = opcode_1 != 4'h0 ? _GEN_1126 : _GEN_818; // @[executor.scala 470:55]
  wire [7:0] _GEN_1587 = opcode_1 != 4'h0 ? _GEN_1127 : _GEN_819; // @[executor.scala 470:55]
  wire [7:0] _GEN_1588 = opcode_1 != 4'h0 ? _GEN_1128 : _GEN_820; // @[executor.scala 470:55]
  wire [7:0] _GEN_1589 = opcode_1 != 4'h0 ? _GEN_1129 : _GEN_821; // @[executor.scala 470:55]
  wire [7:0] _GEN_1590 = opcode_1 != 4'h0 ? _GEN_1134 : _GEN_822; // @[executor.scala 470:55]
  wire [7:0] _GEN_1591 = opcode_1 != 4'h0 ? _GEN_1135 : _GEN_823; // @[executor.scala 470:55]
  wire [7:0] _GEN_1592 = opcode_1 != 4'h0 ? _GEN_1136 : _GEN_824; // @[executor.scala 470:55]
  wire [7:0] _GEN_1593 = opcode_1 != 4'h0 ? _GEN_1137 : _GEN_825; // @[executor.scala 470:55]
  wire [7:0] _GEN_1594 = opcode_1 != 4'h0 ? _GEN_1142 : _GEN_826; // @[executor.scala 470:55]
  wire [7:0] _GEN_1595 = opcode_1 != 4'h0 ? _GEN_1143 : _GEN_827; // @[executor.scala 470:55]
  wire [7:0] _GEN_1596 = opcode_1 != 4'h0 ? _GEN_1144 : _GEN_828; // @[executor.scala 470:55]
  wire [7:0] _GEN_1597 = opcode_1 != 4'h0 ? _GEN_1145 : _GEN_829; // @[executor.scala 470:55]
  wire [7:0] _GEN_1598 = opcode_1 != 4'h0 ? _GEN_1150 : _GEN_830; // @[executor.scala 470:55]
  wire [7:0] _GEN_1599 = opcode_1 != 4'h0 ? _GEN_1151 : _GEN_831; // @[executor.scala 470:55]
  wire [7:0] _GEN_1600 = opcode_1 != 4'h0 ? _GEN_1152 : _GEN_832; // @[executor.scala 470:55]
  wire [7:0] _GEN_1601 = opcode_1 != 4'h0 ? _GEN_1153 : _GEN_833; // @[executor.scala 470:55]
  wire [7:0] _GEN_1602 = opcode_1 != 4'h0 ? _GEN_1158 : _GEN_834; // @[executor.scala 470:55]
  wire [7:0] _GEN_1603 = opcode_1 != 4'h0 ? _GEN_1159 : _GEN_835; // @[executor.scala 470:55]
  wire [7:0] _GEN_1604 = opcode_1 != 4'h0 ? _GEN_1160 : _GEN_836; // @[executor.scala 470:55]
  wire [7:0] _GEN_1605 = opcode_1 != 4'h0 ? _GEN_1161 : _GEN_837; // @[executor.scala 470:55]
  wire [7:0] _GEN_1606 = opcode_1 != 4'h0 ? _GEN_1166 : _GEN_838; // @[executor.scala 470:55]
  wire [7:0] _GEN_1607 = opcode_1 != 4'h0 ? _GEN_1167 : _GEN_839; // @[executor.scala 470:55]
  wire [7:0] _GEN_1608 = opcode_1 != 4'h0 ? _GEN_1168 : _GEN_840; // @[executor.scala 470:55]
  wire [7:0] _GEN_1609 = opcode_1 != 4'h0 ? _GEN_1169 : _GEN_841; // @[executor.scala 470:55]
  wire [7:0] _GEN_1610 = opcode_1 != 4'h0 ? _GEN_1174 : _GEN_842; // @[executor.scala 470:55]
  wire [7:0] _GEN_1611 = opcode_1 != 4'h0 ? _GEN_1175 : _GEN_843; // @[executor.scala 470:55]
  wire [7:0] _GEN_1612 = opcode_1 != 4'h0 ? _GEN_1176 : _GEN_844; // @[executor.scala 470:55]
  wire [7:0] _GEN_1613 = opcode_1 != 4'h0 ? _GEN_1177 : _GEN_845; // @[executor.scala 470:55]
  wire [7:0] _GEN_1614 = opcode_1 != 4'h0 ? _GEN_1182 : _GEN_846; // @[executor.scala 470:55]
  wire [7:0] _GEN_1615 = opcode_1 != 4'h0 ? _GEN_1183 : _GEN_847; // @[executor.scala 470:55]
  wire [7:0] _GEN_1616 = opcode_1 != 4'h0 ? _GEN_1184 : _GEN_848; // @[executor.scala 470:55]
  wire [7:0] _GEN_1617 = opcode_1 != 4'h0 ? _GEN_1185 : _GEN_849; // @[executor.scala 470:55]
  wire [7:0] _GEN_1618 = opcode_1 != 4'h0 ? _GEN_1190 : _GEN_850; // @[executor.scala 470:55]
  wire [7:0] _GEN_1619 = opcode_1 != 4'h0 ? _GEN_1191 : _GEN_851; // @[executor.scala 470:55]
  wire [7:0] _GEN_1620 = opcode_1 != 4'h0 ? _GEN_1192 : _GEN_852; // @[executor.scala 470:55]
  wire [7:0] _GEN_1621 = opcode_1 != 4'h0 ? _GEN_1193 : _GEN_853; // @[executor.scala 470:55]
  wire [7:0] _GEN_1622 = opcode_1 != 4'h0 ? _GEN_1198 : _GEN_854; // @[executor.scala 470:55]
  wire [7:0] _GEN_1623 = opcode_1 != 4'h0 ? _GEN_1199 : _GEN_855; // @[executor.scala 470:55]
  wire [7:0] _GEN_1624 = opcode_1 != 4'h0 ? _GEN_1200 : _GEN_856; // @[executor.scala 470:55]
  wire [7:0] _GEN_1625 = opcode_1 != 4'h0 ? _GEN_1201 : _GEN_857; // @[executor.scala 470:55]
  wire [7:0] _GEN_1626 = opcode_1 != 4'h0 ? _GEN_1206 : _GEN_858; // @[executor.scala 470:55]
  wire [7:0] _GEN_1627 = opcode_1 != 4'h0 ? _GEN_1207 : _GEN_859; // @[executor.scala 470:55]
  wire [7:0] _GEN_1628 = opcode_1 != 4'h0 ? _GEN_1208 : _GEN_860; // @[executor.scala 470:55]
  wire [7:0] _GEN_1629 = opcode_1 != 4'h0 ? _GEN_1209 : _GEN_861; // @[executor.scala 470:55]
  wire [7:0] _GEN_1630 = opcode_1 != 4'h0 ? _GEN_1214 : _GEN_862; // @[executor.scala 470:55]
  wire [7:0] _GEN_1631 = opcode_1 != 4'h0 ? _GEN_1215 : _GEN_863; // @[executor.scala 470:55]
  wire [7:0] _GEN_1632 = opcode_1 != 4'h0 ? _GEN_1216 : _GEN_864; // @[executor.scala 470:55]
  wire [7:0] _GEN_1633 = opcode_1 != 4'h0 ? _GEN_1217 : _GEN_865; // @[executor.scala 470:55]
  wire [7:0] _GEN_1634 = opcode_1 != 4'h0 ? _GEN_1222 : _GEN_866; // @[executor.scala 470:55]
  wire [7:0] _GEN_1635 = opcode_1 != 4'h0 ? _GEN_1223 : _GEN_867; // @[executor.scala 470:55]
  wire [7:0] _GEN_1636 = opcode_1 != 4'h0 ? _GEN_1224 : _GEN_868; // @[executor.scala 470:55]
  wire [7:0] _GEN_1637 = opcode_1 != 4'h0 ? _GEN_1225 : _GEN_869; // @[executor.scala 470:55]
  wire [7:0] _GEN_1638 = opcode_1 != 4'h0 ? _GEN_1230 : _GEN_870; // @[executor.scala 470:55]
  wire [7:0] _GEN_1639 = opcode_1 != 4'h0 ? _GEN_1231 : _GEN_871; // @[executor.scala 470:55]
  wire [7:0] _GEN_1640 = opcode_1 != 4'h0 ? _GEN_1232 : _GEN_872; // @[executor.scala 470:55]
  wire [7:0] _GEN_1641 = opcode_1 != 4'h0 ? _GEN_1233 : _GEN_873; // @[executor.scala 470:55]
  wire [7:0] _GEN_1642 = opcode_1 != 4'h0 ? _GEN_1238 : _GEN_874; // @[executor.scala 470:55]
  wire [7:0] _GEN_1643 = opcode_1 != 4'h0 ? _GEN_1239 : _GEN_875; // @[executor.scala 470:55]
  wire [7:0] _GEN_1644 = opcode_1 != 4'h0 ? _GEN_1240 : _GEN_876; // @[executor.scala 470:55]
  wire [7:0] _GEN_1645 = opcode_1 != 4'h0 ? _GEN_1241 : _GEN_877; // @[executor.scala 470:55]
  wire [7:0] _GEN_1646 = opcode_1 != 4'h0 ? _GEN_1246 : _GEN_878; // @[executor.scala 470:55]
  wire [7:0] _GEN_1647 = opcode_1 != 4'h0 ? _GEN_1247 : _GEN_879; // @[executor.scala 470:55]
  wire [7:0] _GEN_1648 = opcode_1 != 4'h0 ? _GEN_1248 : _GEN_880; // @[executor.scala 470:55]
  wire [7:0] _GEN_1649 = opcode_1 != 4'h0 ? _GEN_1249 : _GEN_881; // @[executor.scala 470:55]
  wire [7:0] _GEN_1650 = opcode_1 != 4'h0 ? _GEN_1254 : _GEN_882; // @[executor.scala 470:55]
  wire [7:0] _GEN_1651 = opcode_1 != 4'h0 ? _GEN_1255 : _GEN_883; // @[executor.scala 470:55]
  wire [7:0] _GEN_1652 = opcode_1 != 4'h0 ? _GEN_1256 : _GEN_884; // @[executor.scala 470:55]
  wire [7:0] _GEN_1653 = opcode_1 != 4'h0 ? _GEN_1257 : _GEN_885; // @[executor.scala 470:55]
  wire [7:0] _GEN_1654 = opcode_1 != 4'h0 ? _GEN_1262 : _GEN_886; // @[executor.scala 470:55]
  wire [7:0] _GEN_1655 = opcode_1 != 4'h0 ? _GEN_1263 : _GEN_887; // @[executor.scala 470:55]
  wire [7:0] _GEN_1656 = opcode_1 != 4'h0 ? _GEN_1264 : _GEN_888; // @[executor.scala 470:55]
  wire [7:0] _GEN_1657 = opcode_1 != 4'h0 ? _GEN_1265 : _GEN_889; // @[executor.scala 470:55]
  wire [7:0] _GEN_1658 = opcode_1 != 4'h0 ? _GEN_1270 : _GEN_890; // @[executor.scala 470:55]
  wire [7:0] _GEN_1659 = opcode_1 != 4'h0 ? _GEN_1271 : _GEN_891; // @[executor.scala 470:55]
  wire [7:0] _GEN_1660 = opcode_1 != 4'h0 ? _GEN_1272 : _GEN_892; // @[executor.scala 470:55]
  wire [7:0] _GEN_1661 = opcode_1 != 4'h0 ? _GEN_1273 : _GEN_893; // @[executor.scala 470:55]
  wire [7:0] _GEN_1662 = opcode_1 != 4'h0 ? _GEN_1278 : _GEN_894; // @[executor.scala 470:55]
  wire [7:0] _GEN_1663 = opcode_1 != 4'h0 ? _GEN_1279 : _GEN_895; // @[executor.scala 470:55]
  wire [7:0] _GEN_1664 = opcode_1 != 4'h0 ? _GEN_1280 : _GEN_896; // @[executor.scala 470:55]
  wire [7:0] _GEN_1665 = opcode_1 != 4'h0 ? _GEN_1281 : _GEN_897; // @[executor.scala 470:55]
  wire [7:0] _GEN_1666 = opcode_1 != 4'h0 ? _GEN_1286 : _GEN_898; // @[executor.scala 470:55]
  wire [7:0] _GEN_1667 = opcode_1 != 4'h0 ? _GEN_1287 : _GEN_899; // @[executor.scala 470:55]
  wire [7:0] _GEN_1668 = opcode_1 != 4'h0 ? _GEN_1288 : _GEN_900; // @[executor.scala 470:55]
  wire [7:0] _GEN_1669 = opcode_1 != 4'h0 ? _GEN_1289 : _GEN_901; // @[executor.scala 470:55]
  wire [7:0] _GEN_1670 = opcode_1 != 4'h0 ? _GEN_1294 : _GEN_902; // @[executor.scala 470:55]
  wire [7:0] _GEN_1671 = opcode_1 != 4'h0 ? _GEN_1295 : _GEN_903; // @[executor.scala 470:55]
  wire [7:0] _GEN_1672 = opcode_1 != 4'h0 ? _GEN_1296 : _GEN_904; // @[executor.scala 470:55]
  wire [7:0] _GEN_1673 = opcode_1 != 4'h0 ? _GEN_1297 : _GEN_905; // @[executor.scala 470:55]
  wire [7:0] _GEN_1674 = opcode_1 != 4'h0 ? _GEN_1302 : _GEN_906; // @[executor.scala 470:55]
  wire [7:0] _GEN_1675 = opcode_1 != 4'h0 ? _GEN_1303 : _GEN_907; // @[executor.scala 470:55]
  wire [7:0] _GEN_1676 = opcode_1 != 4'h0 ? _GEN_1304 : _GEN_908; // @[executor.scala 470:55]
  wire [7:0] _GEN_1677 = opcode_1 != 4'h0 ? _GEN_1305 : _GEN_909; // @[executor.scala 470:55]
  wire [7:0] _GEN_1678 = opcode_1 != 4'h0 ? _GEN_1310 : _GEN_910; // @[executor.scala 470:55]
  wire [7:0] _GEN_1679 = opcode_1 != 4'h0 ? _GEN_1311 : _GEN_911; // @[executor.scala 470:55]
  wire [7:0] _GEN_1680 = opcode_1 != 4'h0 ? _GEN_1312 : _GEN_912; // @[executor.scala 470:55]
  wire [7:0] _GEN_1681 = opcode_1 != 4'h0 ? _GEN_1313 : _GEN_913; // @[executor.scala 470:55]
  wire [7:0] _GEN_1682 = opcode_1 != 4'h0 ? _GEN_1318 : _GEN_914; // @[executor.scala 470:55]
  wire [7:0] _GEN_1683 = opcode_1 != 4'h0 ? _GEN_1319 : _GEN_915; // @[executor.scala 470:55]
  wire [7:0] _GEN_1684 = opcode_1 != 4'h0 ? _GEN_1320 : _GEN_916; // @[executor.scala 470:55]
  wire [7:0] _GEN_1685 = opcode_1 != 4'h0 ? _GEN_1321 : _GEN_917; // @[executor.scala 470:55]
  wire [7:0] _GEN_1686 = opcode_1 != 4'h0 ? _GEN_1326 : _GEN_918; // @[executor.scala 470:55]
  wire [7:0] _GEN_1687 = opcode_1 != 4'h0 ? _GEN_1327 : _GEN_919; // @[executor.scala 470:55]
  wire [7:0] _GEN_1688 = opcode_1 != 4'h0 ? _GEN_1328 : _GEN_920; // @[executor.scala 470:55]
  wire [7:0] _GEN_1689 = opcode_1 != 4'h0 ? _GEN_1329 : _GEN_921; // @[executor.scala 470:55]
  wire [7:0] _GEN_1690 = opcode_1 != 4'h0 ? _GEN_1334 : _GEN_922; // @[executor.scala 470:55]
  wire [7:0] _GEN_1691 = opcode_1 != 4'h0 ? _GEN_1335 : _GEN_923; // @[executor.scala 470:55]
  wire [7:0] _GEN_1692 = opcode_1 != 4'h0 ? _GEN_1336 : _GEN_924; // @[executor.scala 470:55]
  wire [7:0] _GEN_1693 = opcode_1 != 4'h0 ? _GEN_1337 : _GEN_925; // @[executor.scala 470:55]
  wire [7:0] _GEN_1694 = opcode_1 != 4'h0 ? _GEN_1342 : _GEN_926; // @[executor.scala 470:55]
  wire [7:0] _GEN_1695 = opcode_1 != 4'h0 ? _GEN_1343 : _GEN_927; // @[executor.scala 470:55]
  wire [7:0] _GEN_1696 = opcode_1 != 4'h0 ? _GEN_1344 : _GEN_928; // @[executor.scala 470:55]
  wire [7:0] _GEN_1697 = opcode_1 != 4'h0 ? _GEN_1345 : _GEN_929; // @[executor.scala 470:55]
  wire [7:0] _GEN_1698 = opcode_1 != 4'h0 ? _GEN_1350 : _GEN_930; // @[executor.scala 470:55]
  wire [7:0] _GEN_1699 = opcode_1 != 4'h0 ? _GEN_1351 : _GEN_931; // @[executor.scala 470:55]
  wire [7:0] _GEN_1700 = opcode_1 != 4'h0 ? _GEN_1352 : _GEN_932; // @[executor.scala 470:55]
  wire [7:0] _GEN_1701 = opcode_1 != 4'h0 ? _GEN_1353 : _GEN_933; // @[executor.scala 470:55]
  wire [7:0] _GEN_1702 = opcode_1 != 4'h0 ? _GEN_1358 : _GEN_934; // @[executor.scala 470:55]
  wire [7:0] _GEN_1703 = opcode_1 != 4'h0 ? _GEN_1359 : _GEN_935; // @[executor.scala 470:55]
  wire [7:0] _GEN_1704 = opcode_1 != 4'h0 ? _GEN_1360 : _GEN_936; // @[executor.scala 470:55]
  wire [7:0] _GEN_1705 = opcode_1 != 4'h0 ? _GEN_1361 : _GEN_937; // @[executor.scala 470:55]
  wire [7:0] _GEN_1706 = opcode_1 != 4'h0 ? _GEN_1366 : _GEN_938; // @[executor.scala 470:55]
  wire [7:0] _GEN_1707 = opcode_1 != 4'h0 ? _GEN_1367 : _GEN_939; // @[executor.scala 470:55]
  wire [7:0] _GEN_1708 = opcode_1 != 4'h0 ? _GEN_1368 : _GEN_940; // @[executor.scala 470:55]
  wire [7:0] _GEN_1709 = opcode_1 != 4'h0 ? _GEN_1369 : _GEN_941; // @[executor.scala 470:55]
  wire [7:0] _GEN_1710 = opcode_1 != 4'h0 ? _GEN_1374 : _GEN_942; // @[executor.scala 470:55]
  wire [7:0] _GEN_1711 = opcode_1 != 4'h0 ? _GEN_1375 : _GEN_943; // @[executor.scala 470:55]
  wire [7:0] _GEN_1712 = opcode_1 != 4'h0 ? _GEN_1376 : _GEN_944; // @[executor.scala 470:55]
  wire [7:0] _GEN_1713 = opcode_1 != 4'h0 ? _GEN_1377 : _GEN_945; // @[executor.scala 470:55]
  wire [7:0] _GEN_1714 = opcode_1 != 4'h0 ? _GEN_1382 : _GEN_946; // @[executor.scala 470:55]
  wire [7:0] _GEN_1715 = opcode_1 != 4'h0 ? _GEN_1383 : _GEN_947; // @[executor.scala 470:55]
  wire [7:0] _GEN_1716 = opcode_1 != 4'h0 ? _GEN_1384 : _GEN_948; // @[executor.scala 470:55]
  wire [7:0] _GEN_1717 = opcode_1 != 4'h0 ? _GEN_1385 : _GEN_949; // @[executor.scala 470:55]
  wire [7:0] _GEN_1718 = opcode_1 != 4'h0 ? _GEN_1390 : _GEN_950; // @[executor.scala 470:55]
  wire [7:0] _GEN_1719 = opcode_1 != 4'h0 ? _GEN_1391 : _GEN_951; // @[executor.scala 470:55]
  wire [7:0] _GEN_1720 = opcode_1 != 4'h0 ? _GEN_1392 : _GEN_952; // @[executor.scala 470:55]
  wire [7:0] _GEN_1721 = opcode_1 != 4'h0 ? _GEN_1393 : _GEN_953; // @[executor.scala 470:55]
  wire [7:0] _GEN_1722 = opcode_1 != 4'h0 ? _GEN_1398 : _GEN_954; // @[executor.scala 470:55]
  wire [7:0] _GEN_1723 = opcode_1 != 4'h0 ? _GEN_1399 : _GEN_955; // @[executor.scala 470:55]
  wire [7:0] _GEN_1724 = opcode_1 != 4'h0 ? _GEN_1400 : _GEN_956; // @[executor.scala 470:55]
  wire [7:0] _GEN_1725 = opcode_1 != 4'h0 ? _GEN_1401 : _GEN_957; // @[executor.scala 470:55]
  wire [7:0] _GEN_1726 = opcode_1 != 4'h0 ? _GEN_1406 : _GEN_958; // @[executor.scala 470:55]
  wire [7:0] _GEN_1727 = opcode_1 != 4'h0 ? _GEN_1407 : _GEN_959; // @[executor.scala 470:55]
  wire [7:0] _GEN_1728 = opcode_1 != 4'h0 ? _GEN_1408 : _GEN_960; // @[executor.scala 470:55]
  wire [7:0] _GEN_1729 = opcode_1 != 4'h0 ? _GEN_1409 : _GEN_961; // @[executor.scala 470:55]
  wire [7:0] _GEN_1730 = opcode_1 != 4'h0 ? _GEN_1414 : _GEN_962; // @[executor.scala 470:55]
  wire [7:0] _GEN_1731 = opcode_1 != 4'h0 ? _GEN_1415 : _GEN_963; // @[executor.scala 470:55]
  wire [7:0] _GEN_1732 = opcode_1 != 4'h0 ? _GEN_1416 : _GEN_964; // @[executor.scala 470:55]
  wire [7:0] _GEN_1733 = opcode_1 != 4'h0 ? _GEN_1417 : _GEN_965; // @[executor.scala 470:55]
  wire [7:0] _GEN_1734 = opcode_1 != 4'h0 ? _GEN_1422 : _GEN_966; // @[executor.scala 470:55]
  wire [7:0] _GEN_1735 = opcode_1 != 4'h0 ? _GEN_1423 : _GEN_967; // @[executor.scala 470:55]
  wire [7:0] _GEN_1736 = opcode_1 != 4'h0 ? _GEN_1424 : _GEN_968; // @[executor.scala 470:55]
  wire [7:0] _GEN_1737 = opcode_1 != 4'h0 ? _GEN_1425 : _GEN_969; // @[executor.scala 470:55]
  wire [7:0] _GEN_1738 = opcode_1 != 4'h0 ? _GEN_1430 : _GEN_970; // @[executor.scala 470:55]
  wire [7:0] _GEN_1739 = opcode_1 != 4'h0 ? _GEN_1431 : _GEN_971; // @[executor.scala 470:55]
  wire [7:0] _GEN_1740 = opcode_1 != 4'h0 ? _GEN_1432 : _GEN_972; // @[executor.scala 470:55]
  wire [7:0] _GEN_1741 = opcode_1 != 4'h0 ? _GEN_1433 : _GEN_973; // @[executor.scala 470:55]
  wire [7:0] _GEN_1742 = opcode_1 != 4'h0 ? _GEN_1438 : _GEN_974; // @[executor.scala 470:55]
  wire [7:0] _GEN_1743 = opcode_1 != 4'h0 ? _GEN_1439 : _GEN_975; // @[executor.scala 470:55]
  wire [7:0] _GEN_1744 = opcode_1 != 4'h0 ? _GEN_1440 : _GEN_976; // @[executor.scala 470:55]
  wire [7:0] _GEN_1745 = opcode_1 != 4'h0 ? _GEN_1441 : _GEN_977; // @[executor.scala 470:55]
  wire [7:0] _GEN_1746 = opcode_1 != 4'h0 ? _GEN_1446 : _GEN_978; // @[executor.scala 470:55]
  wire [7:0] _GEN_1747 = opcode_1 != 4'h0 ? _GEN_1447 : _GEN_979; // @[executor.scala 470:55]
  wire [7:0] _GEN_1748 = opcode_1 != 4'h0 ? _GEN_1448 : _GEN_980; // @[executor.scala 470:55]
  wire [7:0] _GEN_1749 = opcode_1 != 4'h0 ? _GEN_1449 : _GEN_981; // @[executor.scala 470:55]
  wire [7:0] _GEN_1750 = opcode_1 != 4'h0 ? _GEN_1454 : _GEN_982; // @[executor.scala 470:55]
  wire [7:0] _GEN_1751 = opcode_1 != 4'h0 ? _GEN_1455 : _GEN_983; // @[executor.scala 470:55]
  wire [7:0] _GEN_1752 = opcode_1 != 4'h0 ? _GEN_1456 : _GEN_984; // @[executor.scala 470:55]
  wire [7:0] _GEN_1753 = opcode_1 != 4'h0 ? _GEN_1457 : _GEN_985; // @[executor.scala 470:55]
  wire [7:0] _GEN_1754 = opcode_1 != 4'h0 ? _GEN_1462 : _GEN_986; // @[executor.scala 470:55]
  wire [7:0] _GEN_1755 = opcode_1 != 4'h0 ? _GEN_1463 : _GEN_987; // @[executor.scala 470:55]
  wire [7:0] _GEN_1756 = opcode_1 != 4'h0 ? _GEN_1464 : _GEN_988; // @[executor.scala 470:55]
  wire [7:0] _GEN_1757 = opcode_1 != 4'h0 ? _GEN_1465 : _GEN_989; // @[executor.scala 470:55]
  wire [7:0] _GEN_1758 = opcode_1 != 4'h0 ? _GEN_1470 : _GEN_990; // @[executor.scala 470:55]
  wire [7:0] _GEN_1759 = opcode_1 != 4'h0 ? _GEN_1471 : _GEN_991; // @[executor.scala 470:55]
  wire [7:0] _GEN_1760 = opcode_1 != 4'h0 ? _GEN_1472 : _GEN_992; // @[executor.scala 470:55]
  wire [7:0] _GEN_1761 = opcode_1 != 4'h0 ? _GEN_1473 : _GEN_993; // @[executor.scala 470:55]
  wire [7:0] _GEN_1762 = opcode_1 != 4'h0 ? _GEN_1478 : _GEN_994; // @[executor.scala 470:55]
  wire [7:0] _GEN_1763 = opcode_1 != 4'h0 ? _GEN_1479 : _GEN_995; // @[executor.scala 470:55]
  wire [7:0] _GEN_1764 = opcode_1 != 4'h0 ? _GEN_1480 : _GEN_996; // @[executor.scala 470:55]
  wire [7:0] _GEN_1765 = opcode_1 != 4'h0 ? _GEN_1481 : _GEN_997; // @[executor.scala 470:55]
  wire [7:0] _GEN_1766 = opcode_1 != 4'h0 ? _GEN_1486 : _GEN_998; // @[executor.scala 470:55]
  wire [7:0] _GEN_1767 = opcode_1 != 4'h0 ? _GEN_1487 : _GEN_999; // @[executor.scala 470:55]
  wire [7:0] _GEN_1768 = opcode_1 != 4'h0 ? _GEN_1488 : _GEN_1000; // @[executor.scala 470:55]
  wire [7:0] _GEN_1769 = opcode_1 != 4'h0 ? _GEN_1489 : _GEN_1001; // @[executor.scala 470:55]
  wire [7:0] _GEN_1770 = opcode_1 != 4'h0 ? _GEN_1494 : _GEN_1002; // @[executor.scala 470:55]
  wire [7:0] _GEN_1771 = opcode_1 != 4'h0 ? _GEN_1495 : _GEN_1003; // @[executor.scala 470:55]
  wire [7:0] _GEN_1772 = opcode_1 != 4'h0 ? _GEN_1496 : _GEN_1004; // @[executor.scala 470:55]
  wire [7:0] _GEN_1773 = opcode_1 != 4'h0 ? _GEN_1497 : _GEN_1005; // @[executor.scala 470:55]
  wire [7:0] _GEN_1774 = opcode_1 != 4'h0 ? _GEN_1502 : _GEN_1006; // @[executor.scala 470:55]
  wire [7:0] _GEN_1775 = opcode_1 != 4'h0 ? _GEN_1503 : _GEN_1007; // @[executor.scala 470:55]
  wire [7:0] _GEN_1776 = opcode_1 != 4'h0 ? _GEN_1504 : _GEN_1008; // @[executor.scala 470:55]
  wire [7:0] _GEN_1777 = opcode_1 != 4'h0 ? _GEN_1505 : _GEN_1009; // @[executor.scala 470:55]
  wire [7:0] _GEN_1778 = opcode_1 != 4'h0 ? _GEN_1510 : _GEN_1010; // @[executor.scala 470:55]
  wire [7:0] _GEN_1779 = opcode_1 != 4'h0 ? _GEN_1511 : _GEN_1011; // @[executor.scala 470:55]
  wire [7:0] _GEN_1780 = opcode_1 != 4'h0 ? _GEN_1512 : _GEN_1012; // @[executor.scala 470:55]
  wire [7:0] _GEN_1781 = opcode_1 != 4'h0 ? _GEN_1513 : _GEN_1013; // @[executor.scala 470:55]
  wire [7:0] _GEN_1782 = opcode_1 != 4'h0 ? _GEN_1518 : _GEN_1014; // @[executor.scala 470:55]
  wire [7:0] _GEN_1783 = opcode_1 != 4'h0 ? _GEN_1519 : _GEN_1015; // @[executor.scala 470:55]
  wire [7:0] _GEN_1784 = opcode_1 != 4'h0 ? _GEN_1520 : _GEN_1016; // @[executor.scala 470:55]
  wire [7:0] _GEN_1785 = opcode_1 != 4'h0 ? _GEN_1521 : _GEN_1017; // @[executor.scala 470:55]
  wire [7:0] _GEN_1786 = opcode_1 != 4'h0 ? _GEN_1526 : _GEN_1018; // @[executor.scala 470:55]
  wire [7:0] _GEN_1787 = opcode_1 != 4'h0 ? _GEN_1527 : _GEN_1019; // @[executor.scala 470:55]
  wire [7:0] _GEN_1788 = opcode_1 != 4'h0 ? _GEN_1528 : _GEN_1020; // @[executor.scala 470:55]
  wire [7:0] _GEN_1789 = opcode_1 != 4'h0 ? _GEN_1529 : _GEN_1021; // @[executor.scala 470:55]
  wire [7:0] _GEN_1790 = opcode_1 != 4'h0 ? _GEN_1534 : _GEN_1022; // @[executor.scala 470:55]
  wire [7:0] _GEN_1791 = opcode_1 != 4'h0 ? _GEN_1535 : _GEN_1023; // @[executor.scala 470:55]
  wire [7:0] _GEN_1792 = opcode_1 != 4'h0 ? _GEN_1536 : _GEN_1024; // @[executor.scala 470:55]
  wire [7:0] _GEN_1793 = opcode_1 != 4'h0 ? _GEN_1537 : _GEN_1025; // @[executor.scala 470:55]
  wire [3:0] _GEN_1794 = opcode_1 == 4'hf ? parameter_2_1[13:10] : _GEN_768; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_1795 = opcode_1 == 4'hf ? parameter_2_1[0] : _GEN_769; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_1796 = opcode_1 == 4'hf ? _GEN_770 : _GEN_1538; // @[executor.scala 466:52]
  wire [7:0] _GEN_1797 = opcode_1 == 4'hf ? _GEN_771 : _GEN_1539; // @[executor.scala 466:52]
  wire [7:0] _GEN_1798 = opcode_1 == 4'hf ? _GEN_772 : _GEN_1540; // @[executor.scala 466:52]
  wire [7:0] _GEN_1799 = opcode_1 == 4'hf ? _GEN_773 : _GEN_1541; // @[executor.scala 466:52]
  wire [7:0] _GEN_1800 = opcode_1 == 4'hf ? _GEN_774 : _GEN_1542; // @[executor.scala 466:52]
  wire [7:0] _GEN_1801 = opcode_1 == 4'hf ? _GEN_775 : _GEN_1543; // @[executor.scala 466:52]
  wire [7:0] _GEN_1802 = opcode_1 == 4'hf ? _GEN_776 : _GEN_1544; // @[executor.scala 466:52]
  wire [7:0] _GEN_1803 = opcode_1 == 4'hf ? _GEN_777 : _GEN_1545; // @[executor.scala 466:52]
  wire [7:0] _GEN_1804 = opcode_1 == 4'hf ? _GEN_778 : _GEN_1546; // @[executor.scala 466:52]
  wire [7:0] _GEN_1805 = opcode_1 == 4'hf ? _GEN_779 : _GEN_1547; // @[executor.scala 466:52]
  wire [7:0] _GEN_1806 = opcode_1 == 4'hf ? _GEN_780 : _GEN_1548; // @[executor.scala 466:52]
  wire [7:0] _GEN_1807 = opcode_1 == 4'hf ? _GEN_781 : _GEN_1549; // @[executor.scala 466:52]
  wire [7:0] _GEN_1808 = opcode_1 == 4'hf ? _GEN_782 : _GEN_1550; // @[executor.scala 466:52]
  wire [7:0] _GEN_1809 = opcode_1 == 4'hf ? _GEN_783 : _GEN_1551; // @[executor.scala 466:52]
  wire [7:0] _GEN_1810 = opcode_1 == 4'hf ? _GEN_784 : _GEN_1552; // @[executor.scala 466:52]
  wire [7:0] _GEN_1811 = opcode_1 == 4'hf ? _GEN_785 : _GEN_1553; // @[executor.scala 466:52]
  wire [7:0] _GEN_1812 = opcode_1 == 4'hf ? _GEN_786 : _GEN_1554; // @[executor.scala 466:52]
  wire [7:0] _GEN_1813 = opcode_1 == 4'hf ? _GEN_787 : _GEN_1555; // @[executor.scala 466:52]
  wire [7:0] _GEN_1814 = opcode_1 == 4'hf ? _GEN_788 : _GEN_1556; // @[executor.scala 466:52]
  wire [7:0] _GEN_1815 = opcode_1 == 4'hf ? _GEN_789 : _GEN_1557; // @[executor.scala 466:52]
  wire [7:0] _GEN_1816 = opcode_1 == 4'hf ? _GEN_790 : _GEN_1558; // @[executor.scala 466:52]
  wire [7:0] _GEN_1817 = opcode_1 == 4'hf ? _GEN_791 : _GEN_1559; // @[executor.scala 466:52]
  wire [7:0] _GEN_1818 = opcode_1 == 4'hf ? _GEN_792 : _GEN_1560; // @[executor.scala 466:52]
  wire [7:0] _GEN_1819 = opcode_1 == 4'hf ? _GEN_793 : _GEN_1561; // @[executor.scala 466:52]
  wire [7:0] _GEN_1820 = opcode_1 == 4'hf ? _GEN_794 : _GEN_1562; // @[executor.scala 466:52]
  wire [7:0] _GEN_1821 = opcode_1 == 4'hf ? _GEN_795 : _GEN_1563; // @[executor.scala 466:52]
  wire [7:0] _GEN_1822 = opcode_1 == 4'hf ? _GEN_796 : _GEN_1564; // @[executor.scala 466:52]
  wire [7:0] _GEN_1823 = opcode_1 == 4'hf ? _GEN_797 : _GEN_1565; // @[executor.scala 466:52]
  wire [7:0] _GEN_1824 = opcode_1 == 4'hf ? _GEN_798 : _GEN_1566; // @[executor.scala 466:52]
  wire [7:0] _GEN_1825 = opcode_1 == 4'hf ? _GEN_799 : _GEN_1567; // @[executor.scala 466:52]
  wire [7:0] _GEN_1826 = opcode_1 == 4'hf ? _GEN_800 : _GEN_1568; // @[executor.scala 466:52]
  wire [7:0] _GEN_1827 = opcode_1 == 4'hf ? _GEN_801 : _GEN_1569; // @[executor.scala 466:52]
  wire [7:0] _GEN_1828 = opcode_1 == 4'hf ? _GEN_802 : _GEN_1570; // @[executor.scala 466:52]
  wire [7:0] _GEN_1829 = opcode_1 == 4'hf ? _GEN_803 : _GEN_1571; // @[executor.scala 466:52]
  wire [7:0] _GEN_1830 = opcode_1 == 4'hf ? _GEN_804 : _GEN_1572; // @[executor.scala 466:52]
  wire [7:0] _GEN_1831 = opcode_1 == 4'hf ? _GEN_805 : _GEN_1573; // @[executor.scala 466:52]
  wire [7:0] _GEN_1832 = opcode_1 == 4'hf ? _GEN_806 : _GEN_1574; // @[executor.scala 466:52]
  wire [7:0] _GEN_1833 = opcode_1 == 4'hf ? _GEN_807 : _GEN_1575; // @[executor.scala 466:52]
  wire [7:0] _GEN_1834 = opcode_1 == 4'hf ? _GEN_808 : _GEN_1576; // @[executor.scala 466:52]
  wire [7:0] _GEN_1835 = opcode_1 == 4'hf ? _GEN_809 : _GEN_1577; // @[executor.scala 466:52]
  wire [7:0] _GEN_1836 = opcode_1 == 4'hf ? _GEN_810 : _GEN_1578; // @[executor.scala 466:52]
  wire [7:0] _GEN_1837 = opcode_1 == 4'hf ? _GEN_811 : _GEN_1579; // @[executor.scala 466:52]
  wire [7:0] _GEN_1838 = opcode_1 == 4'hf ? _GEN_812 : _GEN_1580; // @[executor.scala 466:52]
  wire [7:0] _GEN_1839 = opcode_1 == 4'hf ? _GEN_813 : _GEN_1581; // @[executor.scala 466:52]
  wire [7:0] _GEN_1840 = opcode_1 == 4'hf ? _GEN_814 : _GEN_1582; // @[executor.scala 466:52]
  wire [7:0] _GEN_1841 = opcode_1 == 4'hf ? _GEN_815 : _GEN_1583; // @[executor.scala 466:52]
  wire [7:0] _GEN_1842 = opcode_1 == 4'hf ? _GEN_816 : _GEN_1584; // @[executor.scala 466:52]
  wire [7:0] _GEN_1843 = opcode_1 == 4'hf ? _GEN_817 : _GEN_1585; // @[executor.scala 466:52]
  wire [7:0] _GEN_1844 = opcode_1 == 4'hf ? _GEN_818 : _GEN_1586; // @[executor.scala 466:52]
  wire [7:0] _GEN_1845 = opcode_1 == 4'hf ? _GEN_819 : _GEN_1587; // @[executor.scala 466:52]
  wire [7:0] _GEN_1846 = opcode_1 == 4'hf ? _GEN_820 : _GEN_1588; // @[executor.scala 466:52]
  wire [7:0] _GEN_1847 = opcode_1 == 4'hf ? _GEN_821 : _GEN_1589; // @[executor.scala 466:52]
  wire [7:0] _GEN_1848 = opcode_1 == 4'hf ? _GEN_822 : _GEN_1590; // @[executor.scala 466:52]
  wire [7:0] _GEN_1849 = opcode_1 == 4'hf ? _GEN_823 : _GEN_1591; // @[executor.scala 466:52]
  wire [7:0] _GEN_1850 = opcode_1 == 4'hf ? _GEN_824 : _GEN_1592; // @[executor.scala 466:52]
  wire [7:0] _GEN_1851 = opcode_1 == 4'hf ? _GEN_825 : _GEN_1593; // @[executor.scala 466:52]
  wire [7:0] _GEN_1852 = opcode_1 == 4'hf ? _GEN_826 : _GEN_1594; // @[executor.scala 466:52]
  wire [7:0] _GEN_1853 = opcode_1 == 4'hf ? _GEN_827 : _GEN_1595; // @[executor.scala 466:52]
  wire [7:0] _GEN_1854 = opcode_1 == 4'hf ? _GEN_828 : _GEN_1596; // @[executor.scala 466:52]
  wire [7:0] _GEN_1855 = opcode_1 == 4'hf ? _GEN_829 : _GEN_1597; // @[executor.scala 466:52]
  wire [7:0] _GEN_1856 = opcode_1 == 4'hf ? _GEN_830 : _GEN_1598; // @[executor.scala 466:52]
  wire [7:0] _GEN_1857 = opcode_1 == 4'hf ? _GEN_831 : _GEN_1599; // @[executor.scala 466:52]
  wire [7:0] _GEN_1858 = opcode_1 == 4'hf ? _GEN_832 : _GEN_1600; // @[executor.scala 466:52]
  wire [7:0] _GEN_1859 = opcode_1 == 4'hf ? _GEN_833 : _GEN_1601; // @[executor.scala 466:52]
  wire [7:0] _GEN_1860 = opcode_1 == 4'hf ? _GEN_834 : _GEN_1602; // @[executor.scala 466:52]
  wire [7:0] _GEN_1861 = opcode_1 == 4'hf ? _GEN_835 : _GEN_1603; // @[executor.scala 466:52]
  wire [7:0] _GEN_1862 = opcode_1 == 4'hf ? _GEN_836 : _GEN_1604; // @[executor.scala 466:52]
  wire [7:0] _GEN_1863 = opcode_1 == 4'hf ? _GEN_837 : _GEN_1605; // @[executor.scala 466:52]
  wire [7:0] _GEN_1864 = opcode_1 == 4'hf ? _GEN_838 : _GEN_1606; // @[executor.scala 466:52]
  wire [7:0] _GEN_1865 = opcode_1 == 4'hf ? _GEN_839 : _GEN_1607; // @[executor.scala 466:52]
  wire [7:0] _GEN_1866 = opcode_1 == 4'hf ? _GEN_840 : _GEN_1608; // @[executor.scala 466:52]
  wire [7:0] _GEN_1867 = opcode_1 == 4'hf ? _GEN_841 : _GEN_1609; // @[executor.scala 466:52]
  wire [7:0] _GEN_1868 = opcode_1 == 4'hf ? _GEN_842 : _GEN_1610; // @[executor.scala 466:52]
  wire [7:0] _GEN_1869 = opcode_1 == 4'hf ? _GEN_843 : _GEN_1611; // @[executor.scala 466:52]
  wire [7:0] _GEN_1870 = opcode_1 == 4'hf ? _GEN_844 : _GEN_1612; // @[executor.scala 466:52]
  wire [7:0] _GEN_1871 = opcode_1 == 4'hf ? _GEN_845 : _GEN_1613; // @[executor.scala 466:52]
  wire [7:0] _GEN_1872 = opcode_1 == 4'hf ? _GEN_846 : _GEN_1614; // @[executor.scala 466:52]
  wire [7:0] _GEN_1873 = opcode_1 == 4'hf ? _GEN_847 : _GEN_1615; // @[executor.scala 466:52]
  wire [7:0] _GEN_1874 = opcode_1 == 4'hf ? _GEN_848 : _GEN_1616; // @[executor.scala 466:52]
  wire [7:0] _GEN_1875 = opcode_1 == 4'hf ? _GEN_849 : _GEN_1617; // @[executor.scala 466:52]
  wire [7:0] _GEN_1876 = opcode_1 == 4'hf ? _GEN_850 : _GEN_1618; // @[executor.scala 466:52]
  wire [7:0] _GEN_1877 = opcode_1 == 4'hf ? _GEN_851 : _GEN_1619; // @[executor.scala 466:52]
  wire [7:0] _GEN_1878 = opcode_1 == 4'hf ? _GEN_852 : _GEN_1620; // @[executor.scala 466:52]
  wire [7:0] _GEN_1879 = opcode_1 == 4'hf ? _GEN_853 : _GEN_1621; // @[executor.scala 466:52]
  wire [7:0] _GEN_1880 = opcode_1 == 4'hf ? _GEN_854 : _GEN_1622; // @[executor.scala 466:52]
  wire [7:0] _GEN_1881 = opcode_1 == 4'hf ? _GEN_855 : _GEN_1623; // @[executor.scala 466:52]
  wire [7:0] _GEN_1882 = opcode_1 == 4'hf ? _GEN_856 : _GEN_1624; // @[executor.scala 466:52]
  wire [7:0] _GEN_1883 = opcode_1 == 4'hf ? _GEN_857 : _GEN_1625; // @[executor.scala 466:52]
  wire [7:0] _GEN_1884 = opcode_1 == 4'hf ? _GEN_858 : _GEN_1626; // @[executor.scala 466:52]
  wire [7:0] _GEN_1885 = opcode_1 == 4'hf ? _GEN_859 : _GEN_1627; // @[executor.scala 466:52]
  wire [7:0] _GEN_1886 = opcode_1 == 4'hf ? _GEN_860 : _GEN_1628; // @[executor.scala 466:52]
  wire [7:0] _GEN_1887 = opcode_1 == 4'hf ? _GEN_861 : _GEN_1629; // @[executor.scala 466:52]
  wire [7:0] _GEN_1888 = opcode_1 == 4'hf ? _GEN_862 : _GEN_1630; // @[executor.scala 466:52]
  wire [7:0] _GEN_1889 = opcode_1 == 4'hf ? _GEN_863 : _GEN_1631; // @[executor.scala 466:52]
  wire [7:0] _GEN_1890 = opcode_1 == 4'hf ? _GEN_864 : _GEN_1632; // @[executor.scala 466:52]
  wire [7:0] _GEN_1891 = opcode_1 == 4'hf ? _GEN_865 : _GEN_1633; // @[executor.scala 466:52]
  wire [7:0] _GEN_1892 = opcode_1 == 4'hf ? _GEN_866 : _GEN_1634; // @[executor.scala 466:52]
  wire [7:0] _GEN_1893 = opcode_1 == 4'hf ? _GEN_867 : _GEN_1635; // @[executor.scala 466:52]
  wire [7:0] _GEN_1894 = opcode_1 == 4'hf ? _GEN_868 : _GEN_1636; // @[executor.scala 466:52]
  wire [7:0] _GEN_1895 = opcode_1 == 4'hf ? _GEN_869 : _GEN_1637; // @[executor.scala 466:52]
  wire [7:0] _GEN_1896 = opcode_1 == 4'hf ? _GEN_870 : _GEN_1638; // @[executor.scala 466:52]
  wire [7:0] _GEN_1897 = opcode_1 == 4'hf ? _GEN_871 : _GEN_1639; // @[executor.scala 466:52]
  wire [7:0] _GEN_1898 = opcode_1 == 4'hf ? _GEN_872 : _GEN_1640; // @[executor.scala 466:52]
  wire [7:0] _GEN_1899 = opcode_1 == 4'hf ? _GEN_873 : _GEN_1641; // @[executor.scala 466:52]
  wire [7:0] _GEN_1900 = opcode_1 == 4'hf ? _GEN_874 : _GEN_1642; // @[executor.scala 466:52]
  wire [7:0] _GEN_1901 = opcode_1 == 4'hf ? _GEN_875 : _GEN_1643; // @[executor.scala 466:52]
  wire [7:0] _GEN_1902 = opcode_1 == 4'hf ? _GEN_876 : _GEN_1644; // @[executor.scala 466:52]
  wire [7:0] _GEN_1903 = opcode_1 == 4'hf ? _GEN_877 : _GEN_1645; // @[executor.scala 466:52]
  wire [7:0] _GEN_1904 = opcode_1 == 4'hf ? _GEN_878 : _GEN_1646; // @[executor.scala 466:52]
  wire [7:0] _GEN_1905 = opcode_1 == 4'hf ? _GEN_879 : _GEN_1647; // @[executor.scala 466:52]
  wire [7:0] _GEN_1906 = opcode_1 == 4'hf ? _GEN_880 : _GEN_1648; // @[executor.scala 466:52]
  wire [7:0] _GEN_1907 = opcode_1 == 4'hf ? _GEN_881 : _GEN_1649; // @[executor.scala 466:52]
  wire [7:0] _GEN_1908 = opcode_1 == 4'hf ? _GEN_882 : _GEN_1650; // @[executor.scala 466:52]
  wire [7:0] _GEN_1909 = opcode_1 == 4'hf ? _GEN_883 : _GEN_1651; // @[executor.scala 466:52]
  wire [7:0] _GEN_1910 = opcode_1 == 4'hf ? _GEN_884 : _GEN_1652; // @[executor.scala 466:52]
  wire [7:0] _GEN_1911 = opcode_1 == 4'hf ? _GEN_885 : _GEN_1653; // @[executor.scala 466:52]
  wire [7:0] _GEN_1912 = opcode_1 == 4'hf ? _GEN_886 : _GEN_1654; // @[executor.scala 466:52]
  wire [7:0] _GEN_1913 = opcode_1 == 4'hf ? _GEN_887 : _GEN_1655; // @[executor.scala 466:52]
  wire [7:0] _GEN_1914 = opcode_1 == 4'hf ? _GEN_888 : _GEN_1656; // @[executor.scala 466:52]
  wire [7:0] _GEN_1915 = opcode_1 == 4'hf ? _GEN_889 : _GEN_1657; // @[executor.scala 466:52]
  wire [7:0] _GEN_1916 = opcode_1 == 4'hf ? _GEN_890 : _GEN_1658; // @[executor.scala 466:52]
  wire [7:0] _GEN_1917 = opcode_1 == 4'hf ? _GEN_891 : _GEN_1659; // @[executor.scala 466:52]
  wire [7:0] _GEN_1918 = opcode_1 == 4'hf ? _GEN_892 : _GEN_1660; // @[executor.scala 466:52]
  wire [7:0] _GEN_1919 = opcode_1 == 4'hf ? _GEN_893 : _GEN_1661; // @[executor.scala 466:52]
  wire [7:0] _GEN_1920 = opcode_1 == 4'hf ? _GEN_894 : _GEN_1662; // @[executor.scala 466:52]
  wire [7:0] _GEN_1921 = opcode_1 == 4'hf ? _GEN_895 : _GEN_1663; // @[executor.scala 466:52]
  wire [7:0] _GEN_1922 = opcode_1 == 4'hf ? _GEN_896 : _GEN_1664; // @[executor.scala 466:52]
  wire [7:0] _GEN_1923 = opcode_1 == 4'hf ? _GEN_897 : _GEN_1665; // @[executor.scala 466:52]
  wire [7:0] _GEN_1924 = opcode_1 == 4'hf ? _GEN_898 : _GEN_1666; // @[executor.scala 466:52]
  wire [7:0] _GEN_1925 = opcode_1 == 4'hf ? _GEN_899 : _GEN_1667; // @[executor.scala 466:52]
  wire [7:0] _GEN_1926 = opcode_1 == 4'hf ? _GEN_900 : _GEN_1668; // @[executor.scala 466:52]
  wire [7:0] _GEN_1927 = opcode_1 == 4'hf ? _GEN_901 : _GEN_1669; // @[executor.scala 466:52]
  wire [7:0] _GEN_1928 = opcode_1 == 4'hf ? _GEN_902 : _GEN_1670; // @[executor.scala 466:52]
  wire [7:0] _GEN_1929 = opcode_1 == 4'hf ? _GEN_903 : _GEN_1671; // @[executor.scala 466:52]
  wire [7:0] _GEN_1930 = opcode_1 == 4'hf ? _GEN_904 : _GEN_1672; // @[executor.scala 466:52]
  wire [7:0] _GEN_1931 = opcode_1 == 4'hf ? _GEN_905 : _GEN_1673; // @[executor.scala 466:52]
  wire [7:0] _GEN_1932 = opcode_1 == 4'hf ? _GEN_906 : _GEN_1674; // @[executor.scala 466:52]
  wire [7:0] _GEN_1933 = opcode_1 == 4'hf ? _GEN_907 : _GEN_1675; // @[executor.scala 466:52]
  wire [7:0] _GEN_1934 = opcode_1 == 4'hf ? _GEN_908 : _GEN_1676; // @[executor.scala 466:52]
  wire [7:0] _GEN_1935 = opcode_1 == 4'hf ? _GEN_909 : _GEN_1677; // @[executor.scala 466:52]
  wire [7:0] _GEN_1936 = opcode_1 == 4'hf ? _GEN_910 : _GEN_1678; // @[executor.scala 466:52]
  wire [7:0] _GEN_1937 = opcode_1 == 4'hf ? _GEN_911 : _GEN_1679; // @[executor.scala 466:52]
  wire [7:0] _GEN_1938 = opcode_1 == 4'hf ? _GEN_912 : _GEN_1680; // @[executor.scala 466:52]
  wire [7:0] _GEN_1939 = opcode_1 == 4'hf ? _GEN_913 : _GEN_1681; // @[executor.scala 466:52]
  wire [7:0] _GEN_1940 = opcode_1 == 4'hf ? _GEN_914 : _GEN_1682; // @[executor.scala 466:52]
  wire [7:0] _GEN_1941 = opcode_1 == 4'hf ? _GEN_915 : _GEN_1683; // @[executor.scala 466:52]
  wire [7:0] _GEN_1942 = opcode_1 == 4'hf ? _GEN_916 : _GEN_1684; // @[executor.scala 466:52]
  wire [7:0] _GEN_1943 = opcode_1 == 4'hf ? _GEN_917 : _GEN_1685; // @[executor.scala 466:52]
  wire [7:0] _GEN_1944 = opcode_1 == 4'hf ? _GEN_918 : _GEN_1686; // @[executor.scala 466:52]
  wire [7:0] _GEN_1945 = opcode_1 == 4'hf ? _GEN_919 : _GEN_1687; // @[executor.scala 466:52]
  wire [7:0] _GEN_1946 = opcode_1 == 4'hf ? _GEN_920 : _GEN_1688; // @[executor.scala 466:52]
  wire [7:0] _GEN_1947 = opcode_1 == 4'hf ? _GEN_921 : _GEN_1689; // @[executor.scala 466:52]
  wire [7:0] _GEN_1948 = opcode_1 == 4'hf ? _GEN_922 : _GEN_1690; // @[executor.scala 466:52]
  wire [7:0] _GEN_1949 = opcode_1 == 4'hf ? _GEN_923 : _GEN_1691; // @[executor.scala 466:52]
  wire [7:0] _GEN_1950 = opcode_1 == 4'hf ? _GEN_924 : _GEN_1692; // @[executor.scala 466:52]
  wire [7:0] _GEN_1951 = opcode_1 == 4'hf ? _GEN_925 : _GEN_1693; // @[executor.scala 466:52]
  wire [7:0] _GEN_1952 = opcode_1 == 4'hf ? _GEN_926 : _GEN_1694; // @[executor.scala 466:52]
  wire [7:0] _GEN_1953 = opcode_1 == 4'hf ? _GEN_927 : _GEN_1695; // @[executor.scala 466:52]
  wire [7:0] _GEN_1954 = opcode_1 == 4'hf ? _GEN_928 : _GEN_1696; // @[executor.scala 466:52]
  wire [7:0] _GEN_1955 = opcode_1 == 4'hf ? _GEN_929 : _GEN_1697; // @[executor.scala 466:52]
  wire [7:0] _GEN_1956 = opcode_1 == 4'hf ? _GEN_930 : _GEN_1698; // @[executor.scala 466:52]
  wire [7:0] _GEN_1957 = opcode_1 == 4'hf ? _GEN_931 : _GEN_1699; // @[executor.scala 466:52]
  wire [7:0] _GEN_1958 = opcode_1 == 4'hf ? _GEN_932 : _GEN_1700; // @[executor.scala 466:52]
  wire [7:0] _GEN_1959 = opcode_1 == 4'hf ? _GEN_933 : _GEN_1701; // @[executor.scala 466:52]
  wire [7:0] _GEN_1960 = opcode_1 == 4'hf ? _GEN_934 : _GEN_1702; // @[executor.scala 466:52]
  wire [7:0] _GEN_1961 = opcode_1 == 4'hf ? _GEN_935 : _GEN_1703; // @[executor.scala 466:52]
  wire [7:0] _GEN_1962 = opcode_1 == 4'hf ? _GEN_936 : _GEN_1704; // @[executor.scala 466:52]
  wire [7:0] _GEN_1963 = opcode_1 == 4'hf ? _GEN_937 : _GEN_1705; // @[executor.scala 466:52]
  wire [7:0] _GEN_1964 = opcode_1 == 4'hf ? _GEN_938 : _GEN_1706; // @[executor.scala 466:52]
  wire [7:0] _GEN_1965 = opcode_1 == 4'hf ? _GEN_939 : _GEN_1707; // @[executor.scala 466:52]
  wire [7:0] _GEN_1966 = opcode_1 == 4'hf ? _GEN_940 : _GEN_1708; // @[executor.scala 466:52]
  wire [7:0] _GEN_1967 = opcode_1 == 4'hf ? _GEN_941 : _GEN_1709; // @[executor.scala 466:52]
  wire [7:0] _GEN_1968 = opcode_1 == 4'hf ? _GEN_942 : _GEN_1710; // @[executor.scala 466:52]
  wire [7:0] _GEN_1969 = opcode_1 == 4'hf ? _GEN_943 : _GEN_1711; // @[executor.scala 466:52]
  wire [7:0] _GEN_1970 = opcode_1 == 4'hf ? _GEN_944 : _GEN_1712; // @[executor.scala 466:52]
  wire [7:0] _GEN_1971 = opcode_1 == 4'hf ? _GEN_945 : _GEN_1713; // @[executor.scala 466:52]
  wire [7:0] _GEN_1972 = opcode_1 == 4'hf ? _GEN_946 : _GEN_1714; // @[executor.scala 466:52]
  wire [7:0] _GEN_1973 = opcode_1 == 4'hf ? _GEN_947 : _GEN_1715; // @[executor.scala 466:52]
  wire [7:0] _GEN_1974 = opcode_1 == 4'hf ? _GEN_948 : _GEN_1716; // @[executor.scala 466:52]
  wire [7:0] _GEN_1975 = opcode_1 == 4'hf ? _GEN_949 : _GEN_1717; // @[executor.scala 466:52]
  wire [7:0] _GEN_1976 = opcode_1 == 4'hf ? _GEN_950 : _GEN_1718; // @[executor.scala 466:52]
  wire [7:0] _GEN_1977 = opcode_1 == 4'hf ? _GEN_951 : _GEN_1719; // @[executor.scala 466:52]
  wire [7:0] _GEN_1978 = opcode_1 == 4'hf ? _GEN_952 : _GEN_1720; // @[executor.scala 466:52]
  wire [7:0] _GEN_1979 = opcode_1 == 4'hf ? _GEN_953 : _GEN_1721; // @[executor.scala 466:52]
  wire [7:0] _GEN_1980 = opcode_1 == 4'hf ? _GEN_954 : _GEN_1722; // @[executor.scala 466:52]
  wire [7:0] _GEN_1981 = opcode_1 == 4'hf ? _GEN_955 : _GEN_1723; // @[executor.scala 466:52]
  wire [7:0] _GEN_1982 = opcode_1 == 4'hf ? _GEN_956 : _GEN_1724; // @[executor.scala 466:52]
  wire [7:0] _GEN_1983 = opcode_1 == 4'hf ? _GEN_957 : _GEN_1725; // @[executor.scala 466:52]
  wire [7:0] _GEN_1984 = opcode_1 == 4'hf ? _GEN_958 : _GEN_1726; // @[executor.scala 466:52]
  wire [7:0] _GEN_1985 = opcode_1 == 4'hf ? _GEN_959 : _GEN_1727; // @[executor.scala 466:52]
  wire [7:0] _GEN_1986 = opcode_1 == 4'hf ? _GEN_960 : _GEN_1728; // @[executor.scala 466:52]
  wire [7:0] _GEN_1987 = opcode_1 == 4'hf ? _GEN_961 : _GEN_1729; // @[executor.scala 466:52]
  wire [7:0] _GEN_1988 = opcode_1 == 4'hf ? _GEN_962 : _GEN_1730; // @[executor.scala 466:52]
  wire [7:0] _GEN_1989 = opcode_1 == 4'hf ? _GEN_963 : _GEN_1731; // @[executor.scala 466:52]
  wire [7:0] _GEN_1990 = opcode_1 == 4'hf ? _GEN_964 : _GEN_1732; // @[executor.scala 466:52]
  wire [7:0] _GEN_1991 = opcode_1 == 4'hf ? _GEN_965 : _GEN_1733; // @[executor.scala 466:52]
  wire [7:0] _GEN_1992 = opcode_1 == 4'hf ? _GEN_966 : _GEN_1734; // @[executor.scala 466:52]
  wire [7:0] _GEN_1993 = opcode_1 == 4'hf ? _GEN_967 : _GEN_1735; // @[executor.scala 466:52]
  wire [7:0] _GEN_1994 = opcode_1 == 4'hf ? _GEN_968 : _GEN_1736; // @[executor.scala 466:52]
  wire [7:0] _GEN_1995 = opcode_1 == 4'hf ? _GEN_969 : _GEN_1737; // @[executor.scala 466:52]
  wire [7:0] _GEN_1996 = opcode_1 == 4'hf ? _GEN_970 : _GEN_1738; // @[executor.scala 466:52]
  wire [7:0] _GEN_1997 = opcode_1 == 4'hf ? _GEN_971 : _GEN_1739; // @[executor.scala 466:52]
  wire [7:0] _GEN_1998 = opcode_1 == 4'hf ? _GEN_972 : _GEN_1740; // @[executor.scala 466:52]
  wire [7:0] _GEN_1999 = opcode_1 == 4'hf ? _GEN_973 : _GEN_1741; // @[executor.scala 466:52]
  wire [7:0] _GEN_2000 = opcode_1 == 4'hf ? _GEN_974 : _GEN_1742; // @[executor.scala 466:52]
  wire [7:0] _GEN_2001 = opcode_1 == 4'hf ? _GEN_975 : _GEN_1743; // @[executor.scala 466:52]
  wire [7:0] _GEN_2002 = opcode_1 == 4'hf ? _GEN_976 : _GEN_1744; // @[executor.scala 466:52]
  wire [7:0] _GEN_2003 = opcode_1 == 4'hf ? _GEN_977 : _GEN_1745; // @[executor.scala 466:52]
  wire [7:0] _GEN_2004 = opcode_1 == 4'hf ? _GEN_978 : _GEN_1746; // @[executor.scala 466:52]
  wire [7:0] _GEN_2005 = opcode_1 == 4'hf ? _GEN_979 : _GEN_1747; // @[executor.scala 466:52]
  wire [7:0] _GEN_2006 = opcode_1 == 4'hf ? _GEN_980 : _GEN_1748; // @[executor.scala 466:52]
  wire [7:0] _GEN_2007 = opcode_1 == 4'hf ? _GEN_981 : _GEN_1749; // @[executor.scala 466:52]
  wire [7:0] _GEN_2008 = opcode_1 == 4'hf ? _GEN_982 : _GEN_1750; // @[executor.scala 466:52]
  wire [7:0] _GEN_2009 = opcode_1 == 4'hf ? _GEN_983 : _GEN_1751; // @[executor.scala 466:52]
  wire [7:0] _GEN_2010 = opcode_1 == 4'hf ? _GEN_984 : _GEN_1752; // @[executor.scala 466:52]
  wire [7:0] _GEN_2011 = opcode_1 == 4'hf ? _GEN_985 : _GEN_1753; // @[executor.scala 466:52]
  wire [7:0] _GEN_2012 = opcode_1 == 4'hf ? _GEN_986 : _GEN_1754; // @[executor.scala 466:52]
  wire [7:0] _GEN_2013 = opcode_1 == 4'hf ? _GEN_987 : _GEN_1755; // @[executor.scala 466:52]
  wire [7:0] _GEN_2014 = opcode_1 == 4'hf ? _GEN_988 : _GEN_1756; // @[executor.scala 466:52]
  wire [7:0] _GEN_2015 = opcode_1 == 4'hf ? _GEN_989 : _GEN_1757; // @[executor.scala 466:52]
  wire [7:0] _GEN_2016 = opcode_1 == 4'hf ? _GEN_990 : _GEN_1758; // @[executor.scala 466:52]
  wire [7:0] _GEN_2017 = opcode_1 == 4'hf ? _GEN_991 : _GEN_1759; // @[executor.scala 466:52]
  wire [7:0] _GEN_2018 = opcode_1 == 4'hf ? _GEN_992 : _GEN_1760; // @[executor.scala 466:52]
  wire [7:0] _GEN_2019 = opcode_1 == 4'hf ? _GEN_993 : _GEN_1761; // @[executor.scala 466:52]
  wire [7:0] _GEN_2020 = opcode_1 == 4'hf ? _GEN_994 : _GEN_1762; // @[executor.scala 466:52]
  wire [7:0] _GEN_2021 = opcode_1 == 4'hf ? _GEN_995 : _GEN_1763; // @[executor.scala 466:52]
  wire [7:0] _GEN_2022 = opcode_1 == 4'hf ? _GEN_996 : _GEN_1764; // @[executor.scala 466:52]
  wire [7:0] _GEN_2023 = opcode_1 == 4'hf ? _GEN_997 : _GEN_1765; // @[executor.scala 466:52]
  wire [7:0] _GEN_2024 = opcode_1 == 4'hf ? _GEN_998 : _GEN_1766; // @[executor.scala 466:52]
  wire [7:0] _GEN_2025 = opcode_1 == 4'hf ? _GEN_999 : _GEN_1767; // @[executor.scala 466:52]
  wire [7:0] _GEN_2026 = opcode_1 == 4'hf ? _GEN_1000 : _GEN_1768; // @[executor.scala 466:52]
  wire [7:0] _GEN_2027 = opcode_1 == 4'hf ? _GEN_1001 : _GEN_1769; // @[executor.scala 466:52]
  wire [7:0] _GEN_2028 = opcode_1 == 4'hf ? _GEN_1002 : _GEN_1770; // @[executor.scala 466:52]
  wire [7:0] _GEN_2029 = opcode_1 == 4'hf ? _GEN_1003 : _GEN_1771; // @[executor.scala 466:52]
  wire [7:0] _GEN_2030 = opcode_1 == 4'hf ? _GEN_1004 : _GEN_1772; // @[executor.scala 466:52]
  wire [7:0] _GEN_2031 = opcode_1 == 4'hf ? _GEN_1005 : _GEN_1773; // @[executor.scala 466:52]
  wire [7:0] _GEN_2032 = opcode_1 == 4'hf ? _GEN_1006 : _GEN_1774; // @[executor.scala 466:52]
  wire [7:0] _GEN_2033 = opcode_1 == 4'hf ? _GEN_1007 : _GEN_1775; // @[executor.scala 466:52]
  wire [7:0] _GEN_2034 = opcode_1 == 4'hf ? _GEN_1008 : _GEN_1776; // @[executor.scala 466:52]
  wire [7:0] _GEN_2035 = opcode_1 == 4'hf ? _GEN_1009 : _GEN_1777; // @[executor.scala 466:52]
  wire [7:0] _GEN_2036 = opcode_1 == 4'hf ? _GEN_1010 : _GEN_1778; // @[executor.scala 466:52]
  wire [7:0] _GEN_2037 = opcode_1 == 4'hf ? _GEN_1011 : _GEN_1779; // @[executor.scala 466:52]
  wire [7:0] _GEN_2038 = opcode_1 == 4'hf ? _GEN_1012 : _GEN_1780; // @[executor.scala 466:52]
  wire [7:0] _GEN_2039 = opcode_1 == 4'hf ? _GEN_1013 : _GEN_1781; // @[executor.scala 466:52]
  wire [7:0] _GEN_2040 = opcode_1 == 4'hf ? _GEN_1014 : _GEN_1782; // @[executor.scala 466:52]
  wire [7:0] _GEN_2041 = opcode_1 == 4'hf ? _GEN_1015 : _GEN_1783; // @[executor.scala 466:52]
  wire [7:0] _GEN_2042 = opcode_1 == 4'hf ? _GEN_1016 : _GEN_1784; // @[executor.scala 466:52]
  wire [7:0] _GEN_2043 = opcode_1 == 4'hf ? _GEN_1017 : _GEN_1785; // @[executor.scala 466:52]
  wire [7:0] _GEN_2044 = opcode_1 == 4'hf ? _GEN_1018 : _GEN_1786; // @[executor.scala 466:52]
  wire [7:0] _GEN_2045 = opcode_1 == 4'hf ? _GEN_1019 : _GEN_1787; // @[executor.scala 466:52]
  wire [7:0] _GEN_2046 = opcode_1 == 4'hf ? _GEN_1020 : _GEN_1788; // @[executor.scala 466:52]
  wire [7:0] _GEN_2047 = opcode_1 == 4'hf ? _GEN_1021 : _GEN_1789; // @[executor.scala 466:52]
  wire [7:0] _GEN_2048 = opcode_1 == 4'hf ? _GEN_1022 : _GEN_1790; // @[executor.scala 466:52]
  wire [7:0] _GEN_2049 = opcode_1 == 4'hf ? _GEN_1023 : _GEN_1791; // @[executor.scala 466:52]
  wire [7:0] _GEN_2050 = opcode_1 == 4'hf ? _GEN_1024 : _GEN_1792; // @[executor.scala 466:52]
  wire [7:0] _GEN_2051 = opcode_1 == 4'hf ? _GEN_1025 : _GEN_1793; // @[executor.scala 466:52]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_2 = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8594 = {{2'd0}, dst_offset_2}; // @[executor.scala 473:49]
  wire [7:0] byte_512 = field_2[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2052 = mask_2[0] ? byte_512 : _GEN_1796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_513 = field_2[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2053 = mask_2[1] ? byte_513 : _GEN_1797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_514 = field_2[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2054 = mask_2[2] ? byte_514 : _GEN_1798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_515 = field_2[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2055 = mask_2[3] ? byte_515 : _GEN_1799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2056 = _GEN_8594 == 8'h0 ? _GEN_2052 : _GEN_1796; // @[executor.scala 473:84]
  wire [7:0] _GEN_2057 = _GEN_8594 == 8'h0 ? _GEN_2053 : _GEN_1797; // @[executor.scala 473:84]
  wire [7:0] _GEN_2058 = _GEN_8594 == 8'h0 ? _GEN_2054 : _GEN_1798; // @[executor.scala 473:84]
  wire [7:0] _GEN_2059 = _GEN_8594 == 8'h0 ? _GEN_2055 : _GEN_1799; // @[executor.scala 473:84]
  wire [7:0] _GEN_2060 = mask_2[0] ? byte_512 : _GEN_1800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2061 = mask_2[1] ? byte_513 : _GEN_1801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2062 = mask_2[2] ? byte_514 : _GEN_1802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2063 = mask_2[3] ? byte_515 : _GEN_1803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2064 = _GEN_8594 == 8'h1 ? _GEN_2060 : _GEN_1800; // @[executor.scala 473:84]
  wire [7:0] _GEN_2065 = _GEN_8594 == 8'h1 ? _GEN_2061 : _GEN_1801; // @[executor.scala 473:84]
  wire [7:0] _GEN_2066 = _GEN_8594 == 8'h1 ? _GEN_2062 : _GEN_1802; // @[executor.scala 473:84]
  wire [7:0] _GEN_2067 = _GEN_8594 == 8'h1 ? _GEN_2063 : _GEN_1803; // @[executor.scala 473:84]
  wire [7:0] _GEN_2068 = mask_2[0] ? byte_512 : _GEN_1804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2069 = mask_2[1] ? byte_513 : _GEN_1805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2070 = mask_2[2] ? byte_514 : _GEN_1806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2071 = mask_2[3] ? byte_515 : _GEN_1807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2072 = _GEN_8594 == 8'h2 ? _GEN_2068 : _GEN_1804; // @[executor.scala 473:84]
  wire [7:0] _GEN_2073 = _GEN_8594 == 8'h2 ? _GEN_2069 : _GEN_1805; // @[executor.scala 473:84]
  wire [7:0] _GEN_2074 = _GEN_8594 == 8'h2 ? _GEN_2070 : _GEN_1806; // @[executor.scala 473:84]
  wire [7:0] _GEN_2075 = _GEN_8594 == 8'h2 ? _GEN_2071 : _GEN_1807; // @[executor.scala 473:84]
  wire [7:0] _GEN_2076 = mask_2[0] ? byte_512 : _GEN_1808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2077 = mask_2[1] ? byte_513 : _GEN_1809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2078 = mask_2[2] ? byte_514 : _GEN_1810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2079 = mask_2[3] ? byte_515 : _GEN_1811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2080 = _GEN_8594 == 8'h3 ? _GEN_2076 : _GEN_1808; // @[executor.scala 473:84]
  wire [7:0] _GEN_2081 = _GEN_8594 == 8'h3 ? _GEN_2077 : _GEN_1809; // @[executor.scala 473:84]
  wire [7:0] _GEN_2082 = _GEN_8594 == 8'h3 ? _GEN_2078 : _GEN_1810; // @[executor.scala 473:84]
  wire [7:0] _GEN_2083 = _GEN_8594 == 8'h3 ? _GEN_2079 : _GEN_1811; // @[executor.scala 473:84]
  wire [7:0] _GEN_2084 = mask_2[0] ? byte_512 : _GEN_1812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2085 = mask_2[1] ? byte_513 : _GEN_1813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2086 = mask_2[2] ? byte_514 : _GEN_1814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2087 = mask_2[3] ? byte_515 : _GEN_1815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2088 = _GEN_8594 == 8'h4 ? _GEN_2084 : _GEN_1812; // @[executor.scala 473:84]
  wire [7:0] _GEN_2089 = _GEN_8594 == 8'h4 ? _GEN_2085 : _GEN_1813; // @[executor.scala 473:84]
  wire [7:0] _GEN_2090 = _GEN_8594 == 8'h4 ? _GEN_2086 : _GEN_1814; // @[executor.scala 473:84]
  wire [7:0] _GEN_2091 = _GEN_8594 == 8'h4 ? _GEN_2087 : _GEN_1815; // @[executor.scala 473:84]
  wire [7:0] _GEN_2092 = mask_2[0] ? byte_512 : _GEN_1816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2093 = mask_2[1] ? byte_513 : _GEN_1817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2094 = mask_2[2] ? byte_514 : _GEN_1818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2095 = mask_2[3] ? byte_515 : _GEN_1819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2096 = _GEN_8594 == 8'h5 ? _GEN_2092 : _GEN_1816; // @[executor.scala 473:84]
  wire [7:0] _GEN_2097 = _GEN_8594 == 8'h5 ? _GEN_2093 : _GEN_1817; // @[executor.scala 473:84]
  wire [7:0] _GEN_2098 = _GEN_8594 == 8'h5 ? _GEN_2094 : _GEN_1818; // @[executor.scala 473:84]
  wire [7:0] _GEN_2099 = _GEN_8594 == 8'h5 ? _GEN_2095 : _GEN_1819; // @[executor.scala 473:84]
  wire [7:0] _GEN_2100 = mask_2[0] ? byte_512 : _GEN_1820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2101 = mask_2[1] ? byte_513 : _GEN_1821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2102 = mask_2[2] ? byte_514 : _GEN_1822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2103 = mask_2[3] ? byte_515 : _GEN_1823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2104 = _GEN_8594 == 8'h6 ? _GEN_2100 : _GEN_1820; // @[executor.scala 473:84]
  wire [7:0] _GEN_2105 = _GEN_8594 == 8'h6 ? _GEN_2101 : _GEN_1821; // @[executor.scala 473:84]
  wire [7:0] _GEN_2106 = _GEN_8594 == 8'h6 ? _GEN_2102 : _GEN_1822; // @[executor.scala 473:84]
  wire [7:0] _GEN_2107 = _GEN_8594 == 8'h6 ? _GEN_2103 : _GEN_1823; // @[executor.scala 473:84]
  wire [7:0] _GEN_2108 = mask_2[0] ? byte_512 : _GEN_1824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2109 = mask_2[1] ? byte_513 : _GEN_1825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2110 = mask_2[2] ? byte_514 : _GEN_1826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2111 = mask_2[3] ? byte_515 : _GEN_1827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2112 = _GEN_8594 == 8'h7 ? _GEN_2108 : _GEN_1824; // @[executor.scala 473:84]
  wire [7:0] _GEN_2113 = _GEN_8594 == 8'h7 ? _GEN_2109 : _GEN_1825; // @[executor.scala 473:84]
  wire [7:0] _GEN_2114 = _GEN_8594 == 8'h7 ? _GEN_2110 : _GEN_1826; // @[executor.scala 473:84]
  wire [7:0] _GEN_2115 = _GEN_8594 == 8'h7 ? _GEN_2111 : _GEN_1827; // @[executor.scala 473:84]
  wire [7:0] _GEN_2116 = mask_2[0] ? byte_512 : _GEN_1828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2117 = mask_2[1] ? byte_513 : _GEN_1829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2118 = mask_2[2] ? byte_514 : _GEN_1830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2119 = mask_2[3] ? byte_515 : _GEN_1831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2120 = _GEN_8594 == 8'h8 ? _GEN_2116 : _GEN_1828; // @[executor.scala 473:84]
  wire [7:0] _GEN_2121 = _GEN_8594 == 8'h8 ? _GEN_2117 : _GEN_1829; // @[executor.scala 473:84]
  wire [7:0] _GEN_2122 = _GEN_8594 == 8'h8 ? _GEN_2118 : _GEN_1830; // @[executor.scala 473:84]
  wire [7:0] _GEN_2123 = _GEN_8594 == 8'h8 ? _GEN_2119 : _GEN_1831; // @[executor.scala 473:84]
  wire [7:0] _GEN_2124 = mask_2[0] ? byte_512 : _GEN_1832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2125 = mask_2[1] ? byte_513 : _GEN_1833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2126 = mask_2[2] ? byte_514 : _GEN_1834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2127 = mask_2[3] ? byte_515 : _GEN_1835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2128 = _GEN_8594 == 8'h9 ? _GEN_2124 : _GEN_1832; // @[executor.scala 473:84]
  wire [7:0] _GEN_2129 = _GEN_8594 == 8'h9 ? _GEN_2125 : _GEN_1833; // @[executor.scala 473:84]
  wire [7:0] _GEN_2130 = _GEN_8594 == 8'h9 ? _GEN_2126 : _GEN_1834; // @[executor.scala 473:84]
  wire [7:0] _GEN_2131 = _GEN_8594 == 8'h9 ? _GEN_2127 : _GEN_1835; // @[executor.scala 473:84]
  wire [7:0] _GEN_2132 = mask_2[0] ? byte_512 : _GEN_1836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2133 = mask_2[1] ? byte_513 : _GEN_1837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2134 = mask_2[2] ? byte_514 : _GEN_1838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2135 = mask_2[3] ? byte_515 : _GEN_1839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2136 = _GEN_8594 == 8'ha ? _GEN_2132 : _GEN_1836; // @[executor.scala 473:84]
  wire [7:0] _GEN_2137 = _GEN_8594 == 8'ha ? _GEN_2133 : _GEN_1837; // @[executor.scala 473:84]
  wire [7:0] _GEN_2138 = _GEN_8594 == 8'ha ? _GEN_2134 : _GEN_1838; // @[executor.scala 473:84]
  wire [7:0] _GEN_2139 = _GEN_8594 == 8'ha ? _GEN_2135 : _GEN_1839; // @[executor.scala 473:84]
  wire [7:0] _GEN_2140 = mask_2[0] ? byte_512 : _GEN_1840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2141 = mask_2[1] ? byte_513 : _GEN_1841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2142 = mask_2[2] ? byte_514 : _GEN_1842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2143 = mask_2[3] ? byte_515 : _GEN_1843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2144 = _GEN_8594 == 8'hb ? _GEN_2140 : _GEN_1840; // @[executor.scala 473:84]
  wire [7:0] _GEN_2145 = _GEN_8594 == 8'hb ? _GEN_2141 : _GEN_1841; // @[executor.scala 473:84]
  wire [7:0] _GEN_2146 = _GEN_8594 == 8'hb ? _GEN_2142 : _GEN_1842; // @[executor.scala 473:84]
  wire [7:0] _GEN_2147 = _GEN_8594 == 8'hb ? _GEN_2143 : _GEN_1843; // @[executor.scala 473:84]
  wire [7:0] _GEN_2148 = mask_2[0] ? byte_512 : _GEN_1844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2149 = mask_2[1] ? byte_513 : _GEN_1845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2150 = mask_2[2] ? byte_514 : _GEN_1846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2151 = mask_2[3] ? byte_515 : _GEN_1847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2152 = _GEN_8594 == 8'hc ? _GEN_2148 : _GEN_1844; // @[executor.scala 473:84]
  wire [7:0] _GEN_2153 = _GEN_8594 == 8'hc ? _GEN_2149 : _GEN_1845; // @[executor.scala 473:84]
  wire [7:0] _GEN_2154 = _GEN_8594 == 8'hc ? _GEN_2150 : _GEN_1846; // @[executor.scala 473:84]
  wire [7:0] _GEN_2155 = _GEN_8594 == 8'hc ? _GEN_2151 : _GEN_1847; // @[executor.scala 473:84]
  wire [7:0] _GEN_2156 = mask_2[0] ? byte_512 : _GEN_1848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2157 = mask_2[1] ? byte_513 : _GEN_1849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2158 = mask_2[2] ? byte_514 : _GEN_1850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2159 = mask_2[3] ? byte_515 : _GEN_1851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2160 = _GEN_8594 == 8'hd ? _GEN_2156 : _GEN_1848; // @[executor.scala 473:84]
  wire [7:0] _GEN_2161 = _GEN_8594 == 8'hd ? _GEN_2157 : _GEN_1849; // @[executor.scala 473:84]
  wire [7:0] _GEN_2162 = _GEN_8594 == 8'hd ? _GEN_2158 : _GEN_1850; // @[executor.scala 473:84]
  wire [7:0] _GEN_2163 = _GEN_8594 == 8'hd ? _GEN_2159 : _GEN_1851; // @[executor.scala 473:84]
  wire [7:0] _GEN_2164 = mask_2[0] ? byte_512 : _GEN_1852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2165 = mask_2[1] ? byte_513 : _GEN_1853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2166 = mask_2[2] ? byte_514 : _GEN_1854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2167 = mask_2[3] ? byte_515 : _GEN_1855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2168 = _GEN_8594 == 8'he ? _GEN_2164 : _GEN_1852; // @[executor.scala 473:84]
  wire [7:0] _GEN_2169 = _GEN_8594 == 8'he ? _GEN_2165 : _GEN_1853; // @[executor.scala 473:84]
  wire [7:0] _GEN_2170 = _GEN_8594 == 8'he ? _GEN_2166 : _GEN_1854; // @[executor.scala 473:84]
  wire [7:0] _GEN_2171 = _GEN_8594 == 8'he ? _GEN_2167 : _GEN_1855; // @[executor.scala 473:84]
  wire [7:0] _GEN_2172 = mask_2[0] ? byte_512 : _GEN_1856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2173 = mask_2[1] ? byte_513 : _GEN_1857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2174 = mask_2[2] ? byte_514 : _GEN_1858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2175 = mask_2[3] ? byte_515 : _GEN_1859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2176 = _GEN_8594 == 8'hf ? _GEN_2172 : _GEN_1856; // @[executor.scala 473:84]
  wire [7:0] _GEN_2177 = _GEN_8594 == 8'hf ? _GEN_2173 : _GEN_1857; // @[executor.scala 473:84]
  wire [7:0] _GEN_2178 = _GEN_8594 == 8'hf ? _GEN_2174 : _GEN_1858; // @[executor.scala 473:84]
  wire [7:0] _GEN_2179 = _GEN_8594 == 8'hf ? _GEN_2175 : _GEN_1859; // @[executor.scala 473:84]
  wire [7:0] _GEN_2180 = mask_2[0] ? byte_512 : _GEN_1860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2181 = mask_2[1] ? byte_513 : _GEN_1861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2182 = mask_2[2] ? byte_514 : _GEN_1862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2183 = mask_2[3] ? byte_515 : _GEN_1863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2184 = _GEN_8594 == 8'h10 ? _GEN_2180 : _GEN_1860; // @[executor.scala 473:84]
  wire [7:0] _GEN_2185 = _GEN_8594 == 8'h10 ? _GEN_2181 : _GEN_1861; // @[executor.scala 473:84]
  wire [7:0] _GEN_2186 = _GEN_8594 == 8'h10 ? _GEN_2182 : _GEN_1862; // @[executor.scala 473:84]
  wire [7:0] _GEN_2187 = _GEN_8594 == 8'h10 ? _GEN_2183 : _GEN_1863; // @[executor.scala 473:84]
  wire [7:0] _GEN_2188 = mask_2[0] ? byte_512 : _GEN_1864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2189 = mask_2[1] ? byte_513 : _GEN_1865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2190 = mask_2[2] ? byte_514 : _GEN_1866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2191 = mask_2[3] ? byte_515 : _GEN_1867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2192 = _GEN_8594 == 8'h11 ? _GEN_2188 : _GEN_1864; // @[executor.scala 473:84]
  wire [7:0] _GEN_2193 = _GEN_8594 == 8'h11 ? _GEN_2189 : _GEN_1865; // @[executor.scala 473:84]
  wire [7:0] _GEN_2194 = _GEN_8594 == 8'h11 ? _GEN_2190 : _GEN_1866; // @[executor.scala 473:84]
  wire [7:0] _GEN_2195 = _GEN_8594 == 8'h11 ? _GEN_2191 : _GEN_1867; // @[executor.scala 473:84]
  wire [7:0] _GEN_2196 = mask_2[0] ? byte_512 : _GEN_1868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2197 = mask_2[1] ? byte_513 : _GEN_1869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2198 = mask_2[2] ? byte_514 : _GEN_1870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2199 = mask_2[3] ? byte_515 : _GEN_1871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2200 = _GEN_8594 == 8'h12 ? _GEN_2196 : _GEN_1868; // @[executor.scala 473:84]
  wire [7:0] _GEN_2201 = _GEN_8594 == 8'h12 ? _GEN_2197 : _GEN_1869; // @[executor.scala 473:84]
  wire [7:0] _GEN_2202 = _GEN_8594 == 8'h12 ? _GEN_2198 : _GEN_1870; // @[executor.scala 473:84]
  wire [7:0] _GEN_2203 = _GEN_8594 == 8'h12 ? _GEN_2199 : _GEN_1871; // @[executor.scala 473:84]
  wire [7:0] _GEN_2204 = mask_2[0] ? byte_512 : _GEN_1872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2205 = mask_2[1] ? byte_513 : _GEN_1873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2206 = mask_2[2] ? byte_514 : _GEN_1874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2207 = mask_2[3] ? byte_515 : _GEN_1875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2208 = _GEN_8594 == 8'h13 ? _GEN_2204 : _GEN_1872; // @[executor.scala 473:84]
  wire [7:0] _GEN_2209 = _GEN_8594 == 8'h13 ? _GEN_2205 : _GEN_1873; // @[executor.scala 473:84]
  wire [7:0] _GEN_2210 = _GEN_8594 == 8'h13 ? _GEN_2206 : _GEN_1874; // @[executor.scala 473:84]
  wire [7:0] _GEN_2211 = _GEN_8594 == 8'h13 ? _GEN_2207 : _GEN_1875; // @[executor.scala 473:84]
  wire [7:0] _GEN_2212 = mask_2[0] ? byte_512 : _GEN_1876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2213 = mask_2[1] ? byte_513 : _GEN_1877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2214 = mask_2[2] ? byte_514 : _GEN_1878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2215 = mask_2[3] ? byte_515 : _GEN_1879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2216 = _GEN_8594 == 8'h14 ? _GEN_2212 : _GEN_1876; // @[executor.scala 473:84]
  wire [7:0] _GEN_2217 = _GEN_8594 == 8'h14 ? _GEN_2213 : _GEN_1877; // @[executor.scala 473:84]
  wire [7:0] _GEN_2218 = _GEN_8594 == 8'h14 ? _GEN_2214 : _GEN_1878; // @[executor.scala 473:84]
  wire [7:0] _GEN_2219 = _GEN_8594 == 8'h14 ? _GEN_2215 : _GEN_1879; // @[executor.scala 473:84]
  wire [7:0] _GEN_2220 = mask_2[0] ? byte_512 : _GEN_1880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2221 = mask_2[1] ? byte_513 : _GEN_1881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2222 = mask_2[2] ? byte_514 : _GEN_1882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2223 = mask_2[3] ? byte_515 : _GEN_1883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2224 = _GEN_8594 == 8'h15 ? _GEN_2220 : _GEN_1880; // @[executor.scala 473:84]
  wire [7:0] _GEN_2225 = _GEN_8594 == 8'h15 ? _GEN_2221 : _GEN_1881; // @[executor.scala 473:84]
  wire [7:0] _GEN_2226 = _GEN_8594 == 8'h15 ? _GEN_2222 : _GEN_1882; // @[executor.scala 473:84]
  wire [7:0] _GEN_2227 = _GEN_8594 == 8'h15 ? _GEN_2223 : _GEN_1883; // @[executor.scala 473:84]
  wire [7:0] _GEN_2228 = mask_2[0] ? byte_512 : _GEN_1884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2229 = mask_2[1] ? byte_513 : _GEN_1885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2230 = mask_2[2] ? byte_514 : _GEN_1886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2231 = mask_2[3] ? byte_515 : _GEN_1887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2232 = _GEN_8594 == 8'h16 ? _GEN_2228 : _GEN_1884; // @[executor.scala 473:84]
  wire [7:0] _GEN_2233 = _GEN_8594 == 8'h16 ? _GEN_2229 : _GEN_1885; // @[executor.scala 473:84]
  wire [7:0] _GEN_2234 = _GEN_8594 == 8'h16 ? _GEN_2230 : _GEN_1886; // @[executor.scala 473:84]
  wire [7:0] _GEN_2235 = _GEN_8594 == 8'h16 ? _GEN_2231 : _GEN_1887; // @[executor.scala 473:84]
  wire [7:0] _GEN_2236 = mask_2[0] ? byte_512 : _GEN_1888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2237 = mask_2[1] ? byte_513 : _GEN_1889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2238 = mask_2[2] ? byte_514 : _GEN_1890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2239 = mask_2[3] ? byte_515 : _GEN_1891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2240 = _GEN_8594 == 8'h17 ? _GEN_2236 : _GEN_1888; // @[executor.scala 473:84]
  wire [7:0] _GEN_2241 = _GEN_8594 == 8'h17 ? _GEN_2237 : _GEN_1889; // @[executor.scala 473:84]
  wire [7:0] _GEN_2242 = _GEN_8594 == 8'h17 ? _GEN_2238 : _GEN_1890; // @[executor.scala 473:84]
  wire [7:0] _GEN_2243 = _GEN_8594 == 8'h17 ? _GEN_2239 : _GEN_1891; // @[executor.scala 473:84]
  wire [7:0] _GEN_2244 = mask_2[0] ? byte_512 : _GEN_1892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2245 = mask_2[1] ? byte_513 : _GEN_1893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2246 = mask_2[2] ? byte_514 : _GEN_1894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2247 = mask_2[3] ? byte_515 : _GEN_1895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2248 = _GEN_8594 == 8'h18 ? _GEN_2244 : _GEN_1892; // @[executor.scala 473:84]
  wire [7:0] _GEN_2249 = _GEN_8594 == 8'h18 ? _GEN_2245 : _GEN_1893; // @[executor.scala 473:84]
  wire [7:0] _GEN_2250 = _GEN_8594 == 8'h18 ? _GEN_2246 : _GEN_1894; // @[executor.scala 473:84]
  wire [7:0] _GEN_2251 = _GEN_8594 == 8'h18 ? _GEN_2247 : _GEN_1895; // @[executor.scala 473:84]
  wire [7:0] _GEN_2252 = mask_2[0] ? byte_512 : _GEN_1896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2253 = mask_2[1] ? byte_513 : _GEN_1897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2254 = mask_2[2] ? byte_514 : _GEN_1898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2255 = mask_2[3] ? byte_515 : _GEN_1899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2256 = _GEN_8594 == 8'h19 ? _GEN_2252 : _GEN_1896; // @[executor.scala 473:84]
  wire [7:0] _GEN_2257 = _GEN_8594 == 8'h19 ? _GEN_2253 : _GEN_1897; // @[executor.scala 473:84]
  wire [7:0] _GEN_2258 = _GEN_8594 == 8'h19 ? _GEN_2254 : _GEN_1898; // @[executor.scala 473:84]
  wire [7:0] _GEN_2259 = _GEN_8594 == 8'h19 ? _GEN_2255 : _GEN_1899; // @[executor.scala 473:84]
  wire [7:0] _GEN_2260 = mask_2[0] ? byte_512 : _GEN_1900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2261 = mask_2[1] ? byte_513 : _GEN_1901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2262 = mask_2[2] ? byte_514 : _GEN_1902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2263 = mask_2[3] ? byte_515 : _GEN_1903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2264 = _GEN_8594 == 8'h1a ? _GEN_2260 : _GEN_1900; // @[executor.scala 473:84]
  wire [7:0] _GEN_2265 = _GEN_8594 == 8'h1a ? _GEN_2261 : _GEN_1901; // @[executor.scala 473:84]
  wire [7:0] _GEN_2266 = _GEN_8594 == 8'h1a ? _GEN_2262 : _GEN_1902; // @[executor.scala 473:84]
  wire [7:0] _GEN_2267 = _GEN_8594 == 8'h1a ? _GEN_2263 : _GEN_1903; // @[executor.scala 473:84]
  wire [7:0] _GEN_2268 = mask_2[0] ? byte_512 : _GEN_1904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2269 = mask_2[1] ? byte_513 : _GEN_1905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2270 = mask_2[2] ? byte_514 : _GEN_1906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2271 = mask_2[3] ? byte_515 : _GEN_1907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2272 = _GEN_8594 == 8'h1b ? _GEN_2268 : _GEN_1904; // @[executor.scala 473:84]
  wire [7:0] _GEN_2273 = _GEN_8594 == 8'h1b ? _GEN_2269 : _GEN_1905; // @[executor.scala 473:84]
  wire [7:0] _GEN_2274 = _GEN_8594 == 8'h1b ? _GEN_2270 : _GEN_1906; // @[executor.scala 473:84]
  wire [7:0] _GEN_2275 = _GEN_8594 == 8'h1b ? _GEN_2271 : _GEN_1907; // @[executor.scala 473:84]
  wire [7:0] _GEN_2276 = mask_2[0] ? byte_512 : _GEN_1908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2277 = mask_2[1] ? byte_513 : _GEN_1909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2278 = mask_2[2] ? byte_514 : _GEN_1910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2279 = mask_2[3] ? byte_515 : _GEN_1911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2280 = _GEN_8594 == 8'h1c ? _GEN_2276 : _GEN_1908; // @[executor.scala 473:84]
  wire [7:0] _GEN_2281 = _GEN_8594 == 8'h1c ? _GEN_2277 : _GEN_1909; // @[executor.scala 473:84]
  wire [7:0] _GEN_2282 = _GEN_8594 == 8'h1c ? _GEN_2278 : _GEN_1910; // @[executor.scala 473:84]
  wire [7:0] _GEN_2283 = _GEN_8594 == 8'h1c ? _GEN_2279 : _GEN_1911; // @[executor.scala 473:84]
  wire [7:0] _GEN_2284 = mask_2[0] ? byte_512 : _GEN_1912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2285 = mask_2[1] ? byte_513 : _GEN_1913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2286 = mask_2[2] ? byte_514 : _GEN_1914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2287 = mask_2[3] ? byte_515 : _GEN_1915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2288 = _GEN_8594 == 8'h1d ? _GEN_2284 : _GEN_1912; // @[executor.scala 473:84]
  wire [7:0] _GEN_2289 = _GEN_8594 == 8'h1d ? _GEN_2285 : _GEN_1913; // @[executor.scala 473:84]
  wire [7:0] _GEN_2290 = _GEN_8594 == 8'h1d ? _GEN_2286 : _GEN_1914; // @[executor.scala 473:84]
  wire [7:0] _GEN_2291 = _GEN_8594 == 8'h1d ? _GEN_2287 : _GEN_1915; // @[executor.scala 473:84]
  wire [7:0] _GEN_2292 = mask_2[0] ? byte_512 : _GEN_1916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2293 = mask_2[1] ? byte_513 : _GEN_1917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2294 = mask_2[2] ? byte_514 : _GEN_1918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2295 = mask_2[3] ? byte_515 : _GEN_1919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2296 = _GEN_8594 == 8'h1e ? _GEN_2292 : _GEN_1916; // @[executor.scala 473:84]
  wire [7:0] _GEN_2297 = _GEN_8594 == 8'h1e ? _GEN_2293 : _GEN_1917; // @[executor.scala 473:84]
  wire [7:0] _GEN_2298 = _GEN_8594 == 8'h1e ? _GEN_2294 : _GEN_1918; // @[executor.scala 473:84]
  wire [7:0] _GEN_2299 = _GEN_8594 == 8'h1e ? _GEN_2295 : _GEN_1919; // @[executor.scala 473:84]
  wire [7:0] _GEN_2300 = mask_2[0] ? byte_512 : _GEN_1920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2301 = mask_2[1] ? byte_513 : _GEN_1921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2302 = mask_2[2] ? byte_514 : _GEN_1922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2303 = mask_2[3] ? byte_515 : _GEN_1923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2304 = _GEN_8594 == 8'h1f ? _GEN_2300 : _GEN_1920; // @[executor.scala 473:84]
  wire [7:0] _GEN_2305 = _GEN_8594 == 8'h1f ? _GEN_2301 : _GEN_1921; // @[executor.scala 473:84]
  wire [7:0] _GEN_2306 = _GEN_8594 == 8'h1f ? _GEN_2302 : _GEN_1922; // @[executor.scala 473:84]
  wire [7:0] _GEN_2307 = _GEN_8594 == 8'h1f ? _GEN_2303 : _GEN_1923; // @[executor.scala 473:84]
  wire [7:0] _GEN_2308 = mask_2[0] ? byte_512 : _GEN_1924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2309 = mask_2[1] ? byte_513 : _GEN_1925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2310 = mask_2[2] ? byte_514 : _GEN_1926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2311 = mask_2[3] ? byte_515 : _GEN_1927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2312 = _GEN_8594 == 8'h20 ? _GEN_2308 : _GEN_1924; // @[executor.scala 473:84]
  wire [7:0] _GEN_2313 = _GEN_8594 == 8'h20 ? _GEN_2309 : _GEN_1925; // @[executor.scala 473:84]
  wire [7:0] _GEN_2314 = _GEN_8594 == 8'h20 ? _GEN_2310 : _GEN_1926; // @[executor.scala 473:84]
  wire [7:0] _GEN_2315 = _GEN_8594 == 8'h20 ? _GEN_2311 : _GEN_1927; // @[executor.scala 473:84]
  wire [7:0] _GEN_2316 = mask_2[0] ? byte_512 : _GEN_1928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2317 = mask_2[1] ? byte_513 : _GEN_1929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2318 = mask_2[2] ? byte_514 : _GEN_1930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2319 = mask_2[3] ? byte_515 : _GEN_1931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2320 = _GEN_8594 == 8'h21 ? _GEN_2316 : _GEN_1928; // @[executor.scala 473:84]
  wire [7:0] _GEN_2321 = _GEN_8594 == 8'h21 ? _GEN_2317 : _GEN_1929; // @[executor.scala 473:84]
  wire [7:0] _GEN_2322 = _GEN_8594 == 8'h21 ? _GEN_2318 : _GEN_1930; // @[executor.scala 473:84]
  wire [7:0] _GEN_2323 = _GEN_8594 == 8'h21 ? _GEN_2319 : _GEN_1931; // @[executor.scala 473:84]
  wire [7:0] _GEN_2324 = mask_2[0] ? byte_512 : _GEN_1932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2325 = mask_2[1] ? byte_513 : _GEN_1933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2326 = mask_2[2] ? byte_514 : _GEN_1934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2327 = mask_2[3] ? byte_515 : _GEN_1935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2328 = _GEN_8594 == 8'h22 ? _GEN_2324 : _GEN_1932; // @[executor.scala 473:84]
  wire [7:0] _GEN_2329 = _GEN_8594 == 8'h22 ? _GEN_2325 : _GEN_1933; // @[executor.scala 473:84]
  wire [7:0] _GEN_2330 = _GEN_8594 == 8'h22 ? _GEN_2326 : _GEN_1934; // @[executor.scala 473:84]
  wire [7:0] _GEN_2331 = _GEN_8594 == 8'h22 ? _GEN_2327 : _GEN_1935; // @[executor.scala 473:84]
  wire [7:0] _GEN_2332 = mask_2[0] ? byte_512 : _GEN_1936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2333 = mask_2[1] ? byte_513 : _GEN_1937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2334 = mask_2[2] ? byte_514 : _GEN_1938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2335 = mask_2[3] ? byte_515 : _GEN_1939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2336 = _GEN_8594 == 8'h23 ? _GEN_2332 : _GEN_1936; // @[executor.scala 473:84]
  wire [7:0] _GEN_2337 = _GEN_8594 == 8'h23 ? _GEN_2333 : _GEN_1937; // @[executor.scala 473:84]
  wire [7:0] _GEN_2338 = _GEN_8594 == 8'h23 ? _GEN_2334 : _GEN_1938; // @[executor.scala 473:84]
  wire [7:0] _GEN_2339 = _GEN_8594 == 8'h23 ? _GEN_2335 : _GEN_1939; // @[executor.scala 473:84]
  wire [7:0] _GEN_2340 = mask_2[0] ? byte_512 : _GEN_1940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2341 = mask_2[1] ? byte_513 : _GEN_1941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2342 = mask_2[2] ? byte_514 : _GEN_1942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2343 = mask_2[3] ? byte_515 : _GEN_1943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2344 = _GEN_8594 == 8'h24 ? _GEN_2340 : _GEN_1940; // @[executor.scala 473:84]
  wire [7:0] _GEN_2345 = _GEN_8594 == 8'h24 ? _GEN_2341 : _GEN_1941; // @[executor.scala 473:84]
  wire [7:0] _GEN_2346 = _GEN_8594 == 8'h24 ? _GEN_2342 : _GEN_1942; // @[executor.scala 473:84]
  wire [7:0] _GEN_2347 = _GEN_8594 == 8'h24 ? _GEN_2343 : _GEN_1943; // @[executor.scala 473:84]
  wire [7:0] _GEN_2348 = mask_2[0] ? byte_512 : _GEN_1944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2349 = mask_2[1] ? byte_513 : _GEN_1945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2350 = mask_2[2] ? byte_514 : _GEN_1946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2351 = mask_2[3] ? byte_515 : _GEN_1947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2352 = _GEN_8594 == 8'h25 ? _GEN_2348 : _GEN_1944; // @[executor.scala 473:84]
  wire [7:0] _GEN_2353 = _GEN_8594 == 8'h25 ? _GEN_2349 : _GEN_1945; // @[executor.scala 473:84]
  wire [7:0] _GEN_2354 = _GEN_8594 == 8'h25 ? _GEN_2350 : _GEN_1946; // @[executor.scala 473:84]
  wire [7:0] _GEN_2355 = _GEN_8594 == 8'h25 ? _GEN_2351 : _GEN_1947; // @[executor.scala 473:84]
  wire [7:0] _GEN_2356 = mask_2[0] ? byte_512 : _GEN_1948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2357 = mask_2[1] ? byte_513 : _GEN_1949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2358 = mask_2[2] ? byte_514 : _GEN_1950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2359 = mask_2[3] ? byte_515 : _GEN_1951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2360 = _GEN_8594 == 8'h26 ? _GEN_2356 : _GEN_1948; // @[executor.scala 473:84]
  wire [7:0] _GEN_2361 = _GEN_8594 == 8'h26 ? _GEN_2357 : _GEN_1949; // @[executor.scala 473:84]
  wire [7:0] _GEN_2362 = _GEN_8594 == 8'h26 ? _GEN_2358 : _GEN_1950; // @[executor.scala 473:84]
  wire [7:0] _GEN_2363 = _GEN_8594 == 8'h26 ? _GEN_2359 : _GEN_1951; // @[executor.scala 473:84]
  wire [7:0] _GEN_2364 = mask_2[0] ? byte_512 : _GEN_1952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2365 = mask_2[1] ? byte_513 : _GEN_1953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2366 = mask_2[2] ? byte_514 : _GEN_1954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2367 = mask_2[3] ? byte_515 : _GEN_1955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2368 = _GEN_8594 == 8'h27 ? _GEN_2364 : _GEN_1952; // @[executor.scala 473:84]
  wire [7:0] _GEN_2369 = _GEN_8594 == 8'h27 ? _GEN_2365 : _GEN_1953; // @[executor.scala 473:84]
  wire [7:0] _GEN_2370 = _GEN_8594 == 8'h27 ? _GEN_2366 : _GEN_1954; // @[executor.scala 473:84]
  wire [7:0] _GEN_2371 = _GEN_8594 == 8'h27 ? _GEN_2367 : _GEN_1955; // @[executor.scala 473:84]
  wire [7:0] _GEN_2372 = mask_2[0] ? byte_512 : _GEN_1956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2373 = mask_2[1] ? byte_513 : _GEN_1957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2374 = mask_2[2] ? byte_514 : _GEN_1958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2375 = mask_2[3] ? byte_515 : _GEN_1959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2376 = _GEN_8594 == 8'h28 ? _GEN_2372 : _GEN_1956; // @[executor.scala 473:84]
  wire [7:0] _GEN_2377 = _GEN_8594 == 8'h28 ? _GEN_2373 : _GEN_1957; // @[executor.scala 473:84]
  wire [7:0] _GEN_2378 = _GEN_8594 == 8'h28 ? _GEN_2374 : _GEN_1958; // @[executor.scala 473:84]
  wire [7:0] _GEN_2379 = _GEN_8594 == 8'h28 ? _GEN_2375 : _GEN_1959; // @[executor.scala 473:84]
  wire [7:0] _GEN_2380 = mask_2[0] ? byte_512 : _GEN_1960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2381 = mask_2[1] ? byte_513 : _GEN_1961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2382 = mask_2[2] ? byte_514 : _GEN_1962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2383 = mask_2[3] ? byte_515 : _GEN_1963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2384 = _GEN_8594 == 8'h29 ? _GEN_2380 : _GEN_1960; // @[executor.scala 473:84]
  wire [7:0] _GEN_2385 = _GEN_8594 == 8'h29 ? _GEN_2381 : _GEN_1961; // @[executor.scala 473:84]
  wire [7:0] _GEN_2386 = _GEN_8594 == 8'h29 ? _GEN_2382 : _GEN_1962; // @[executor.scala 473:84]
  wire [7:0] _GEN_2387 = _GEN_8594 == 8'h29 ? _GEN_2383 : _GEN_1963; // @[executor.scala 473:84]
  wire [7:0] _GEN_2388 = mask_2[0] ? byte_512 : _GEN_1964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2389 = mask_2[1] ? byte_513 : _GEN_1965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2390 = mask_2[2] ? byte_514 : _GEN_1966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2391 = mask_2[3] ? byte_515 : _GEN_1967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2392 = _GEN_8594 == 8'h2a ? _GEN_2388 : _GEN_1964; // @[executor.scala 473:84]
  wire [7:0] _GEN_2393 = _GEN_8594 == 8'h2a ? _GEN_2389 : _GEN_1965; // @[executor.scala 473:84]
  wire [7:0] _GEN_2394 = _GEN_8594 == 8'h2a ? _GEN_2390 : _GEN_1966; // @[executor.scala 473:84]
  wire [7:0] _GEN_2395 = _GEN_8594 == 8'h2a ? _GEN_2391 : _GEN_1967; // @[executor.scala 473:84]
  wire [7:0] _GEN_2396 = mask_2[0] ? byte_512 : _GEN_1968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2397 = mask_2[1] ? byte_513 : _GEN_1969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2398 = mask_2[2] ? byte_514 : _GEN_1970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2399 = mask_2[3] ? byte_515 : _GEN_1971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2400 = _GEN_8594 == 8'h2b ? _GEN_2396 : _GEN_1968; // @[executor.scala 473:84]
  wire [7:0] _GEN_2401 = _GEN_8594 == 8'h2b ? _GEN_2397 : _GEN_1969; // @[executor.scala 473:84]
  wire [7:0] _GEN_2402 = _GEN_8594 == 8'h2b ? _GEN_2398 : _GEN_1970; // @[executor.scala 473:84]
  wire [7:0] _GEN_2403 = _GEN_8594 == 8'h2b ? _GEN_2399 : _GEN_1971; // @[executor.scala 473:84]
  wire [7:0] _GEN_2404 = mask_2[0] ? byte_512 : _GEN_1972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2405 = mask_2[1] ? byte_513 : _GEN_1973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2406 = mask_2[2] ? byte_514 : _GEN_1974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2407 = mask_2[3] ? byte_515 : _GEN_1975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2408 = _GEN_8594 == 8'h2c ? _GEN_2404 : _GEN_1972; // @[executor.scala 473:84]
  wire [7:0] _GEN_2409 = _GEN_8594 == 8'h2c ? _GEN_2405 : _GEN_1973; // @[executor.scala 473:84]
  wire [7:0] _GEN_2410 = _GEN_8594 == 8'h2c ? _GEN_2406 : _GEN_1974; // @[executor.scala 473:84]
  wire [7:0] _GEN_2411 = _GEN_8594 == 8'h2c ? _GEN_2407 : _GEN_1975; // @[executor.scala 473:84]
  wire [7:0] _GEN_2412 = mask_2[0] ? byte_512 : _GEN_1976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2413 = mask_2[1] ? byte_513 : _GEN_1977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2414 = mask_2[2] ? byte_514 : _GEN_1978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2415 = mask_2[3] ? byte_515 : _GEN_1979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2416 = _GEN_8594 == 8'h2d ? _GEN_2412 : _GEN_1976; // @[executor.scala 473:84]
  wire [7:0] _GEN_2417 = _GEN_8594 == 8'h2d ? _GEN_2413 : _GEN_1977; // @[executor.scala 473:84]
  wire [7:0] _GEN_2418 = _GEN_8594 == 8'h2d ? _GEN_2414 : _GEN_1978; // @[executor.scala 473:84]
  wire [7:0] _GEN_2419 = _GEN_8594 == 8'h2d ? _GEN_2415 : _GEN_1979; // @[executor.scala 473:84]
  wire [7:0] _GEN_2420 = mask_2[0] ? byte_512 : _GEN_1980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2421 = mask_2[1] ? byte_513 : _GEN_1981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2422 = mask_2[2] ? byte_514 : _GEN_1982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2423 = mask_2[3] ? byte_515 : _GEN_1983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2424 = _GEN_8594 == 8'h2e ? _GEN_2420 : _GEN_1980; // @[executor.scala 473:84]
  wire [7:0] _GEN_2425 = _GEN_8594 == 8'h2e ? _GEN_2421 : _GEN_1981; // @[executor.scala 473:84]
  wire [7:0] _GEN_2426 = _GEN_8594 == 8'h2e ? _GEN_2422 : _GEN_1982; // @[executor.scala 473:84]
  wire [7:0] _GEN_2427 = _GEN_8594 == 8'h2e ? _GEN_2423 : _GEN_1983; // @[executor.scala 473:84]
  wire [7:0] _GEN_2428 = mask_2[0] ? byte_512 : _GEN_1984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2429 = mask_2[1] ? byte_513 : _GEN_1985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2430 = mask_2[2] ? byte_514 : _GEN_1986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2431 = mask_2[3] ? byte_515 : _GEN_1987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2432 = _GEN_8594 == 8'h2f ? _GEN_2428 : _GEN_1984; // @[executor.scala 473:84]
  wire [7:0] _GEN_2433 = _GEN_8594 == 8'h2f ? _GEN_2429 : _GEN_1985; // @[executor.scala 473:84]
  wire [7:0] _GEN_2434 = _GEN_8594 == 8'h2f ? _GEN_2430 : _GEN_1986; // @[executor.scala 473:84]
  wire [7:0] _GEN_2435 = _GEN_8594 == 8'h2f ? _GEN_2431 : _GEN_1987; // @[executor.scala 473:84]
  wire [7:0] _GEN_2436 = mask_2[0] ? byte_512 : _GEN_1988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2437 = mask_2[1] ? byte_513 : _GEN_1989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2438 = mask_2[2] ? byte_514 : _GEN_1990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2439 = mask_2[3] ? byte_515 : _GEN_1991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2440 = _GEN_8594 == 8'h30 ? _GEN_2436 : _GEN_1988; // @[executor.scala 473:84]
  wire [7:0] _GEN_2441 = _GEN_8594 == 8'h30 ? _GEN_2437 : _GEN_1989; // @[executor.scala 473:84]
  wire [7:0] _GEN_2442 = _GEN_8594 == 8'h30 ? _GEN_2438 : _GEN_1990; // @[executor.scala 473:84]
  wire [7:0] _GEN_2443 = _GEN_8594 == 8'h30 ? _GEN_2439 : _GEN_1991; // @[executor.scala 473:84]
  wire [7:0] _GEN_2444 = mask_2[0] ? byte_512 : _GEN_1992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2445 = mask_2[1] ? byte_513 : _GEN_1993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2446 = mask_2[2] ? byte_514 : _GEN_1994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2447 = mask_2[3] ? byte_515 : _GEN_1995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2448 = _GEN_8594 == 8'h31 ? _GEN_2444 : _GEN_1992; // @[executor.scala 473:84]
  wire [7:0] _GEN_2449 = _GEN_8594 == 8'h31 ? _GEN_2445 : _GEN_1993; // @[executor.scala 473:84]
  wire [7:0] _GEN_2450 = _GEN_8594 == 8'h31 ? _GEN_2446 : _GEN_1994; // @[executor.scala 473:84]
  wire [7:0] _GEN_2451 = _GEN_8594 == 8'h31 ? _GEN_2447 : _GEN_1995; // @[executor.scala 473:84]
  wire [7:0] _GEN_2452 = mask_2[0] ? byte_512 : _GEN_1996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2453 = mask_2[1] ? byte_513 : _GEN_1997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2454 = mask_2[2] ? byte_514 : _GEN_1998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2455 = mask_2[3] ? byte_515 : _GEN_1999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2456 = _GEN_8594 == 8'h32 ? _GEN_2452 : _GEN_1996; // @[executor.scala 473:84]
  wire [7:0] _GEN_2457 = _GEN_8594 == 8'h32 ? _GEN_2453 : _GEN_1997; // @[executor.scala 473:84]
  wire [7:0] _GEN_2458 = _GEN_8594 == 8'h32 ? _GEN_2454 : _GEN_1998; // @[executor.scala 473:84]
  wire [7:0] _GEN_2459 = _GEN_8594 == 8'h32 ? _GEN_2455 : _GEN_1999; // @[executor.scala 473:84]
  wire [7:0] _GEN_2460 = mask_2[0] ? byte_512 : _GEN_2000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2461 = mask_2[1] ? byte_513 : _GEN_2001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2462 = mask_2[2] ? byte_514 : _GEN_2002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2463 = mask_2[3] ? byte_515 : _GEN_2003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2464 = _GEN_8594 == 8'h33 ? _GEN_2460 : _GEN_2000; // @[executor.scala 473:84]
  wire [7:0] _GEN_2465 = _GEN_8594 == 8'h33 ? _GEN_2461 : _GEN_2001; // @[executor.scala 473:84]
  wire [7:0] _GEN_2466 = _GEN_8594 == 8'h33 ? _GEN_2462 : _GEN_2002; // @[executor.scala 473:84]
  wire [7:0] _GEN_2467 = _GEN_8594 == 8'h33 ? _GEN_2463 : _GEN_2003; // @[executor.scala 473:84]
  wire [7:0] _GEN_2468 = mask_2[0] ? byte_512 : _GEN_2004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2469 = mask_2[1] ? byte_513 : _GEN_2005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2470 = mask_2[2] ? byte_514 : _GEN_2006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2471 = mask_2[3] ? byte_515 : _GEN_2007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2472 = _GEN_8594 == 8'h34 ? _GEN_2468 : _GEN_2004; // @[executor.scala 473:84]
  wire [7:0] _GEN_2473 = _GEN_8594 == 8'h34 ? _GEN_2469 : _GEN_2005; // @[executor.scala 473:84]
  wire [7:0] _GEN_2474 = _GEN_8594 == 8'h34 ? _GEN_2470 : _GEN_2006; // @[executor.scala 473:84]
  wire [7:0] _GEN_2475 = _GEN_8594 == 8'h34 ? _GEN_2471 : _GEN_2007; // @[executor.scala 473:84]
  wire [7:0] _GEN_2476 = mask_2[0] ? byte_512 : _GEN_2008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2477 = mask_2[1] ? byte_513 : _GEN_2009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2478 = mask_2[2] ? byte_514 : _GEN_2010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2479 = mask_2[3] ? byte_515 : _GEN_2011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2480 = _GEN_8594 == 8'h35 ? _GEN_2476 : _GEN_2008; // @[executor.scala 473:84]
  wire [7:0] _GEN_2481 = _GEN_8594 == 8'h35 ? _GEN_2477 : _GEN_2009; // @[executor.scala 473:84]
  wire [7:0] _GEN_2482 = _GEN_8594 == 8'h35 ? _GEN_2478 : _GEN_2010; // @[executor.scala 473:84]
  wire [7:0] _GEN_2483 = _GEN_8594 == 8'h35 ? _GEN_2479 : _GEN_2011; // @[executor.scala 473:84]
  wire [7:0] _GEN_2484 = mask_2[0] ? byte_512 : _GEN_2012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2485 = mask_2[1] ? byte_513 : _GEN_2013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2486 = mask_2[2] ? byte_514 : _GEN_2014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2487 = mask_2[3] ? byte_515 : _GEN_2015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2488 = _GEN_8594 == 8'h36 ? _GEN_2484 : _GEN_2012; // @[executor.scala 473:84]
  wire [7:0] _GEN_2489 = _GEN_8594 == 8'h36 ? _GEN_2485 : _GEN_2013; // @[executor.scala 473:84]
  wire [7:0] _GEN_2490 = _GEN_8594 == 8'h36 ? _GEN_2486 : _GEN_2014; // @[executor.scala 473:84]
  wire [7:0] _GEN_2491 = _GEN_8594 == 8'h36 ? _GEN_2487 : _GEN_2015; // @[executor.scala 473:84]
  wire [7:0] _GEN_2492 = mask_2[0] ? byte_512 : _GEN_2016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2493 = mask_2[1] ? byte_513 : _GEN_2017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2494 = mask_2[2] ? byte_514 : _GEN_2018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2495 = mask_2[3] ? byte_515 : _GEN_2019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2496 = _GEN_8594 == 8'h37 ? _GEN_2492 : _GEN_2016; // @[executor.scala 473:84]
  wire [7:0] _GEN_2497 = _GEN_8594 == 8'h37 ? _GEN_2493 : _GEN_2017; // @[executor.scala 473:84]
  wire [7:0] _GEN_2498 = _GEN_8594 == 8'h37 ? _GEN_2494 : _GEN_2018; // @[executor.scala 473:84]
  wire [7:0] _GEN_2499 = _GEN_8594 == 8'h37 ? _GEN_2495 : _GEN_2019; // @[executor.scala 473:84]
  wire [7:0] _GEN_2500 = mask_2[0] ? byte_512 : _GEN_2020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2501 = mask_2[1] ? byte_513 : _GEN_2021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2502 = mask_2[2] ? byte_514 : _GEN_2022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2503 = mask_2[3] ? byte_515 : _GEN_2023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2504 = _GEN_8594 == 8'h38 ? _GEN_2500 : _GEN_2020; // @[executor.scala 473:84]
  wire [7:0] _GEN_2505 = _GEN_8594 == 8'h38 ? _GEN_2501 : _GEN_2021; // @[executor.scala 473:84]
  wire [7:0] _GEN_2506 = _GEN_8594 == 8'h38 ? _GEN_2502 : _GEN_2022; // @[executor.scala 473:84]
  wire [7:0] _GEN_2507 = _GEN_8594 == 8'h38 ? _GEN_2503 : _GEN_2023; // @[executor.scala 473:84]
  wire [7:0] _GEN_2508 = mask_2[0] ? byte_512 : _GEN_2024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2509 = mask_2[1] ? byte_513 : _GEN_2025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2510 = mask_2[2] ? byte_514 : _GEN_2026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2511 = mask_2[3] ? byte_515 : _GEN_2027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2512 = _GEN_8594 == 8'h39 ? _GEN_2508 : _GEN_2024; // @[executor.scala 473:84]
  wire [7:0] _GEN_2513 = _GEN_8594 == 8'h39 ? _GEN_2509 : _GEN_2025; // @[executor.scala 473:84]
  wire [7:0] _GEN_2514 = _GEN_8594 == 8'h39 ? _GEN_2510 : _GEN_2026; // @[executor.scala 473:84]
  wire [7:0] _GEN_2515 = _GEN_8594 == 8'h39 ? _GEN_2511 : _GEN_2027; // @[executor.scala 473:84]
  wire [7:0] _GEN_2516 = mask_2[0] ? byte_512 : _GEN_2028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2517 = mask_2[1] ? byte_513 : _GEN_2029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2518 = mask_2[2] ? byte_514 : _GEN_2030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2519 = mask_2[3] ? byte_515 : _GEN_2031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2520 = _GEN_8594 == 8'h3a ? _GEN_2516 : _GEN_2028; // @[executor.scala 473:84]
  wire [7:0] _GEN_2521 = _GEN_8594 == 8'h3a ? _GEN_2517 : _GEN_2029; // @[executor.scala 473:84]
  wire [7:0] _GEN_2522 = _GEN_8594 == 8'h3a ? _GEN_2518 : _GEN_2030; // @[executor.scala 473:84]
  wire [7:0] _GEN_2523 = _GEN_8594 == 8'h3a ? _GEN_2519 : _GEN_2031; // @[executor.scala 473:84]
  wire [7:0] _GEN_2524 = mask_2[0] ? byte_512 : _GEN_2032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2525 = mask_2[1] ? byte_513 : _GEN_2033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2526 = mask_2[2] ? byte_514 : _GEN_2034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2527 = mask_2[3] ? byte_515 : _GEN_2035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2528 = _GEN_8594 == 8'h3b ? _GEN_2524 : _GEN_2032; // @[executor.scala 473:84]
  wire [7:0] _GEN_2529 = _GEN_8594 == 8'h3b ? _GEN_2525 : _GEN_2033; // @[executor.scala 473:84]
  wire [7:0] _GEN_2530 = _GEN_8594 == 8'h3b ? _GEN_2526 : _GEN_2034; // @[executor.scala 473:84]
  wire [7:0] _GEN_2531 = _GEN_8594 == 8'h3b ? _GEN_2527 : _GEN_2035; // @[executor.scala 473:84]
  wire [7:0] _GEN_2532 = mask_2[0] ? byte_512 : _GEN_2036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2533 = mask_2[1] ? byte_513 : _GEN_2037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2534 = mask_2[2] ? byte_514 : _GEN_2038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2535 = mask_2[3] ? byte_515 : _GEN_2039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2536 = _GEN_8594 == 8'h3c ? _GEN_2532 : _GEN_2036; // @[executor.scala 473:84]
  wire [7:0] _GEN_2537 = _GEN_8594 == 8'h3c ? _GEN_2533 : _GEN_2037; // @[executor.scala 473:84]
  wire [7:0] _GEN_2538 = _GEN_8594 == 8'h3c ? _GEN_2534 : _GEN_2038; // @[executor.scala 473:84]
  wire [7:0] _GEN_2539 = _GEN_8594 == 8'h3c ? _GEN_2535 : _GEN_2039; // @[executor.scala 473:84]
  wire [7:0] _GEN_2540 = mask_2[0] ? byte_512 : _GEN_2040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2541 = mask_2[1] ? byte_513 : _GEN_2041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2542 = mask_2[2] ? byte_514 : _GEN_2042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2543 = mask_2[3] ? byte_515 : _GEN_2043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2544 = _GEN_8594 == 8'h3d ? _GEN_2540 : _GEN_2040; // @[executor.scala 473:84]
  wire [7:0] _GEN_2545 = _GEN_8594 == 8'h3d ? _GEN_2541 : _GEN_2041; // @[executor.scala 473:84]
  wire [7:0] _GEN_2546 = _GEN_8594 == 8'h3d ? _GEN_2542 : _GEN_2042; // @[executor.scala 473:84]
  wire [7:0] _GEN_2547 = _GEN_8594 == 8'h3d ? _GEN_2543 : _GEN_2043; // @[executor.scala 473:84]
  wire [7:0] _GEN_2548 = mask_2[0] ? byte_512 : _GEN_2044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2549 = mask_2[1] ? byte_513 : _GEN_2045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2550 = mask_2[2] ? byte_514 : _GEN_2046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2551 = mask_2[3] ? byte_515 : _GEN_2047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2552 = _GEN_8594 == 8'h3e ? _GEN_2548 : _GEN_2044; // @[executor.scala 473:84]
  wire [7:0] _GEN_2553 = _GEN_8594 == 8'h3e ? _GEN_2549 : _GEN_2045; // @[executor.scala 473:84]
  wire [7:0] _GEN_2554 = _GEN_8594 == 8'h3e ? _GEN_2550 : _GEN_2046; // @[executor.scala 473:84]
  wire [7:0] _GEN_2555 = _GEN_8594 == 8'h3e ? _GEN_2551 : _GEN_2047; // @[executor.scala 473:84]
  wire [7:0] _GEN_2556 = mask_2[0] ? byte_512 : _GEN_2048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2557 = mask_2[1] ? byte_513 : _GEN_2049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2558 = mask_2[2] ? byte_514 : _GEN_2050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2559 = mask_2[3] ? byte_515 : _GEN_2051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2560 = _GEN_8594 == 8'h3f ? _GEN_2556 : _GEN_2048; // @[executor.scala 473:84]
  wire [7:0] _GEN_2561 = _GEN_8594 == 8'h3f ? _GEN_2557 : _GEN_2049; // @[executor.scala 473:84]
  wire [7:0] _GEN_2562 = _GEN_8594 == 8'h3f ? _GEN_2558 : _GEN_2050; // @[executor.scala 473:84]
  wire [7:0] _GEN_2563 = _GEN_8594 == 8'h3f ? _GEN_2559 : _GEN_2051; // @[executor.scala 473:84]
  wire [7:0] _GEN_2564 = opcode_2 != 4'h0 ? _GEN_2056 : _GEN_1796; // @[executor.scala 470:55]
  wire [7:0] _GEN_2565 = opcode_2 != 4'h0 ? _GEN_2057 : _GEN_1797; // @[executor.scala 470:55]
  wire [7:0] _GEN_2566 = opcode_2 != 4'h0 ? _GEN_2058 : _GEN_1798; // @[executor.scala 470:55]
  wire [7:0] _GEN_2567 = opcode_2 != 4'h0 ? _GEN_2059 : _GEN_1799; // @[executor.scala 470:55]
  wire [7:0] _GEN_2568 = opcode_2 != 4'h0 ? _GEN_2064 : _GEN_1800; // @[executor.scala 470:55]
  wire [7:0] _GEN_2569 = opcode_2 != 4'h0 ? _GEN_2065 : _GEN_1801; // @[executor.scala 470:55]
  wire [7:0] _GEN_2570 = opcode_2 != 4'h0 ? _GEN_2066 : _GEN_1802; // @[executor.scala 470:55]
  wire [7:0] _GEN_2571 = opcode_2 != 4'h0 ? _GEN_2067 : _GEN_1803; // @[executor.scala 470:55]
  wire [7:0] _GEN_2572 = opcode_2 != 4'h0 ? _GEN_2072 : _GEN_1804; // @[executor.scala 470:55]
  wire [7:0] _GEN_2573 = opcode_2 != 4'h0 ? _GEN_2073 : _GEN_1805; // @[executor.scala 470:55]
  wire [7:0] _GEN_2574 = opcode_2 != 4'h0 ? _GEN_2074 : _GEN_1806; // @[executor.scala 470:55]
  wire [7:0] _GEN_2575 = opcode_2 != 4'h0 ? _GEN_2075 : _GEN_1807; // @[executor.scala 470:55]
  wire [7:0] _GEN_2576 = opcode_2 != 4'h0 ? _GEN_2080 : _GEN_1808; // @[executor.scala 470:55]
  wire [7:0] _GEN_2577 = opcode_2 != 4'h0 ? _GEN_2081 : _GEN_1809; // @[executor.scala 470:55]
  wire [7:0] _GEN_2578 = opcode_2 != 4'h0 ? _GEN_2082 : _GEN_1810; // @[executor.scala 470:55]
  wire [7:0] _GEN_2579 = opcode_2 != 4'h0 ? _GEN_2083 : _GEN_1811; // @[executor.scala 470:55]
  wire [7:0] _GEN_2580 = opcode_2 != 4'h0 ? _GEN_2088 : _GEN_1812; // @[executor.scala 470:55]
  wire [7:0] _GEN_2581 = opcode_2 != 4'h0 ? _GEN_2089 : _GEN_1813; // @[executor.scala 470:55]
  wire [7:0] _GEN_2582 = opcode_2 != 4'h0 ? _GEN_2090 : _GEN_1814; // @[executor.scala 470:55]
  wire [7:0] _GEN_2583 = opcode_2 != 4'h0 ? _GEN_2091 : _GEN_1815; // @[executor.scala 470:55]
  wire [7:0] _GEN_2584 = opcode_2 != 4'h0 ? _GEN_2096 : _GEN_1816; // @[executor.scala 470:55]
  wire [7:0] _GEN_2585 = opcode_2 != 4'h0 ? _GEN_2097 : _GEN_1817; // @[executor.scala 470:55]
  wire [7:0] _GEN_2586 = opcode_2 != 4'h0 ? _GEN_2098 : _GEN_1818; // @[executor.scala 470:55]
  wire [7:0] _GEN_2587 = opcode_2 != 4'h0 ? _GEN_2099 : _GEN_1819; // @[executor.scala 470:55]
  wire [7:0] _GEN_2588 = opcode_2 != 4'h0 ? _GEN_2104 : _GEN_1820; // @[executor.scala 470:55]
  wire [7:0] _GEN_2589 = opcode_2 != 4'h0 ? _GEN_2105 : _GEN_1821; // @[executor.scala 470:55]
  wire [7:0] _GEN_2590 = opcode_2 != 4'h0 ? _GEN_2106 : _GEN_1822; // @[executor.scala 470:55]
  wire [7:0] _GEN_2591 = opcode_2 != 4'h0 ? _GEN_2107 : _GEN_1823; // @[executor.scala 470:55]
  wire [7:0] _GEN_2592 = opcode_2 != 4'h0 ? _GEN_2112 : _GEN_1824; // @[executor.scala 470:55]
  wire [7:0] _GEN_2593 = opcode_2 != 4'h0 ? _GEN_2113 : _GEN_1825; // @[executor.scala 470:55]
  wire [7:0] _GEN_2594 = opcode_2 != 4'h0 ? _GEN_2114 : _GEN_1826; // @[executor.scala 470:55]
  wire [7:0] _GEN_2595 = opcode_2 != 4'h0 ? _GEN_2115 : _GEN_1827; // @[executor.scala 470:55]
  wire [7:0] _GEN_2596 = opcode_2 != 4'h0 ? _GEN_2120 : _GEN_1828; // @[executor.scala 470:55]
  wire [7:0] _GEN_2597 = opcode_2 != 4'h0 ? _GEN_2121 : _GEN_1829; // @[executor.scala 470:55]
  wire [7:0] _GEN_2598 = opcode_2 != 4'h0 ? _GEN_2122 : _GEN_1830; // @[executor.scala 470:55]
  wire [7:0] _GEN_2599 = opcode_2 != 4'h0 ? _GEN_2123 : _GEN_1831; // @[executor.scala 470:55]
  wire [7:0] _GEN_2600 = opcode_2 != 4'h0 ? _GEN_2128 : _GEN_1832; // @[executor.scala 470:55]
  wire [7:0] _GEN_2601 = opcode_2 != 4'h0 ? _GEN_2129 : _GEN_1833; // @[executor.scala 470:55]
  wire [7:0] _GEN_2602 = opcode_2 != 4'h0 ? _GEN_2130 : _GEN_1834; // @[executor.scala 470:55]
  wire [7:0] _GEN_2603 = opcode_2 != 4'h0 ? _GEN_2131 : _GEN_1835; // @[executor.scala 470:55]
  wire [7:0] _GEN_2604 = opcode_2 != 4'h0 ? _GEN_2136 : _GEN_1836; // @[executor.scala 470:55]
  wire [7:0] _GEN_2605 = opcode_2 != 4'h0 ? _GEN_2137 : _GEN_1837; // @[executor.scala 470:55]
  wire [7:0] _GEN_2606 = opcode_2 != 4'h0 ? _GEN_2138 : _GEN_1838; // @[executor.scala 470:55]
  wire [7:0] _GEN_2607 = opcode_2 != 4'h0 ? _GEN_2139 : _GEN_1839; // @[executor.scala 470:55]
  wire [7:0] _GEN_2608 = opcode_2 != 4'h0 ? _GEN_2144 : _GEN_1840; // @[executor.scala 470:55]
  wire [7:0] _GEN_2609 = opcode_2 != 4'h0 ? _GEN_2145 : _GEN_1841; // @[executor.scala 470:55]
  wire [7:0] _GEN_2610 = opcode_2 != 4'h0 ? _GEN_2146 : _GEN_1842; // @[executor.scala 470:55]
  wire [7:0] _GEN_2611 = opcode_2 != 4'h0 ? _GEN_2147 : _GEN_1843; // @[executor.scala 470:55]
  wire [7:0] _GEN_2612 = opcode_2 != 4'h0 ? _GEN_2152 : _GEN_1844; // @[executor.scala 470:55]
  wire [7:0] _GEN_2613 = opcode_2 != 4'h0 ? _GEN_2153 : _GEN_1845; // @[executor.scala 470:55]
  wire [7:0] _GEN_2614 = opcode_2 != 4'h0 ? _GEN_2154 : _GEN_1846; // @[executor.scala 470:55]
  wire [7:0] _GEN_2615 = opcode_2 != 4'h0 ? _GEN_2155 : _GEN_1847; // @[executor.scala 470:55]
  wire [7:0] _GEN_2616 = opcode_2 != 4'h0 ? _GEN_2160 : _GEN_1848; // @[executor.scala 470:55]
  wire [7:0] _GEN_2617 = opcode_2 != 4'h0 ? _GEN_2161 : _GEN_1849; // @[executor.scala 470:55]
  wire [7:0] _GEN_2618 = opcode_2 != 4'h0 ? _GEN_2162 : _GEN_1850; // @[executor.scala 470:55]
  wire [7:0] _GEN_2619 = opcode_2 != 4'h0 ? _GEN_2163 : _GEN_1851; // @[executor.scala 470:55]
  wire [7:0] _GEN_2620 = opcode_2 != 4'h0 ? _GEN_2168 : _GEN_1852; // @[executor.scala 470:55]
  wire [7:0] _GEN_2621 = opcode_2 != 4'h0 ? _GEN_2169 : _GEN_1853; // @[executor.scala 470:55]
  wire [7:0] _GEN_2622 = opcode_2 != 4'h0 ? _GEN_2170 : _GEN_1854; // @[executor.scala 470:55]
  wire [7:0] _GEN_2623 = opcode_2 != 4'h0 ? _GEN_2171 : _GEN_1855; // @[executor.scala 470:55]
  wire [7:0] _GEN_2624 = opcode_2 != 4'h0 ? _GEN_2176 : _GEN_1856; // @[executor.scala 470:55]
  wire [7:0] _GEN_2625 = opcode_2 != 4'h0 ? _GEN_2177 : _GEN_1857; // @[executor.scala 470:55]
  wire [7:0] _GEN_2626 = opcode_2 != 4'h0 ? _GEN_2178 : _GEN_1858; // @[executor.scala 470:55]
  wire [7:0] _GEN_2627 = opcode_2 != 4'h0 ? _GEN_2179 : _GEN_1859; // @[executor.scala 470:55]
  wire [7:0] _GEN_2628 = opcode_2 != 4'h0 ? _GEN_2184 : _GEN_1860; // @[executor.scala 470:55]
  wire [7:0] _GEN_2629 = opcode_2 != 4'h0 ? _GEN_2185 : _GEN_1861; // @[executor.scala 470:55]
  wire [7:0] _GEN_2630 = opcode_2 != 4'h0 ? _GEN_2186 : _GEN_1862; // @[executor.scala 470:55]
  wire [7:0] _GEN_2631 = opcode_2 != 4'h0 ? _GEN_2187 : _GEN_1863; // @[executor.scala 470:55]
  wire [7:0] _GEN_2632 = opcode_2 != 4'h0 ? _GEN_2192 : _GEN_1864; // @[executor.scala 470:55]
  wire [7:0] _GEN_2633 = opcode_2 != 4'h0 ? _GEN_2193 : _GEN_1865; // @[executor.scala 470:55]
  wire [7:0] _GEN_2634 = opcode_2 != 4'h0 ? _GEN_2194 : _GEN_1866; // @[executor.scala 470:55]
  wire [7:0] _GEN_2635 = opcode_2 != 4'h0 ? _GEN_2195 : _GEN_1867; // @[executor.scala 470:55]
  wire [7:0] _GEN_2636 = opcode_2 != 4'h0 ? _GEN_2200 : _GEN_1868; // @[executor.scala 470:55]
  wire [7:0] _GEN_2637 = opcode_2 != 4'h0 ? _GEN_2201 : _GEN_1869; // @[executor.scala 470:55]
  wire [7:0] _GEN_2638 = opcode_2 != 4'h0 ? _GEN_2202 : _GEN_1870; // @[executor.scala 470:55]
  wire [7:0] _GEN_2639 = opcode_2 != 4'h0 ? _GEN_2203 : _GEN_1871; // @[executor.scala 470:55]
  wire [7:0] _GEN_2640 = opcode_2 != 4'h0 ? _GEN_2208 : _GEN_1872; // @[executor.scala 470:55]
  wire [7:0] _GEN_2641 = opcode_2 != 4'h0 ? _GEN_2209 : _GEN_1873; // @[executor.scala 470:55]
  wire [7:0] _GEN_2642 = opcode_2 != 4'h0 ? _GEN_2210 : _GEN_1874; // @[executor.scala 470:55]
  wire [7:0] _GEN_2643 = opcode_2 != 4'h0 ? _GEN_2211 : _GEN_1875; // @[executor.scala 470:55]
  wire [7:0] _GEN_2644 = opcode_2 != 4'h0 ? _GEN_2216 : _GEN_1876; // @[executor.scala 470:55]
  wire [7:0] _GEN_2645 = opcode_2 != 4'h0 ? _GEN_2217 : _GEN_1877; // @[executor.scala 470:55]
  wire [7:0] _GEN_2646 = opcode_2 != 4'h0 ? _GEN_2218 : _GEN_1878; // @[executor.scala 470:55]
  wire [7:0] _GEN_2647 = opcode_2 != 4'h0 ? _GEN_2219 : _GEN_1879; // @[executor.scala 470:55]
  wire [7:0] _GEN_2648 = opcode_2 != 4'h0 ? _GEN_2224 : _GEN_1880; // @[executor.scala 470:55]
  wire [7:0] _GEN_2649 = opcode_2 != 4'h0 ? _GEN_2225 : _GEN_1881; // @[executor.scala 470:55]
  wire [7:0] _GEN_2650 = opcode_2 != 4'h0 ? _GEN_2226 : _GEN_1882; // @[executor.scala 470:55]
  wire [7:0] _GEN_2651 = opcode_2 != 4'h0 ? _GEN_2227 : _GEN_1883; // @[executor.scala 470:55]
  wire [7:0] _GEN_2652 = opcode_2 != 4'h0 ? _GEN_2232 : _GEN_1884; // @[executor.scala 470:55]
  wire [7:0] _GEN_2653 = opcode_2 != 4'h0 ? _GEN_2233 : _GEN_1885; // @[executor.scala 470:55]
  wire [7:0] _GEN_2654 = opcode_2 != 4'h0 ? _GEN_2234 : _GEN_1886; // @[executor.scala 470:55]
  wire [7:0] _GEN_2655 = opcode_2 != 4'h0 ? _GEN_2235 : _GEN_1887; // @[executor.scala 470:55]
  wire [7:0] _GEN_2656 = opcode_2 != 4'h0 ? _GEN_2240 : _GEN_1888; // @[executor.scala 470:55]
  wire [7:0] _GEN_2657 = opcode_2 != 4'h0 ? _GEN_2241 : _GEN_1889; // @[executor.scala 470:55]
  wire [7:0] _GEN_2658 = opcode_2 != 4'h0 ? _GEN_2242 : _GEN_1890; // @[executor.scala 470:55]
  wire [7:0] _GEN_2659 = opcode_2 != 4'h0 ? _GEN_2243 : _GEN_1891; // @[executor.scala 470:55]
  wire [7:0] _GEN_2660 = opcode_2 != 4'h0 ? _GEN_2248 : _GEN_1892; // @[executor.scala 470:55]
  wire [7:0] _GEN_2661 = opcode_2 != 4'h0 ? _GEN_2249 : _GEN_1893; // @[executor.scala 470:55]
  wire [7:0] _GEN_2662 = opcode_2 != 4'h0 ? _GEN_2250 : _GEN_1894; // @[executor.scala 470:55]
  wire [7:0] _GEN_2663 = opcode_2 != 4'h0 ? _GEN_2251 : _GEN_1895; // @[executor.scala 470:55]
  wire [7:0] _GEN_2664 = opcode_2 != 4'h0 ? _GEN_2256 : _GEN_1896; // @[executor.scala 470:55]
  wire [7:0] _GEN_2665 = opcode_2 != 4'h0 ? _GEN_2257 : _GEN_1897; // @[executor.scala 470:55]
  wire [7:0] _GEN_2666 = opcode_2 != 4'h0 ? _GEN_2258 : _GEN_1898; // @[executor.scala 470:55]
  wire [7:0] _GEN_2667 = opcode_2 != 4'h0 ? _GEN_2259 : _GEN_1899; // @[executor.scala 470:55]
  wire [7:0] _GEN_2668 = opcode_2 != 4'h0 ? _GEN_2264 : _GEN_1900; // @[executor.scala 470:55]
  wire [7:0] _GEN_2669 = opcode_2 != 4'h0 ? _GEN_2265 : _GEN_1901; // @[executor.scala 470:55]
  wire [7:0] _GEN_2670 = opcode_2 != 4'h0 ? _GEN_2266 : _GEN_1902; // @[executor.scala 470:55]
  wire [7:0] _GEN_2671 = opcode_2 != 4'h0 ? _GEN_2267 : _GEN_1903; // @[executor.scala 470:55]
  wire [7:0] _GEN_2672 = opcode_2 != 4'h0 ? _GEN_2272 : _GEN_1904; // @[executor.scala 470:55]
  wire [7:0] _GEN_2673 = opcode_2 != 4'h0 ? _GEN_2273 : _GEN_1905; // @[executor.scala 470:55]
  wire [7:0] _GEN_2674 = opcode_2 != 4'h0 ? _GEN_2274 : _GEN_1906; // @[executor.scala 470:55]
  wire [7:0] _GEN_2675 = opcode_2 != 4'h0 ? _GEN_2275 : _GEN_1907; // @[executor.scala 470:55]
  wire [7:0] _GEN_2676 = opcode_2 != 4'h0 ? _GEN_2280 : _GEN_1908; // @[executor.scala 470:55]
  wire [7:0] _GEN_2677 = opcode_2 != 4'h0 ? _GEN_2281 : _GEN_1909; // @[executor.scala 470:55]
  wire [7:0] _GEN_2678 = opcode_2 != 4'h0 ? _GEN_2282 : _GEN_1910; // @[executor.scala 470:55]
  wire [7:0] _GEN_2679 = opcode_2 != 4'h0 ? _GEN_2283 : _GEN_1911; // @[executor.scala 470:55]
  wire [7:0] _GEN_2680 = opcode_2 != 4'h0 ? _GEN_2288 : _GEN_1912; // @[executor.scala 470:55]
  wire [7:0] _GEN_2681 = opcode_2 != 4'h0 ? _GEN_2289 : _GEN_1913; // @[executor.scala 470:55]
  wire [7:0] _GEN_2682 = opcode_2 != 4'h0 ? _GEN_2290 : _GEN_1914; // @[executor.scala 470:55]
  wire [7:0] _GEN_2683 = opcode_2 != 4'h0 ? _GEN_2291 : _GEN_1915; // @[executor.scala 470:55]
  wire [7:0] _GEN_2684 = opcode_2 != 4'h0 ? _GEN_2296 : _GEN_1916; // @[executor.scala 470:55]
  wire [7:0] _GEN_2685 = opcode_2 != 4'h0 ? _GEN_2297 : _GEN_1917; // @[executor.scala 470:55]
  wire [7:0] _GEN_2686 = opcode_2 != 4'h0 ? _GEN_2298 : _GEN_1918; // @[executor.scala 470:55]
  wire [7:0] _GEN_2687 = opcode_2 != 4'h0 ? _GEN_2299 : _GEN_1919; // @[executor.scala 470:55]
  wire [7:0] _GEN_2688 = opcode_2 != 4'h0 ? _GEN_2304 : _GEN_1920; // @[executor.scala 470:55]
  wire [7:0] _GEN_2689 = opcode_2 != 4'h0 ? _GEN_2305 : _GEN_1921; // @[executor.scala 470:55]
  wire [7:0] _GEN_2690 = opcode_2 != 4'h0 ? _GEN_2306 : _GEN_1922; // @[executor.scala 470:55]
  wire [7:0] _GEN_2691 = opcode_2 != 4'h0 ? _GEN_2307 : _GEN_1923; // @[executor.scala 470:55]
  wire [7:0] _GEN_2692 = opcode_2 != 4'h0 ? _GEN_2312 : _GEN_1924; // @[executor.scala 470:55]
  wire [7:0] _GEN_2693 = opcode_2 != 4'h0 ? _GEN_2313 : _GEN_1925; // @[executor.scala 470:55]
  wire [7:0] _GEN_2694 = opcode_2 != 4'h0 ? _GEN_2314 : _GEN_1926; // @[executor.scala 470:55]
  wire [7:0] _GEN_2695 = opcode_2 != 4'h0 ? _GEN_2315 : _GEN_1927; // @[executor.scala 470:55]
  wire [7:0] _GEN_2696 = opcode_2 != 4'h0 ? _GEN_2320 : _GEN_1928; // @[executor.scala 470:55]
  wire [7:0] _GEN_2697 = opcode_2 != 4'h0 ? _GEN_2321 : _GEN_1929; // @[executor.scala 470:55]
  wire [7:0] _GEN_2698 = opcode_2 != 4'h0 ? _GEN_2322 : _GEN_1930; // @[executor.scala 470:55]
  wire [7:0] _GEN_2699 = opcode_2 != 4'h0 ? _GEN_2323 : _GEN_1931; // @[executor.scala 470:55]
  wire [7:0] _GEN_2700 = opcode_2 != 4'h0 ? _GEN_2328 : _GEN_1932; // @[executor.scala 470:55]
  wire [7:0] _GEN_2701 = opcode_2 != 4'h0 ? _GEN_2329 : _GEN_1933; // @[executor.scala 470:55]
  wire [7:0] _GEN_2702 = opcode_2 != 4'h0 ? _GEN_2330 : _GEN_1934; // @[executor.scala 470:55]
  wire [7:0] _GEN_2703 = opcode_2 != 4'h0 ? _GEN_2331 : _GEN_1935; // @[executor.scala 470:55]
  wire [7:0] _GEN_2704 = opcode_2 != 4'h0 ? _GEN_2336 : _GEN_1936; // @[executor.scala 470:55]
  wire [7:0] _GEN_2705 = opcode_2 != 4'h0 ? _GEN_2337 : _GEN_1937; // @[executor.scala 470:55]
  wire [7:0] _GEN_2706 = opcode_2 != 4'h0 ? _GEN_2338 : _GEN_1938; // @[executor.scala 470:55]
  wire [7:0] _GEN_2707 = opcode_2 != 4'h0 ? _GEN_2339 : _GEN_1939; // @[executor.scala 470:55]
  wire [7:0] _GEN_2708 = opcode_2 != 4'h0 ? _GEN_2344 : _GEN_1940; // @[executor.scala 470:55]
  wire [7:0] _GEN_2709 = opcode_2 != 4'h0 ? _GEN_2345 : _GEN_1941; // @[executor.scala 470:55]
  wire [7:0] _GEN_2710 = opcode_2 != 4'h0 ? _GEN_2346 : _GEN_1942; // @[executor.scala 470:55]
  wire [7:0] _GEN_2711 = opcode_2 != 4'h0 ? _GEN_2347 : _GEN_1943; // @[executor.scala 470:55]
  wire [7:0] _GEN_2712 = opcode_2 != 4'h0 ? _GEN_2352 : _GEN_1944; // @[executor.scala 470:55]
  wire [7:0] _GEN_2713 = opcode_2 != 4'h0 ? _GEN_2353 : _GEN_1945; // @[executor.scala 470:55]
  wire [7:0] _GEN_2714 = opcode_2 != 4'h0 ? _GEN_2354 : _GEN_1946; // @[executor.scala 470:55]
  wire [7:0] _GEN_2715 = opcode_2 != 4'h0 ? _GEN_2355 : _GEN_1947; // @[executor.scala 470:55]
  wire [7:0] _GEN_2716 = opcode_2 != 4'h0 ? _GEN_2360 : _GEN_1948; // @[executor.scala 470:55]
  wire [7:0] _GEN_2717 = opcode_2 != 4'h0 ? _GEN_2361 : _GEN_1949; // @[executor.scala 470:55]
  wire [7:0] _GEN_2718 = opcode_2 != 4'h0 ? _GEN_2362 : _GEN_1950; // @[executor.scala 470:55]
  wire [7:0] _GEN_2719 = opcode_2 != 4'h0 ? _GEN_2363 : _GEN_1951; // @[executor.scala 470:55]
  wire [7:0] _GEN_2720 = opcode_2 != 4'h0 ? _GEN_2368 : _GEN_1952; // @[executor.scala 470:55]
  wire [7:0] _GEN_2721 = opcode_2 != 4'h0 ? _GEN_2369 : _GEN_1953; // @[executor.scala 470:55]
  wire [7:0] _GEN_2722 = opcode_2 != 4'h0 ? _GEN_2370 : _GEN_1954; // @[executor.scala 470:55]
  wire [7:0] _GEN_2723 = opcode_2 != 4'h0 ? _GEN_2371 : _GEN_1955; // @[executor.scala 470:55]
  wire [7:0] _GEN_2724 = opcode_2 != 4'h0 ? _GEN_2376 : _GEN_1956; // @[executor.scala 470:55]
  wire [7:0] _GEN_2725 = opcode_2 != 4'h0 ? _GEN_2377 : _GEN_1957; // @[executor.scala 470:55]
  wire [7:0] _GEN_2726 = opcode_2 != 4'h0 ? _GEN_2378 : _GEN_1958; // @[executor.scala 470:55]
  wire [7:0] _GEN_2727 = opcode_2 != 4'h0 ? _GEN_2379 : _GEN_1959; // @[executor.scala 470:55]
  wire [7:0] _GEN_2728 = opcode_2 != 4'h0 ? _GEN_2384 : _GEN_1960; // @[executor.scala 470:55]
  wire [7:0] _GEN_2729 = opcode_2 != 4'h0 ? _GEN_2385 : _GEN_1961; // @[executor.scala 470:55]
  wire [7:0] _GEN_2730 = opcode_2 != 4'h0 ? _GEN_2386 : _GEN_1962; // @[executor.scala 470:55]
  wire [7:0] _GEN_2731 = opcode_2 != 4'h0 ? _GEN_2387 : _GEN_1963; // @[executor.scala 470:55]
  wire [7:0] _GEN_2732 = opcode_2 != 4'h0 ? _GEN_2392 : _GEN_1964; // @[executor.scala 470:55]
  wire [7:0] _GEN_2733 = opcode_2 != 4'h0 ? _GEN_2393 : _GEN_1965; // @[executor.scala 470:55]
  wire [7:0] _GEN_2734 = opcode_2 != 4'h0 ? _GEN_2394 : _GEN_1966; // @[executor.scala 470:55]
  wire [7:0] _GEN_2735 = opcode_2 != 4'h0 ? _GEN_2395 : _GEN_1967; // @[executor.scala 470:55]
  wire [7:0] _GEN_2736 = opcode_2 != 4'h0 ? _GEN_2400 : _GEN_1968; // @[executor.scala 470:55]
  wire [7:0] _GEN_2737 = opcode_2 != 4'h0 ? _GEN_2401 : _GEN_1969; // @[executor.scala 470:55]
  wire [7:0] _GEN_2738 = opcode_2 != 4'h0 ? _GEN_2402 : _GEN_1970; // @[executor.scala 470:55]
  wire [7:0] _GEN_2739 = opcode_2 != 4'h0 ? _GEN_2403 : _GEN_1971; // @[executor.scala 470:55]
  wire [7:0] _GEN_2740 = opcode_2 != 4'h0 ? _GEN_2408 : _GEN_1972; // @[executor.scala 470:55]
  wire [7:0] _GEN_2741 = opcode_2 != 4'h0 ? _GEN_2409 : _GEN_1973; // @[executor.scala 470:55]
  wire [7:0] _GEN_2742 = opcode_2 != 4'h0 ? _GEN_2410 : _GEN_1974; // @[executor.scala 470:55]
  wire [7:0] _GEN_2743 = opcode_2 != 4'h0 ? _GEN_2411 : _GEN_1975; // @[executor.scala 470:55]
  wire [7:0] _GEN_2744 = opcode_2 != 4'h0 ? _GEN_2416 : _GEN_1976; // @[executor.scala 470:55]
  wire [7:0] _GEN_2745 = opcode_2 != 4'h0 ? _GEN_2417 : _GEN_1977; // @[executor.scala 470:55]
  wire [7:0] _GEN_2746 = opcode_2 != 4'h0 ? _GEN_2418 : _GEN_1978; // @[executor.scala 470:55]
  wire [7:0] _GEN_2747 = opcode_2 != 4'h0 ? _GEN_2419 : _GEN_1979; // @[executor.scala 470:55]
  wire [7:0] _GEN_2748 = opcode_2 != 4'h0 ? _GEN_2424 : _GEN_1980; // @[executor.scala 470:55]
  wire [7:0] _GEN_2749 = opcode_2 != 4'h0 ? _GEN_2425 : _GEN_1981; // @[executor.scala 470:55]
  wire [7:0] _GEN_2750 = opcode_2 != 4'h0 ? _GEN_2426 : _GEN_1982; // @[executor.scala 470:55]
  wire [7:0] _GEN_2751 = opcode_2 != 4'h0 ? _GEN_2427 : _GEN_1983; // @[executor.scala 470:55]
  wire [7:0] _GEN_2752 = opcode_2 != 4'h0 ? _GEN_2432 : _GEN_1984; // @[executor.scala 470:55]
  wire [7:0] _GEN_2753 = opcode_2 != 4'h0 ? _GEN_2433 : _GEN_1985; // @[executor.scala 470:55]
  wire [7:0] _GEN_2754 = opcode_2 != 4'h0 ? _GEN_2434 : _GEN_1986; // @[executor.scala 470:55]
  wire [7:0] _GEN_2755 = opcode_2 != 4'h0 ? _GEN_2435 : _GEN_1987; // @[executor.scala 470:55]
  wire [7:0] _GEN_2756 = opcode_2 != 4'h0 ? _GEN_2440 : _GEN_1988; // @[executor.scala 470:55]
  wire [7:0] _GEN_2757 = opcode_2 != 4'h0 ? _GEN_2441 : _GEN_1989; // @[executor.scala 470:55]
  wire [7:0] _GEN_2758 = opcode_2 != 4'h0 ? _GEN_2442 : _GEN_1990; // @[executor.scala 470:55]
  wire [7:0] _GEN_2759 = opcode_2 != 4'h0 ? _GEN_2443 : _GEN_1991; // @[executor.scala 470:55]
  wire [7:0] _GEN_2760 = opcode_2 != 4'h0 ? _GEN_2448 : _GEN_1992; // @[executor.scala 470:55]
  wire [7:0] _GEN_2761 = opcode_2 != 4'h0 ? _GEN_2449 : _GEN_1993; // @[executor.scala 470:55]
  wire [7:0] _GEN_2762 = opcode_2 != 4'h0 ? _GEN_2450 : _GEN_1994; // @[executor.scala 470:55]
  wire [7:0] _GEN_2763 = opcode_2 != 4'h0 ? _GEN_2451 : _GEN_1995; // @[executor.scala 470:55]
  wire [7:0] _GEN_2764 = opcode_2 != 4'h0 ? _GEN_2456 : _GEN_1996; // @[executor.scala 470:55]
  wire [7:0] _GEN_2765 = opcode_2 != 4'h0 ? _GEN_2457 : _GEN_1997; // @[executor.scala 470:55]
  wire [7:0] _GEN_2766 = opcode_2 != 4'h0 ? _GEN_2458 : _GEN_1998; // @[executor.scala 470:55]
  wire [7:0] _GEN_2767 = opcode_2 != 4'h0 ? _GEN_2459 : _GEN_1999; // @[executor.scala 470:55]
  wire [7:0] _GEN_2768 = opcode_2 != 4'h0 ? _GEN_2464 : _GEN_2000; // @[executor.scala 470:55]
  wire [7:0] _GEN_2769 = opcode_2 != 4'h0 ? _GEN_2465 : _GEN_2001; // @[executor.scala 470:55]
  wire [7:0] _GEN_2770 = opcode_2 != 4'h0 ? _GEN_2466 : _GEN_2002; // @[executor.scala 470:55]
  wire [7:0] _GEN_2771 = opcode_2 != 4'h0 ? _GEN_2467 : _GEN_2003; // @[executor.scala 470:55]
  wire [7:0] _GEN_2772 = opcode_2 != 4'h0 ? _GEN_2472 : _GEN_2004; // @[executor.scala 470:55]
  wire [7:0] _GEN_2773 = opcode_2 != 4'h0 ? _GEN_2473 : _GEN_2005; // @[executor.scala 470:55]
  wire [7:0] _GEN_2774 = opcode_2 != 4'h0 ? _GEN_2474 : _GEN_2006; // @[executor.scala 470:55]
  wire [7:0] _GEN_2775 = opcode_2 != 4'h0 ? _GEN_2475 : _GEN_2007; // @[executor.scala 470:55]
  wire [7:0] _GEN_2776 = opcode_2 != 4'h0 ? _GEN_2480 : _GEN_2008; // @[executor.scala 470:55]
  wire [7:0] _GEN_2777 = opcode_2 != 4'h0 ? _GEN_2481 : _GEN_2009; // @[executor.scala 470:55]
  wire [7:0] _GEN_2778 = opcode_2 != 4'h0 ? _GEN_2482 : _GEN_2010; // @[executor.scala 470:55]
  wire [7:0] _GEN_2779 = opcode_2 != 4'h0 ? _GEN_2483 : _GEN_2011; // @[executor.scala 470:55]
  wire [7:0] _GEN_2780 = opcode_2 != 4'h0 ? _GEN_2488 : _GEN_2012; // @[executor.scala 470:55]
  wire [7:0] _GEN_2781 = opcode_2 != 4'h0 ? _GEN_2489 : _GEN_2013; // @[executor.scala 470:55]
  wire [7:0] _GEN_2782 = opcode_2 != 4'h0 ? _GEN_2490 : _GEN_2014; // @[executor.scala 470:55]
  wire [7:0] _GEN_2783 = opcode_2 != 4'h0 ? _GEN_2491 : _GEN_2015; // @[executor.scala 470:55]
  wire [7:0] _GEN_2784 = opcode_2 != 4'h0 ? _GEN_2496 : _GEN_2016; // @[executor.scala 470:55]
  wire [7:0] _GEN_2785 = opcode_2 != 4'h0 ? _GEN_2497 : _GEN_2017; // @[executor.scala 470:55]
  wire [7:0] _GEN_2786 = opcode_2 != 4'h0 ? _GEN_2498 : _GEN_2018; // @[executor.scala 470:55]
  wire [7:0] _GEN_2787 = opcode_2 != 4'h0 ? _GEN_2499 : _GEN_2019; // @[executor.scala 470:55]
  wire [7:0] _GEN_2788 = opcode_2 != 4'h0 ? _GEN_2504 : _GEN_2020; // @[executor.scala 470:55]
  wire [7:0] _GEN_2789 = opcode_2 != 4'h0 ? _GEN_2505 : _GEN_2021; // @[executor.scala 470:55]
  wire [7:0] _GEN_2790 = opcode_2 != 4'h0 ? _GEN_2506 : _GEN_2022; // @[executor.scala 470:55]
  wire [7:0] _GEN_2791 = opcode_2 != 4'h0 ? _GEN_2507 : _GEN_2023; // @[executor.scala 470:55]
  wire [7:0] _GEN_2792 = opcode_2 != 4'h0 ? _GEN_2512 : _GEN_2024; // @[executor.scala 470:55]
  wire [7:0] _GEN_2793 = opcode_2 != 4'h0 ? _GEN_2513 : _GEN_2025; // @[executor.scala 470:55]
  wire [7:0] _GEN_2794 = opcode_2 != 4'h0 ? _GEN_2514 : _GEN_2026; // @[executor.scala 470:55]
  wire [7:0] _GEN_2795 = opcode_2 != 4'h0 ? _GEN_2515 : _GEN_2027; // @[executor.scala 470:55]
  wire [7:0] _GEN_2796 = opcode_2 != 4'h0 ? _GEN_2520 : _GEN_2028; // @[executor.scala 470:55]
  wire [7:0] _GEN_2797 = opcode_2 != 4'h0 ? _GEN_2521 : _GEN_2029; // @[executor.scala 470:55]
  wire [7:0] _GEN_2798 = opcode_2 != 4'h0 ? _GEN_2522 : _GEN_2030; // @[executor.scala 470:55]
  wire [7:0] _GEN_2799 = opcode_2 != 4'h0 ? _GEN_2523 : _GEN_2031; // @[executor.scala 470:55]
  wire [7:0] _GEN_2800 = opcode_2 != 4'h0 ? _GEN_2528 : _GEN_2032; // @[executor.scala 470:55]
  wire [7:0] _GEN_2801 = opcode_2 != 4'h0 ? _GEN_2529 : _GEN_2033; // @[executor.scala 470:55]
  wire [7:0] _GEN_2802 = opcode_2 != 4'h0 ? _GEN_2530 : _GEN_2034; // @[executor.scala 470:55]
  wire [7:0] _GEN_2803 = opcode_2 != 4'h0 ? _GEN_2531 : _GEN_2035; // @[executor.scala 470:55]
  wire [7:0] _GEN_2804 = opcode_2 != 4'h0 ? _GEN_2536 : _GEN_2036; // @[executor.scala 470:55]
  wire [7:0] _GEN_2805 = opcode_2 != 4'h0 ? _GEN_2537 : _GEN_2037; // @[executor.scala 470:55]
  wire [7:0] _GEN_2806 = opcode_2 != 4'h0 ? _GEN_2538 : _GEN_2038; // @[executor.scala 470:55]
  wire [7:0] _GEN_2807 = opcode_2 != 4'h0 ? _GEN_2539 : _GEN_2039; // @[executor.scala 470:55]
  wire [7:0] _GEN_2808 = opcode_2 != 4'h0 ? _GEN_2544 : _GEN_2040; // @[executor.scala 470:55]
  wire [7:0] _GEN_2809 = opcode_2 != 4'h0 ? _GEN_2545 : _GEN_2041; // @[executor.scala 470:55]
  wire [7:0] _GEN_2810 = opcode_2 != 4'h0 ? _GEN_2546 : _GEN_2042; // @[executor.scala 470:55]
  wire [7:0] _GEN_2811 = opcode_2 != 4'h0 ? _GEN_2547 : _GEN_2043; // @[executor.scala 470:55]
  wire [7:0] _GEN_2812 = opcode_2 != 4'h0 ? _GEN_2552 : _GEN_2044; // @[executor.scala 470:55]
  wire [7:0] _GEN_2813 = opcode_2 != 4'h0 ? _GEN_2553 : _GEN_2045; // @[executor.scala 470:55]
  wire [7:0] _GEN_2814 = opcode_2 != 4'h0 ? _GEN_2554 : _GEN_2046; // @[executor.scala 470:55]
  wire [7:0] _GEN_2815 = opcode_2 != 4'h0 ? _GEN_2555 : _GEN_2047; // @[executor.scala 470:55]
  wire [7:0] _GEN_2816 = opcode_2 != 4'h0 ? _GEN_2560 : _GEN_2048; // @[executor.scala 470:55]
  wire [7:0] _GEN_2817 = opcode_2 != 4'h0 ? _GEN_2561 : _GEN_2049; // @[executor.scala 470:55]
  wire [7:0] _GEN_2818 = opcode_2 != 4'h0 ? _GEN_2562 : _GEN_2050; // @[executor.scala 470:55]
  wire [7:0] _GEN_2819 = opcode_2 != 4'h0 ? _GEN_2563 : _GEN_2051; // @[executor.scala 470:55]
  wire [3:0] _GEN_2820 = opcode_2 == 4'hf ? parameter_2_2[13:10] : _GEN_1794; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_2821 = opcode_2 == 4'hf ? parameter_2_2[0] : _GEN_1795; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_2822 = opcode_2 == 4'hf ? _GEN_1796 : _GEN_2564; // @[executor.scala 466:52]
  wire [7:0] _GEN_2823 = opcode_2 == 4'hf ? _GEN_1797 : _GEN_2565; // @[executor.scala 466:52]
  wire [7:0] _GEN_2824 = opcode_2 == 4'hf ? _GEN_1798 : _GEN_2566; // @[executor.scala 466:52]
  wire [7:0] _GEN_2825 = opcode_2 == 4'hf ? _GEN_1799 : _GEN_2567; // @[executor.scala 466:52]
  wire [7:0] _GEN_2826 = opcode_2 == 4'hf ? _GEN_1800 : _GEN_2568; // @[executor.scala 466:52]
  wire [7:0] _GEN_2827 = opcode_2 == 4'hf ? _GEN_1801 : _GEN_2569; // @[executor.scala 466:52]
  wire [7:0] _GEN_2828 = opcode_2 == 4'hf ? _GEN_1802 : _GEN_2570; // @[executor.scala 466:52]
  wire [7:0] _GEN_2829 = opcode_2 == 4'hf ? _GEN_1803 : _GEN_2571; // @[executor.scala 466:52]
  wire [7:0] _GEN_2830 = opcode_2 == 4'hf ? _GEN_1804 : _GEN_2572; // @[executor.scala 466:52]
  wire [7:0] _GEN_2831 = opcode_2 == 4'hf ? _GEN_1805 : _GEN_2573; // @[executor.scala 466:52]
  wire [7:0] _GEN_2832 = opcode_2 == 4'hf ? _GEN_1806 : _GEN_2574; // @[executor.scala 466:52]
  wire [7:0] _GEN_2833 = opcode_2 == 4'hf ? _GEN_1807 : _GEN_2575; // @[executor.scala 466:52]
  wire [7:0] _GEN_2834 = opcode_2 == 4'hf ? _GEN_1808 : _GEN_2576; // @[executor.scala 466:52]
  wire [7:0] _GEN_2835 = opcode_2 == 4'hf ? _GEN_1809 : _GEN_2577; // @[executor.scala 466:52]
  wire [7:0] _GEN_2836 = opcode_2 == 4'hf ? _GEN_1810 : _GEN_2578; // @[executor.scala 466:52]
  wire [7:0] _GEN_2837 = opcode_2 == 4'hf ? _GEN_1811 : _GEN_2579; // @[executor.scala 466:52]
  wire [7:0] _GEN_2838 = opcode_2 == 4'hf ? _GEN_1812 : _GEN_2580; // @[executor.scala 466:52]
  wire [7:0] _GEN_2839 = opcode_2 == 4'hf ? _GEN_1813 : _GEN_2581; // @[executor.scala 466:52]
  wire [7:0] _GEN_2840 = opcode_2 == 4'hf ? _GEN_1814 : _GEN_2582; // @[executor.scala 466:52]
  wire [7:0] _GEN_2841 = opcode_2 == 4'hf ? _GEN_1815 : _GEN_2583; // @[executor.scala 466:52]
  wire [7:0] _GEN_2842 = opcode_2 == 4'hf ? _GEN_1816 : _GEN_2584; // @[executor.scala 466:52]
  wire [7:0] _GEN_2843 = opcode_2 == 4'hf ? _GEN_1817 : _GEN_2585; // @[executor.scala 466:52]
  wire [7:0] _GEN_2844 = opcode_2 == 4'hf ? _GEN_1818 : _GEN_2586; // @[executor.scala 466:52]
  wire [7:0] _GEN_2845 = opcode_2 == 4'hf ? _GEN_1819 : _GEN_2587; // @[executor.scala 466:52]
  wire [7:0] _GEN_2846 = opcode_2 == 4'hf ? _GEN_1820 : _GEN_2588; // @[executor.scala 466:52]
  wire [7:0] _GEN_2847 = opcode_2 == 4'hf ? _GEN_1821 : _GEN_2589; // @[executor.scala 466:52]
  wire [7:0] _GEN_2848 = opcode_2 == 4'hf ? _GEN_1822 : _GEN_2590; // @[executor.scala 466:52]
  wire [7:0] _GEN_2849 = opcode_2 == 4'hf ? _GEN_1823 : _GEN_2591; // @[executor.scala 466:52]
  wire [7:0] _GEN_2850 = opcode_2 == 4'hf ? _GEN_1824 : _GEN_2592; // @[executor.scala 466:52]
  wire [7:0] _GEN_2851 = opcode_2 == 4'hf ? _GEN_1825 : _GEN_2593; // @[executor.scala 466:52]
  wire [7:0] _GEN_2852 = opcode_2 == 4'hf ? _GEN_1826 : _GEN_2594; // @[executor.scala 466:52]
  wire [7:0] _GEN_2853 = opcode_2 == 4'hf ? _GEN_1827 : _GEN_2595; // @[executor.scala 466:52]
  wire [7:0] _GEN_2854 = opcode_2 == 4'hf ? _GEN_1828 : _GEN_2596; // @[executor.scala 466:52]
  wire [7:0] _GEN_2855 = opcode_2 == 4'hf ? _GEN_1829 : _GEN_2597; // @[executor.scala 466:52]
  wire [7:0] _GEN_2856 = opcode_2 == 4'hf ? _GEN_1830 : _GEN_2598; // @[executor.scala 466:52]
  wire [7:0] _GEN_2857 = opcode_2 == 4'hf ? _GEN_1831 : _GEN_2599; // @[executor.scala 466:52]
  wire [7:0] _GEN_2858 = opcode_2 == 4'hf ? _GEN_1832 : _GEN_2600; // @[executor.scala 466:52]
  wire [7:0] _GEN_2859 = opcode_2 == 4'hf ? _GEN_1833 : _GEN_2601; // @[executor.scala 466:52]
  wire [7:0] _GEN_2860 = opcode_2 == 4'hf ? _GEN_1834 : _GEN_2602; // @[executor.scala 466:52]
  wire [7:0] _GEN_2861 = opcode_2 == 4'hf ? _GEN_1835 : _GEN_2603; // @[executor.scala 466:52]
  wire [7:0] _GEN_2862 = opcode_2 == 4'hf ? _GEN_1836 : _GEN_2604; // @[executor.scala 466:52]
  wire [7:0] _GEN_2863 = opcode_2 == 4'hf ? _GEN_1837 : _GEN_2605; // @[executor.scala 466:52]
  wire [7:0] _GEN_2864 = opcode_2 == 4'hf ? _GEN_1838 : _GEN_2606; // @[executor.scala 466:52]
  wire [7:0] _GEN_2865 = opcode_2 == 4'hf ? _GEN_1839 : _GEN_2607; // @[executor.scala 466:52]
  wire [7:0] _GEN_2866 = opcode_2 == 4'hf ? _GEN_1840 : _GEN_2608; // @[executor.scala 466:52]
  wire [7:0] _GEN_2867 = opcode_2 == 4'hf ? _GEN_1841 : _GEN_2609; // @[executor.scala 466:52]
  wire [7:0] _GEN_2868 = opcode_2 == 4'hf ? _GEN_1842 : _GEN_2610; // @[executor.scala 466:52]
  wire [7:0] _GEN_2869 = opcode_2 == 4'hf ? _GEN_1843 : _GEN_2611; // @[executor.scala 466:52]
  wire [7:0] _GEN_2870 = opcode_2 == 4'hf ? _GEN_1844 : _GEN_2612; // @[executor.scala 466:52]
  wire [7:0] _GEN_2871 = opcode_2 == 4'hf ? _GEN_1845 : _GEN_2613; // @[executor.scala 466:52]
  wire [7:0] _GEN_2872 = opcode_2 == 4'hf ? _GEN_1846 : _GEN_2614; // @[executor.scala 466:52]
  wire [7:0] _GEN_2873 = opcode_2 == 4'hf ? _GEN_1847 : _GEN_2615; // @[executor.scala 466:52]
  wire [7:0] _GEN_2874 = opcode_2 == 4'hf ? _GEN_1848 : _GEN_2616; // @[executor.scala 466:52]
  wire [7:0] _GEN_2875 = opcode_2 == 4'hf ? _GEN_1849 : _GEN_2617; // @[executor.scala 466:52]
  wire [7:0] _GEN_2876 = opcode_2 == 4'hf ? _GEN_1850 : _GEN_2618; // @[executor.scala 466:52]
  wire [7:0] _GEN_2877 = opcode_2 == 4'hf ? _GEN_1851 : _GEN_2619; // @[executor.scala 466:52]
  wire [7:0] _GEN_2878 = opcode_2 == 4'hf ? _GEN_1852 : _GEN_2620; // @[executor.scala 466:52]
  wire [7:0] _GEN_2879 = opcode_2 == 4'hf ? _GEN_1853 : _GEN_2621; // @[executor.scala 466:52]
  wire [7:0] _GEN_2880 = opcode_2 == 4'hf ? _GEN_1854 : _GEN_2622; // @[executor.scala 466:52]
  wire [7:0] _GEN_2881 = opcode_2 == 4'hf ? _GEN_1855 : _GEN_2623; // @[executor.scala 466:52]
  wire [7:0] _GEN_2882 = opcode_2 == 4'hf ? _GEN_1856 : _GEN_2624; // @[executor.scala 466:52]
  wire [7:0] _GEN_2883 = opcode_2 == 4'hf ? _GEN_1857 : _GEN_2625; // @[executor.scala 466:52]
  wire [7:0] _GEN_2884 = opcode_2 == 4'hf ? _GEN_1858 : _GEN_2626; // @[executor.scala 466:52]
  wire [7:0] _GEN_2885 = opcode_2 == 4'hf ? _GEN_1859 : _GEN_2627; // @[executor.scala 466:52]
  wire [7:0] _GEN_2886 = opcode_2 == 4'hf ? _GEN_1860 : _GEN_2628; // @[executor.scala 466:52]
  wire [7:0] _GEN_2887 = opcode_2 == 4'hf ? _GEN_1861 : _GEN_2629; // @[executor.scala 466:52]
  wire [7:0] _GEN_2888 = opcode_2 == 4'hf ? _GEN_1862 : _GEN_2630; // @[executor.scala 466:52]
  wire [7:0] _GEN_2889 = opcode_2 == 4'hf ? _GEN_1863 : _GEN_2631; // @[executor.scala 466:52]
  wire [7:0] _GEN_2890 = opcode_2 == 4'hf ? _GEN_1864 : _GEN_2632; // @[executor.scala 466:52]
  wire [7:0] _GEN_2891 = opcode_2 == 4'hf ? _GEN_1865 : _GEN_2633; // @[executor.scala 466:52]
  wire [7:0] _GEN_2892 = opcode_2 == 4'hf ? _GEN_1866 : _GEN_2634; // @[executor.scala 466:52]
  wire [7:0] _GEN_2893 = opcode_2 == 4'hf ? _GEN_1867 : _GEN_2635; // @[executor.scala 466:52]
  wire [7:0] _GEN_2894 = opcode_2 == 4'hf ? _GEN_1868 : _GEN_2636; // @[executor.scala 466:52]
  wire [7:0] _GEN_2895 = opcode_2 == 4'hf ? _GEN_1869 : _GEN_2637; // @[executor.scala 466:52]
  wire [7:0] _GEN_2896 = opcode_2 == 4'hf ? _GEN_1870 : _GEN_2638; // @[executor.scala 466:52]
  wire [7:0] _GEN_2897 = opcode_2 == 4'hf ? _GEN_1871 : _GEN_2639; // @[executor.scala 466:52]
  wire [7:0] _GEN_2898 = opcode_2 == 4'hf ? _GEN_1872 : _GEN_2640; // @[executor.scala 466:52]
  wire [7:0] _GEN_2899 = opcode_2 == 4'hf ? _GEN_1873 : _GEN_2641; // @[executor.scala 466:52]
  wire [7:0] _GEN_2900 = opcode_2 == 4'hf ? _GEN_1874 : _GEN_2642; // @[executor.scala 466:52]
  wire [7:0] _GEN_2901 = opcode_2 == 4'hf ? _GEN_1875 : _GEN_2643; // @[executor.scala 466:52]
  wire [7:0] _GEN_2902 = opcode_2 == 4'hf ? _GEN_1876 : _GEN_2644; // @[executor.scala 466:52]
  wire [7:0] _GEN_2903 = opcode_2 == 4'hf ? _GEN_1877 : _GEN_2645; // @[executor.scala 466:52]
  wire [7:0] _GEN_2904 = opcode_2 == 4'hf ? _GEN_1878 : _GEN_2646; // @[executor.scala 466:52]
  wire [7:0] _GEN_2905 = opcode_2 == 4'hf ? _GEN_1879 : _GEN_2647; // @[executor.scala 466:52]
  wire [7:0] _GEN_2906 = opcode_2 == 4'hf ? _GEN_1880 : _GEN_2648; // @[executor.scala 466:52]
  wire [7:0] _GEN_2907 = opcode_2 == 4'hf ? _GEN_1881 : _GEN_2649; // @[executor.scala 466:52]
  wire [7:0] _GEN_2908 = opcode_2 == 4'hf ? _GEN_1882 : _GEN_2650; // @[executor.scala 466:52]
  wire [7:0] _GEN_2909 = opcode_2 == 4'hf ? _GEN_1883 : _GEN_2651; // @[executor.scala 466:52]
  wire [7:0] _GEN_2910 = opcode_2 == 4'hf ? _GEN_1884 : _GEN_2652; // @[executor.scala 466:52]
  wire [7:0] _GEN_2911 = opcode_2 == 4'hf ? _GEN_1885 : _GEN_2653; // @[executor.scala 466:52]
  wire [7:0] _GEN_2912 = opcode_2 == 4'hf ? _GEN_1886 : _GEN_2654; // @[executor.scala 466:52]
  wire [7:0] _GEN_2913 = opcode_2 == 4'hf ? _GEN_1887 : _GEN_2655; // @[executor.scala 466:52]
  wire [7:0] _GEN_2914 = opcode_2 == 4'hf ? _GEN_1888 : _GEN_2656; // @[executor.scala 466:52]
  wire [7:0] _GEN_2915 = opcode_2 == 4'hf ? _GEN_1889 : _GEN_2657; // @[executor.scala 466:52]
  wire [7:0] _GEN_2916 = opcode_2 == 4'hf ? _GEN_1890 : _GEN_2658; // @[executor.scala 466:52]
  wire [7:0] _GEN_2917 = opcode_2 == 4'hf ? _GEN_1891 : _GEN_2659; // @[executor.scala 466:52]
  wire [7:0] _GEN_2918 = opcode_2 == 4'hf ? _GEN_1892 : _GEN_2660; // @[executor.scala 466:52]
  wire [7:0] _GEN_2919 = opcode_2 == 4'hf ? _GEN_1893 : _GEN_2661; // @[executor.scala 466:52]
  wire [7:0] _GEN_2920 = opcode_2 == 4'hf ? _GEN_1894 : _GEN_2662; // @[executor.scala 466:52]
  wire [7:0] _GEN_2921 = opcode_2 == 4'hf ? _GEN_1895 : _GEN_2663; // @[executor.scala 466:52]
  wire [7:0] _GEN_2922 = opcode_2 == 4'hf ? _GEN_1896 : _GEN_2664; // @[executor.scala 466:52]
  wire [7:0] _GEN_2923 = opcode_2 == 4'hf ? _GEN_1897 : _GEN_2665; // @[executor.scala 466:52]
  wire [7:0] _GEN_2924 = opcode_2 == 4'hf ? _GEN_1898 : _GEN_2666; // @[executor.scala 466:52]
  wire [7:0] _GEN_2925 = opcode_2 == 4'hf ? _GEN_1899 : _GEN_2667; // @[executor.scala 466:52]
  wire [7:0] _GEN_2926 = opcode_2 == 4'hf ? _GEN_1900 : _GEN_2668; // @[executor.scala 466:52]
  wire [7:0] _GEN_2927 = opcode_2 == 4'hf ? _GEN_1901 : _GEN_2669; // @[executor.scala 466:52]
  wire [7:0] _GEN_2928 = opcode_2 == 4'hf ? _GEN_1902 : _GEN_2670; // @[executor.scala 466:52]
  wire [7:0] _GEN_2929 = opcode_2 == 4'hf ? _GEN_1903 : _GEN_2671; // @[executor.scala 466:52]
  wire [7:0] _GEN_2930 = opcode_2 == 4'hf ? _GEN_1904 : _GEN_2672; // @[executor.scala 466:52]
  wire [7:0] _GEN_2931 = opcode_2 == 4'hf ? _GEN_1905 : _GEN_2673; // @[executor.scala 466:52]
  wire [7:0] _GEN_2932 = opcode_2 == 4'hf ? _GEN_1906 : _GEN_2674; // @[executor.scala 466:52]
  wire [7:0] _GEN_2933 = opcode_2 == 4'hf ? _GEN_1907 : _GEN_2675; // @[executor.scala 466:52]
  wire [7:0] _GEN_2934 = opcode_2 == 4'hf ? _GEN_1908 : _GEN_2676; // @[executor.scala 466:52]
  wire [7:0] _GEN_2935 = opcode_2 == 4'hf ? _GEN_1909 : _GEN_2677; // @[executor.scala 466:52]
  wire [7:0] _GEN_2936 = opcode_2 == 4'hf ? _GEN_1910 : _GEN_2678; // @[executor.scala 466:52]
  wire [7:0] _GEN_2937 = opcode_2 == 4'hf ? _GEN_1911 : _GEN_2679; // @[executor.scala 466:52]
  wire [7:0] _GEN_2938 = opcode_2 == 4'hf ? _GEN_1912 : _GEN_2680; // @[executor.scala 466:52]
  wire [7:0] _GEN_2939 = opcode_2 == 4'hf ? _GEN_1913 : _GEN_2681; // @[executor.scala 466:52]
  wire [7:0] _GEN_2940 = opcode_2 == 4'hf ? _GEN_1914 : _GEN_2682; // @[executor.scala 466:52]
  wire [7:0] _GEN_2941 = opcode_2 == 4'hf ? _GEN_1915 : _GEN_2683; // @[executor.scala 466:52]
  wire [7:0] _GEN_2942 = opcode_2 == 4'hf ? _GEN_1916 : _GEN_2684; // @[executor.scala 466:52]
  wire [7:0] _GEN_2943 = opcode_2 == 4'hf ? _GEN_1917 : _GEN_2685; // @[executor.scala 466:52]
  wire [7:0] _GEN_2944 = opcode_2 == 4'hf ? _GEN_1918 : _GEN_2686; // @[executor.scala 466:52]
  wire [7:0] _GEN_2945 = opcode_2 == 4'hf ? _GEN_1919 : _GEN_2687; // @[executor.scala 466:52]
  wire [7:0] _GEN_2946 = opcode_2 == 4'hf ? _GEN_1920 : _GEN_2688; // @[executor.scala 466:52]
  wire [7:0] _GEN_2947 = opcode_2 == 4'hf ? _GEN_1921 : _GEN_2689; // @[executor.scala 466:52]
  wire [7:0] _GEN_2948 = opcode_2 == 4'hf ? _GEN_1922 : _GEN_2690; // @[executor.scala 466:52]
  wire [7:0] _GEN_2949 = opcode_2 == 4'hf ? _GEN_1923 : _GEN_2691; // @[executor.scala 466:52]
  wire [7:0] _GEN_2950 = opcode_2 == 4'hf ? _GEN_1924 : _GEN_2692; // @[executor.scala 466:52]
  wire [7:0] _GEN_2951 = opcode_2 == 4'hf ? _GEN_1925 : _GEN_2693; // @[executor.scala 466:52]
  wire [7:0] _GEN_2952 = opcode_2 == 4'hf ? _GEN_1926 : _GEN_2694; // @[executor.scala 466:52]
  wire [7:0] _GEN_2953 = opcode_2 == 4'hf ? _GEN_1927 : _GEN_2695; // @[executor.scala 466:52]
  wire [7:0] _GEN_2954 = opcode_2 == 4'hf ? _GEN_1928 : _GEN_2696; // @[executor.scala 466:52]
  wire [7:0] _GEN_2955 = opcode_2 == 4'hf ? _GEN_1929 : _GEN_2697; // @[executor.scala 466:52]
  wire [7:0] _GEN_2956 = opcode_2 == 4'hf ? _GEN_1930 : _GEN_2698; // @[executor.scala 466:52]
  wire [7:0] _GEN_2957 = opcode_2 == 4'hf ? _GEN_1931 : _GEN_2699; // @[executor.scala 466:52]
  wire [7:0] _GEN_2958 = opcode_2 == 4'hf ? _GEN_1932 : _GEN_2700; // @[executor.scala 466:52]
  wire [7:0] _GEN_2959 = opcode_2 == 4'hf ? _GEN_1933 : _GEN_2701; // @[executor.scala 466:52]
  wire [7:0] _GEN_2960 = opcode_2 == 4'hf ? _GEN_1934 : _GEN_2702; // @[executor.scala 466:52]
  wire [7:0] _GEN_2961 = opcode_2 == 4'hf ? _GEN_1935 : _GEN_2703; // @[executor.scala 466:52]
  wire [7:0] _GEN_2962 = opcode_2 == 4'hf ? _GEN_1936 : _GEN_2704; // @[executor.scala 466:52]
  wire [7:0] _GEN_2963 = opcode_2 == 4'hf ? _GEN_1937 : _GEN_2705; // @[executor.scala 466:52]
  wire [7:0] _GEN_2964 = opcode_2 == 4'hf ? _GEN_1938 : _GEN_2706; // @[executor.scala 466:52]
  wire [7:0] _GEN_2965 = opcode_2 == 4'hf ? _GEN_1939 : _GEN_2707; // @[executor.scala 466:52]
  wire [7:0] _GEN_2966 = opcode_2 == 4'hf ? _GEN_1940 : _GEN_2708; // @[executor.scala 466:52]
  wire [7:0] _GEN_2967 = opcode_2 == 4'hf ? _GEN_1941 : _GEN_2709; // @[executor.scala 466:52]
  wire [7:0] _GEN_2968 = opcode_2 == 4'hf ? _GEN_1942 : _GEN_2710; // @[executor.scala 466:52]
  wire [7:0] _GEN_2969 = opcode_2 == 4'hf ? _GEN_1943 : _GEN_2711; // @[executor.scala 466:52]
  wire [7:0] _GEN_2970 = opcode_2 == 4'hf ? _GEN_1944 : _GEN_2712; // @[executor.scala 466:52]
  wire [7:0] _GEN_2971 = opcode_2 == 4'hf ? _GEN_1945 : _GEN_2713; // @[executor.scala 466:52]
  wire [7:0] _GEN_2972 = opcode_2 == 4'hf ? _GEN_1946 : _GEN_2714; // @[executor.scala 466:52]
  wire [7:0] _GEN_2973 = opcode_2 == 4'hf ? _GEN_1947 : _GEN_2715; // @[executor.scala 466:52]
  wire [7:0] _GEN_2974 = opcode_2 == 4'hf ? _GEN_1948 : _GEN_2716; // @[executor.scala 466:52]
  wire [7:0] _GEN_2975 = opcode_2 == 4'hf ? _GEN_1949 : _GEN_2717; // @[executor.scala 466:52]
  wire [7:0] _GEN_2976 = opcode_2 == 4'hf ? _GEN_1950 : _GEN_2718; // @[executor.scala 466:52]
  wire [7:0] _GEN_2977 = opcode_2 == 4'hf ? _GEN_1951 : _GEN_2719; // @[executor.scala 466:52]
  wire [7:0] _GEN_2978 = opcode_2 == 4'hf ? _GEN_1952 : _GEN_2720; // @[executor.scala 466:52]
  wire [7:0] _GEN_2979 = opcode_2 == 4'hf ? _GEN_1953 : _GEN_2721; // @[executor.scala 466:52]
  wire [7:0] _GEN_2980 = opcode_2 == 4'hf ? _GEN_1954 : _GEN_2722; // @[executor.scala 466:52]
  wire [7:0] _GEN_2981 = opcode_2 == 4'hf ? _GEN_1955 : _GEN_2723; // @[executor.scala 466:52]
  wire [7:0] _GEN_2982 = opcode_2 == 4'hf ? _GEN_1956 : _GEN_2724; // @[executor.scala 466:52]
  wire [7:0] _GEN_2983 = opcode_2 == 4'hf ? _GEN_1957 : _GEN_2725; // @[executor.scala 466:52]
  wire [7:0] _GEN_2984 = opcode_2 == 4'hf ? _GEN_1958 : _GEN_2726; // @[executor.scala 466:52]
  wire [7:0] _GEN_2985 = opcode_2 == 4'hf ? _GEN_1959 : _GEN_2727; // @[executor.scala 466:52]
  wire [7:0] _GEN_2986 = opcode_2 == 4'hf ? _GEN_1960 : _GEN_2728; // @[executor.scala 466:52]
  wire [7:0] _GEN_2987 = opcode_2 == 4'hf ? _GEN_1961 : _GEN_2729; // @[executor.scala 466:52]
  wire [7:0] _GEN_2988 = opcode_2 == 4'hf ? _GEN_1962 : _GEN_2730; // @[executor.scala 466:52]
  wire [7:0] _GEN_2989 = opcode_2 == 4'hf ? _GEN_1963 : _GEN_2731; // @[executor.scala 466:52]
  wire [7:0] _GEN_2990 = opcode_2 == 4'hf ? _GEN_1964 : _GEN_2732; // @[executor.scala 466:52]
  wire [7:0] _GEN_2991 = opcode_2 == 4'hf ? _GEN_1965 : _GEN_2733; // @[executor.scala 466:52]
  wire [7:0] _GEN_2992 = opcode_2 == 4'hf ? _GEN_1966 : _GEN_2734; // @[executor.scala 466:52]
  wire [7:0] _GEN_2993 = opcode_2 == 4'hf ? _GEN_1967 : _GEN_2735; // @[executor.scala 466:52]
  wire [7:0] _GEN_2994 = opcode_2 == 4'hf ? _GEN_1968 : _GEN_2736; // @[executor.scala 466:52]
  wire [7:0] _GEN_2995 = opcode_2 == 4'hf ? _GEN_1969 : _GEN_2737; // @[executor.scala 466:52]
  wire [7:0] _GEN_2996 = opcode_2 == 4'hf ? _GEN_1970 : _GEN_2738; // @[executor.scala 466:52]
  wire [7:0] _GEN_2997 = opcode_2 == 4'hf ? _GEN_1971 : _GEN_2739; // @[executor.scala 466:52]
  wire [7:0] _GEN_2998 = opcode_2 == 4'hf ? _GEN_1972 : _GEN_2740; // @[executor.scala 466:52]
  wire [7:0] _GEN_2999 = opcode_2 == 4'hf ? _GEN_1973 : _GEN_2741; // @[executor.scala 466:52]
  wire [7:0] _GEN_3000 = opcode_2 == 4'hf ? _GEN_1974 : _GEN_2742; // @[executor.scala 466:52]
  wire [7:0] _GEN_3001 = opcode_2 == 4'hf ? _GEN_1975 : _GEN_2743; // @[executor.scala 466:52]
  wire [7:0] _GEN_3002 = opcode_2 == 4'hf ? _GEN_1976 : _GEN_2744; // @[executor.scala 466:52]
  wire [7:0] _GEN_3003 = opcode_2 == 4'hf ? _GEN_1977 : _GEN_2745; // @[executor.scala 466:52]
  wire [7:0] _GEN_3004 = opcode_2 == 4'hf ? _GEN_1978 : _GEN_2746; // @[executor.scala 466:52]
  wire [7:0] _GEN_3005 = opcode_2 == 4'hf ? _GEN_1979 : _GEN_2747; // @[executor.scala 466:52]
  wire [7:0] _GEN_3006 = opcode_2 == 4'hf ? _GEN_1980 : _GEN_2748; // @[executor.scala 466:52]
  wire [7:0] _GEN_3007 = opcode_2 == 4'hf ? _GEN_1981 : _GEN_2749; // @[executor.scala 466:52]
  wire [7:0] _GEN_3008 = opcode_2 == 4'hf ? _GEN_1982 : _GEN_2750; // @[executor.scala 466:52]
  wire [7:0] _GEN_3009 = opcode_2 == 4'hf ? _GEN_1983 : _GEN_2751; // @[executor.scala 466:52]
  wire [7:0] _GEN_3010 = opcode_2 == 4'hf ? _GEN_1984 : _GEN_2752; // @[executor.scala 466:52]
  wire [7:0] _GEN_3011 = opcode_2 == 4'hf ? _GEN_1985 : _GEN_2753; // @[executor.scala 466:52]
  wire [7:0] _GEN_3012 = opcode_2 == 4'hf ? _GEN_1986 : _GEN_2754; // @[executor.scala 466:52]
  wire [7:0] _GEN_3013 = opcode_2 == 4'hf ? _GEN_1987 : _GEN_2755; // @[executor.scala 466:52]
  wire [7:0] _GEN_3014 = opcode_2 == 4'hf ? _GEN_1988 : _GEN_2756; // @[executor.scala 466:52]
  wire [7:0] _GEN_3015 = opcode_2 == 4'hf ? _GEN_1989 : _GEN_2757; // @[executor.scala 466:52]
  wire [7:0] _GEN_3016 = opcode_2 == 4'hf ? _GEN_1990 : _GEN_2758; // @[executor.scala 466:52]
  wire [7:0] _GEN_3017 = opcode_2 == 4'hf ? _GEN_1991 : _GEN_2759; // @[executor.scala 466:52]
  wire [7:0] _GEN_3018 = opcode_2 == 4'hf ? _GEN_1992 : _GEN_2760; // @[executor.scala 466:52]
  wire [7:0] _GEN_3019 = opcode_2 == 4'hf ? _GEN_1993 : _GEN_2761; // @[executor.scala 466:52]
  wire [7:0] _GEN_3020 = opcode_2 == 4'hf ? _GEN_1994 : _GEN_2762; // @[executor.scala 466:52]
  wire [7:0] _GEN_3021 = opcode_2 == 4'hf ? _GEN_1995 : _GEN_2763; // @[executor.scala 466:52]
  wire [7:0] _GEN_3022 = opcode_2 == 4'hf ? _GEN_1996 : _GEN_2764; // @[executor.scala 466:52]
  wire [7:0] _GEN_3023 = opcode_2 == 4'hf ? _GEN_1997 : _GEN_2765; // @[executor.scala 466:52]
  wire [7:0] _GEN_3024 = opcode_2 == 4'hf ? _GEN_1998 : _GEN_2766; // @[executor.scala 466:52]
  wire [7:0] _GEN_3025 = opcode_2 == 4'hf ? _GEN_1999 : _GEN_2767; // @[executor.scala 466:52]
  wire [7:0] _GEN_3026 = opcode_2 == 4'hf ? _GEN_2000 : _GEN_2768; // @[executor.scala 466:52]
  wire [7:0] _GEN_3027 = opcode_2 == 4'hf ? _GEN_2001 : _GEN_2769; // @[executor.scala 466:52]
  wire [7:0] _GEN_3028 = opcode_2 == 4'hf ? _GEN_2002 : _GEN_2770; // @[executor.scala 466:52]
  wire [7:0] _GEN_3029 = opcode_2 == 4'hf ? _GEN_2003 : _GEN_2771; // @[executor.scala 466:52]
  wire [7:0] _GEN_3030 = opcode_2 == 4'hf ? _GEN_2004 : _GEN_2772; // @[executor.scala 466:52]
  wire [7:0] _GEN_3031 = opcode_2 == 4'hf ? _GEN_2005 : _GEN_2773; // @[executor.scala 466:52]
  wire [7:0] _GEN_3032 = opcode_2 == 4'hf ? _GEN_2006 : _GEN_2774; // @[executor.scala 466:52]
  wire [7:0] _GEN_3033 = opcode_2 == 4'hf ? _GEN_2007 : _GEN_2775; // @[executor.scala 466:52]
  wire [7:0] _GEN_3034 = opcode_2 == 4'hf ? _GEN_2008 : _GEN_2776; // @[executor.scala 466:52]
  wire [7:0] _GEN_3035 = opcode_2 == 4'hf ? _GEN_2009 : _GEN_2777; // @[executor.scala 466:52]
  wire [7:0] _GEN_3036 = opcode_2 == 4'hf ? _GEN_2010 : _GEN_2778; // @[executor.scala 466:52]
  wire [7:0] _GEN_3037 = opcode_2 == 4'hf ? _GEN_2011 : _GEN_2779; // @[executor.scala 466:52]
  wire [7:0] _GEN_3038 = opcode_2 == 4'hf ? _GEN_2012 : _GEN_2780; // @[executor.scala 466:52]
  wire [7:0] _GEN_3039 = opcode_2 == 4'hf ? _GEN_2013 : _GEN_2781; // @[executor.scala 466:52]
  wire [7:0] _GEN_3040 = opcode_2 == 4'hf ? _GEN_2014 : _GEN_2782; // @[executor.scala 466:52]
  wire [7:0] _GEN_3041 = opcode_2 == 4'hf ? _GEN_2015 : _GEN_2783; // @[executor.scala 466:52]
  wire [7:0] _GEN_3042 = opcode_2 == 4'hf ? _GEN_2016 : _GEN_2784; // @[executor.scala 466:52]
  wire [7:0] _GEN_3043 = opcode_2 == 4'hf ? _GEN_2017 : _GEN_2785; // @[executor.scala 466:52]
  wire [7:0] _GEN_3044 = opcode_2 == 4'hf ? _GEN_2018 : _GEN_2786; // @[executor.scala 466:52]
  wire [7:0] _GEN_3045 = opcode_2 == 4'hf ? _GEN_2019 : _GEN_2787; // @[executor.scala 466:52]
  wire [7:0] _GEN_3046 = opcode_2 == 4'hf ? _GEN_2020 : _GEN_2788; // @[executor.scala 466:52]
  wire [7:0] _GEN_3047 = opcode_2 == 4'hf ? _GEN_2021 : _GEN_2789; // @[executor.scala 466:52]
  wire [7:0] _GEN_3048 = opcode_2 == 4'hf ? _GEN_2022 : _GEN_2790; // @[executor.scala 466:52]
  wire [7:0] _GEN_3049 = opcode_2 == 4'hf ? _GEN_2023 : _GEN_2791; // @[executor.scala 466:52]
  wire [7:0] _GEN_3050 = opcode_2 == 4'hf ? _GEN_2024 : _GEN_2792; // @[executor.scala 466:52]
  wire [7:0] _GEN_3051 = opcode_2 == 4'hf ? _GEN_2025 : _GEN_2793; // @[executor.scala 466:52]
  wire [7:0] _GEN_3052 = opcode_2 == 4'hf ? _GEN_2026 : _GEN_2794; // @[executor.scala 466:52]
  wire [7:0] _GEN_3053 = opcode_2 == 4'hf ? _GEN_2027 : _GEN_2795; // @[executor.scala 466:52]
  wire [7:0] _GEN_3054 = opcode_2 == 4'hf ? _GEN_2028 : _GEN_2796; // @[executor.scala 466:52]
  wire [7:0] _GEN_3055 = opcode_2 == 4'hf ? _GEN_2029 : _GEN_2797; // @[executor.scala 466:52]
  wire [7:0] _GEN_3056 = opcode_2 == 4'hf ? _GEN_2030 : _GEN_2798; // @[executor.scala 466:52]
  wire [7:0] _GEN_3057 = opcode_2 == 4'hf ? _GEN_2031 : _GEN_2799; // @[executor.scala 466:52]
  wire [7:0] _GEN_3058 = opcode_2 == 4'hf ? _GEN_2032 : _GEN_2800; // @[executor.scala 466:52]
  wire [7:0] _GEN_3059 = opcode_2 == 4'hf ? _GEN_2033 : _GEN_2801; // @[executor.scala 466:52]
  wire [7:0] _GEN_3060 = opcode_2 == 4'hf ? _GEN_2034 : _GEN_2802; // @[executor.scala 466:52]
  wire [7:0] _GEN_3061 = opcode_2 == 4'hf ? _GEN_2035 : _GEN_2803; // @[executor.scala 466:52]
  wire [7:0] _GEN_3062 = opcode_2 == 4'hf ? _GEN_2036 : _GEN_2804; // @[executor.scala 466:52]
  wire [7:0] _GEN_3063 = opcode_2 == 4'hf ? _GEN_2037 : _GEN_2805; // @[executor.scala 466:52]
  wire [7:0] _GEN_3064 = opcode_2 == 4'hf ? _GEN_2038 : _GEN_2806; // @[executor.scala 466:52]
  wire [7:0] _GEN_3065 = opcode_2 == 4'hf ? _GEN_2039 : _GEN_2807; // @[executor.scala 466:52]
  wire [7:0] _GEN_3066 = opcode_2 == 4'hf ? _GEN_2040 : _GEN_2808; // @[executor.scala 466:52]
  wire [7:0] _GEN_3067 = opcode_2 == 4'hf ? _GEN_2041 : _GEN_2809; // @[executor.scala 466:52]
  wire [7:0] _GEN_3068 = opcode_2 == 4'hf ? _GEN_2042 : _GEN_2810; // @[executor.scala 466:52]
  wire [7:0] _GEN_3069 = opcode_2 == 4'hf ? _GEN_2043 : _GEN_2811; // @[executor.scala 466:52]
  wire [7:0] _GEN_3070 = opcode_2 == 4'hf ? _GEN_2044 : _GEN_2812; // @[executor.scala 466:52]
  wire [7:0] _GEN_3071 = opcode_2 == 4'hf ? _GEN_2045 : _GEN_2813; // @[executor.scala 466:52]
  wire [7:0] _GEN_3072 = opcode_2 == 4'hf ? _GEN_2046 : _GEN_2814; // @[executor.scala 466:52]
  wire [7:0] _GEN_3073 = opcode_2 == 4'hf ? _GEN_2047 : _GEN_2815; // @[executor.scala 466:52]
  wire [7:0] _GEN_3074 = opcode_2 == 4'hf ? _GEN_2048 : _GEN_2816; // @[executor.scala 466:52]
  wire [7:0] _GEN_3075 = opcode_2 == 4'hf ? _GEN_2049 : _GEN_2817; // @[executor.scala 466:52]
  wire [7:0] _GEN_3076 = opcode_2 == 4'hf ? _GEN_2050 : _GEN_2818; // @[executor.scala 466:52]
  wire [7:0] _GEN_3077 = opcode_2 == 4'hf ? _GEN_2051 : _GEN_2819; // @[executor.scala 466:52]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_3 = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8658 = {{2'd0}, dst_offset_3}; // @[executor.scala 473:49]
  wire [7:0] byte_768 = field_3[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3078 = mask_3[0] ? byte_768 : _GEN_2822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_769 = field_3[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3079 = mask_3[1] ? byte_769 : _GEN_2823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_770 = field_3[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3080 = mask_3[2] ? byte_770 : _GEN_2824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_771 = field_3[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3081 = mask_3[3] ? byte_771 : _GEN_2825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3082 = _GEN_8658 == 8'h0 ? _GEN_3078 : _GEN_2822; // @[executor.scala 473:84]
  wire [7:0] _GEN_3083 = _GEN_8658 == 8'h0 ? _GEN_3079 : _GEN_2823; // @[executor.scala 473:84]
  wire [7:0] _GEN_3084 = _GEN_8658 == 8'h0 ? _GEN_3080 : _GEN_2824; // @[executor.scala 473:84]
  wire [7:0] _GEN_3085 = _GEN_8658 == 8'h0 ? _GEN_3081 : _GEN_2825; // @[executor.scala 473:84]
  wire [7:0] _GEN_3086 = mask_3[0] ? byte_768 : _GEN_2826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3087 = mask_3[1] ? byte_769 : _GEN_2827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3088 = mask_3[2] ? byte_770 : _GEN_2828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3089 = mask_3[3] ? byte_771 : _GEN_2829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3090 = _GEN_8658 == 8'h1 ? _GEN_3086 : _GEN_2826; // @[executor.scala 473:84]
  wire [7:0] _GEN_3091 = _GEN_8658 == 8'h1 ? _GEN_3087 : _GEN_2827; // @[executor.scala 473:84]
  wire [7:0] _GEN_3092 = _GEN_8658 == 8'h1 ? _GEN_3088 : _GEN_2828; // @[executor.scala 473:84]
  wire [7:0] _GEN_3093 = _GEN_8658 == 8'h1 ? _GEN_3089 : _GEN_2829; // @[executor.scala 473:84]
  wire [7:0] _GEN_3094 = mask_3[0] ? byte_768 : _GEN_2830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3095 = mask_3[1] ? byte_769 : _GEN_2831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3096 = mask_3[2] ? byte_770 : _GEN_2832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3097 = mask_3[3] ? byte_771 : _GEN_2833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3098 = _GEN_8658 == 8'h2 ? _GEN_3094 : _GEN_2830; // @[executor.scala 473:84]
  wire [7:0] _GEN_3099 = _GEN_8658 == 8'h2 ? _GEN_3095 : _GEN_2831; // @[executor.scala 473:84]
  wire [7:0] _GEN_3100 = _GEN_8658 == 8'h2 ? _GEN_3096 : _GEN_2832; // @[executor.scala 473:84]
  wire [7:0] _GEN_3101 = _GEN_8658 == 8'h2 ? _GEN_3097 : _GEN_2833; // @[executor.scala 473:84]
  wire [7:0] _GEN_3102 = mask_3[0] ? byte_768 : _GEN_2834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3103 = mask_3[1] ? byte_769 : _GEN_2835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3104 = mask_3[2] ? byte_770 : _GEN_2836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3105 = mask_3[3] ? byte_771 : _GEN_2837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3106 = _GEN_8658 == 8'h3 ? _GEN_3102 : _GEN_2834; // @[executor.scala 473:84]
  wire [7:0] _GEN_3107 = _GEN_8658 == 8'h3 ? _GEN_3103 : _GEN_2835; // @[executor.scala 473:84]
  wire [7:0] _GEN_3108 = _GEN_8658 == 8'h3 ? _GEN_3104 : _GEN_2836; // @[executor.scala 473:84]
  wire [7:0] _GEN_3109 = _GEN_8658 == 8'h3 ? _GEN_3105 : _GEN_2837; // @[executor.scala 473:84]
  wire [7:0] _GEN_3110 = mask_3[0] ? byte_768 : _GEN_2838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3111 = mask_3[1] ? byte_769 : _GEN_2839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3112 = mask_3[2] ? byte_770 : _GEN_2840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3113 = mask_3[3] ? byte_771 : _GEN_2841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3114 = _GEN_8658 == 8'h4 ? _GEN_3110 : _GEN_2838; // @[executor.scala 473:84]
  wire [7:0] _GEN_3115 = _GEN_8658 == 8'h4 ? _GEN_3111 : _GEN_2839; // @[executor.scala 473:84]
  wire [7:0] _GEN_3116 = _GEN_8658 == 8'h4 ? _GEN_3112 : _GEN_2840; // @[executor.scala 473:84]
  wire [7:0] _GEN_3117 = _GEN_8658 == 8'h4 ? _GEN_3113 : _GEN_2841; // @[executor.scala 473:84]
  wire [7:0] _GEN_3118 = mask_3[0] ? byte_768 : _GEN_2842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3119 = mask_3[1] ? byte_769 : _GEN_2843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3120 = mask_3[2] ? byte_770 : _GEN_2844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3121 = mask_3[3] ? byte_771 : _GEN_2845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3122 = _GEN_8658 == 8'h5 ? _GEN_3118 : _GEN_2842; // @[executor.scala 473:84]
  wire [7:0] _GEN_3123 = _GEN_8658 == 8'h5 ? _GEN_3119 : _GEN_2843; // @[executor.scala 473:84]
  wire [7:0] _GEN_3124 = _GEN_8658 == 8'h5 ? _GEN_3120 : _GEN_2844; // @[executor.scala 473:84]
  wire [7:0] _GEN_3125 = _GEN_8658 == 8'h5 ? _GEN_3121 : _GEN_2845; // @[executor.scala 473:84]
  wire [7:0] _GEN_3126 = mask_3[0] ? byte_768 : _GEN_2846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3127 = mask_3[1] ? byte_769 : _GEN_2847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3128 = mask_3[2] ? byte_770 : _GEN_2848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3129 = mask_3[3] ? byte_771 : _GEN_2849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3130 = _GEN_8658 == 8'h6 ? _GEN_3126 : _GEN_2846; // @[executor.scala 473:84]
  wire [7:0] _GEN_3131 = _GEN_8658 == 8'h6 ? _GEN_3127 : _GEN_2847; // @[executor.scala 473:84]
  wire [7:0] _GEN_3132 = _GEN_8658 == 8'h6 ? _GEN_3128 : _GEN_2848; // @[executor.scala 473:84]
  wire [7:0] _GEN_3133 = _GEN_8658 == 8'h6 ? _GEN_3129 : _GEN_2849; // @[executor.scala 473:84]
  wire [7:0] _GEN_3134 = mask_3[0] ? byte_768 : _GEN_2850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3135 = mask_3[1] ? byte_769 : _GEN_2851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3136 = mask_3[2] ? byte_770 : _GEN_2852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3137 = mask_3[3] ? byte_771 : _GEN_2853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3138 = _GEN_8658 == 8'h7 ? _GEN_3134 : _GEN_2850; // @[executor.scala 473:84]
  wire [7:0] _GEN_3139 = _GEN_8658 == 8'h7 ? _GEN_3135 : _GEN_2851; // @[executor.scala 473:84]
  wire [7:0] _GEN_3140 = _GEN_8658 == 8'h7 ? _GEN_3136 : _GEN_2852; // @[executor.scala 473:84]
  wire [7:0] _GEN_3141 = _GEN_8658 == 8'h7 ? _GEN_3137 : _GEN_2853; // @[executor.scala 473:84]
  wire [7:0] _GEN_3142 = mask_3[0] ? byte_768 : _GEN_2854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3143 = mask_3[1] ? byte_769 : _GEN_2855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3144 = mask_3[2] ? byte_770 : _GEN_2856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3145 = mask_3[3] ? byte_771 : _GEN_2857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3146 = _GEN_8658 == 8'h8 ? _GEN_3142 : _GEN_2854; // @[executor.scala 473:84]
  wire [7:0] _GEN_3147 = _GEN_8658 == 8'h8 ? _GEN_3143 : _GEN_2855; // @[executor.scala 473:84]
  wire [7:0] _GEN_3148 = _GEN_8658 == 8'h8 ? _GEN_3144 : _GEN_2856; // @[executor.scala 473:84]
  wire [7:0] _GEN_3149 = _GEN_8658 == 8'h8 ? _GEN_3145 : _GEN_2857; // @[executor.scala 473:84]
  wire [7:0] _GEN_3150 = mask_3[0] ? byte_768 : _GEN_2858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3151 = mask_3[1] ? byte_769 : _GEN_2859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3152 = mask_3[2] ? byte_770 : _GEN_2860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3153 = mask_3[3] ? byte_771 : _GEN_2861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3154 = _GEN_8658 == 8'h9 ? _GEN_3150 : _GEN_2858; // @[executor.scala 473:84]
  wire [7:0] _GEN_3155 = _GEN_8658 == 8'h9 ? _GEN_3151 : _GEN_2859; // @[executor.scala 473:84]
  wire [7:0] _GEN_3156 = _GEN_8658 == 8'h9 ? _GEN_3152 : _GEN_2860; // @[executor.scala 473:84]
  wire [7:0] _GEN_3157 = _GEN_8658 == 8'h9 ? _GEN_3153 : _GEN_2861; // @[executor.scala 473:84]
  wire [7:0] _GEN_3158 = mask_3[0] ? byte_768 : _GEN_2862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3159 = mask_3[1] ? byte_769 : _GEN_2863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3160 = mask_3[2] ? byte_770 : _GEN_2864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3161 = mask_3[3] ? byte_771 : _GEN_2865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3162 = _GEN_8658 == 8'ha ? _GEN_3158 : _GEN_2862; // @[executor.scala 473:84]
  wire [7:0] _GEN_3163 = _GEN_8658 == 8'ha ? _GEN_3159 : _GEN_2863; // @[executor.scala 473:84]
  wire [7:0] _GEN_3164 = _GEN_8658 == 8'ha ? _GEN_3160 : _GEN_2864; // @[executor.scala 473:84]
  wire [7:0] _GEN_3165 = _GEN_8658 == 8'ha ? _GEN_3161 : _GEN_2865; // @[executor.scala 473:84]
  wire [7:0] _GEN_3166 = mask_3[0] ? byte_768 : _GEN_2866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3167 = mask_3[1] ? byte_769 : _GEN_2867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3168 = mask_3[2] ? byte_770 : _GEN_2868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3169 = mask_3[3] ? byte_771 : _GEN_2869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3170 = _GEN_8658 == 8'hb ? _GEN_3166 : _GEN_2866; // @[executor.scala 473:84]
  wire [7:0] _GEN_3171 = _GEN_8658 == 8'hb ? _GEN_3167 : _GEN_2867; // @[executor.scala 473:84]
  wire [7:0] _GEN_3172 = _GEN_8658 == 8'hb ? _GEN_3168 : _GEN_2868; // @[executor.scala 473:84]
  wire [7:0] _GEN_3173 = _GEN_8658 == 8'hb ? _GEN_3169 : _GEN_2869; // @[executor.scala 473:84]
  wire [7:0] _GEN_3174 = mask_3[0] ? byte_768 : _GEN_2870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3175 = mask_3[1] ? byte_769 : _GEN_2871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3176 = mask_3[2] ? byte_770 : _GEN_2872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3177 = mask_3[3] ? byte_771 : _GEN_2873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3178 = _GEN_8658 == 8'hc ? _GEN_3174 : _GEN_2870; // @[executor.scala 473:84]
  wire [7:0] _GEN_3179 = _GEN_8658 == 8'hc ? _GEN_3175 : _GEN_2871; // @[executor.scala 473:84]
  wire [7:0] _GEN_3180 = _GEN_8658 == 8'hc ? _GEN_3176 : _GEN_2872; // @[executor.scala 473:84]
  wire [7:0] _GEN_3181 = _GEN_8658 == 8'hc ? _GEN_3177 : _GEN_2873; // @[executor.scala 473:84]
  wire [7:0] _GEN_3182 = mask_3[0] ? byte_768 : _GEN_2874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3183 = mask_3[1] ? byte_769 : _GEN_2875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3184 = mask_3[2] ? byte_770 : _GEN_2876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3185 = mask_3[3] ? byte_771 : _GEN_2877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3186 = _GEN_8658 == 8'hd ? _GEN_3182 : _GEN_2874; // @[executor.scala 473:84]
  wire [7:0] _GEN_3187 = _GEN_8658 == 8'hd ? _GEN_3183 : _GEN_2875; // @[executor.scala 473:84]
  wire [7:0] _GEN_3188 = _GEN_8658 == 8'hd ? _GEN_3184 : _GEN_2876; // @[executor.scala 473:84]
  wire [7:0] _GEN_3189 = _GEN_8658 == 8'hd ? _GEN_3185 : _GEN_2877; // @[executor.scala 473:84]
  wire [7:0] _GEN_3190 = mask_3[0] ? byte_768 : _GEN_2878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3191 = mask_3[1] ? byte_769 : _GEN_2879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3192 = mask_3[2] ? byte_770 : _GEN_2880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3193 = mask_3[3] ? byte_771 : _GEN_2881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3194 = _GEN_8658 == 8'he ? _GEN_3190 : _GEN_2878; // @[executor.scala 473:84]
  wire [7:0] _GEN_3195 = _GEN_8658 == 8'he ? _GEN_3191 : _GEN_2879; // @[executor.scala 473:84]
  wire [7:0] _GEN_3196 = _GEN_8658 == 8'he ? _GEN_3192 : _GEN_2880; // @[executor.scala 473:84]
  wire [7:0] _GEN_3197 = _GEN_8658 == 8'he ? _GEN_3193 : _GEN_2881; // @[executor.scala 473:84]
  wire [7:0] _GEN_3198 = mask_3[0] ? byte_768 : _GEN_2882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3199 = mask_3[1] ? byte_769 : _GEN_2883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3200 = mask_3[2] ? byte_770 : _GEN_2884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3201 = mask_3[3] ? byte_771 : _GEN_2885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3202 = _GEN_8658 == 8'hf ? _GEN_3198 : _GEN_2882; // @[executor.scala 473:84]
  wire [7:0] _GEN_3203 = _GEN_8658 == 8'hf ? _GEN_3199 : _GEN_2883; // @[executor.scala 473:84]
  wire [7:0] _GEN_3204 = _GEN_8658 == 8'hf ? _GEN_3200 : _GEN_2884; // @[executor.scala 473:84]
  wire [7:0] _GEN_3205 = _GEN_8658 == 8'hf ? _GEN_3201 : _GEN_2885; // @[executor.scala 473:84]
  wire [7:0] _GEN_3206 = mask_3[0] ? byte_768 : _GEN_2886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3207 = mask_3[1] ? byte_769 : _GEN_2887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3208 = mask_3[2] ? byte_770 : _GEN_2888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3209 = mask_3[3] ? byte_771 : _GEN_2889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3210 = _GEN_8658 == 8'h10 ? _GEN_3206 : _GEN_2886; // @[executor.scala 473:84]
  wire [7:0] _GEN_3211 = _GEN_8658 == 8'h10 ? _GEN_3207 : _GEN_2887; // @[executor.scala 473:84]
  wire [7:0] _GEN_3212 = _GEN_8658 == 8'h10 ? _GEN_3208 : _GEN_2888; // @[executor.scala 473:84]
  wire [7:0] _GEN_3213 = _GEN_8658 == 8'h10 ? _GEN_3209 : _GEN_2889; // @[executor.scala 473:84]
  wire [7:0] _GEN_3214 = mask_3[0] ? byte_768 : _GEN_2890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3215 = mask_3[1] ? byte_769 : _GEN_2891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3216 = mask_3[2] ? byte_770 : _GEN_2892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3217 = mask_3[3] ? byte_771 : _GEN_2893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3218 = _GEN_8658 == 8'h11 ? _GEN_3214 : _GEN_2890; // @[executor.scala 473:84]
  wire [7:0] _GEN_3219 = _GEN_8658 == 8'h11 ? _GEN_3215 : _GEN_2891; // @[executor.scala 473:84]
  wire [7:0] _GEN_3220 = _GEN_8658 == 8'h11 ? _GEN_3216 : _GEN_2892; // @[executor.scala 473:84]
  wire [7:0] _GEN_3221 = _GEN_8658 == 8'h11 ? _GEN_3217 : _GEN_2893; // @[executor.scala 473:84]
  wire [7:0] _GEN_3222 = mask_3[0] ? byte_768 : _GEN_2894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3223 = mask_3[1] ? byte_769 : _GEN_2895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3224 = mask_3[2] ? byte_770 : _GEN_2896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3225 = mask_3[3] ? byte_771 : _GEN_2897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3226 = _GEN_8658 == 8'h12 ? _GEN_3222 : _GEN_2894; // @[executor.scala 473:84]
  wire [7:0] _GEN_3227 = _GEN_8658 == 8'h12 ? _GEN_3223 : _GEN_2895; // @[executor.scala 473:84]
  wire [7:0] _GEN_3228 = _GEN_8658 == 8'h12 ? _GEN_3224 : _GEN_2896; // @[executor.scala 473:84]
  wire [7:0] _GEN_3229 = _GEN_8658 == 8'h12 ? _GEN_3225 : _GEN_2897; // @[executor.scala 473:84]
  wire [7:0] _GEN_3230 = mask_3[0] ? byte_768 : _GEN_2898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3231 = mask_3[1] ? byte_769 : _GEN_2899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3232 = mask_3[2] ? byte_770 : _GEN_2900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3233 = mask_3[3] ? byte_771 : _GEN_2901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3234 = _GEN_8658 == 8'h13 ? _GEN_3230 : _GEN_2898; // @[executor.scala 473:84]
  wire [7:0] _GEN_3235 = _GEN_8658 == 8'h13 ? _GEN_3231 : _GEN_2899; // @[executor.scala 473:84]
  wire [7:0] _GEN_3236 = _GEN_8658 == 8'h13 ? _GEN_3232 : _GEN_2900; // @[executor.scala 473:84]
  wire [7:0] _GEN_3237 = _GEN_8658 == 8'h13 ? _GEN_3233 : _GEN_2901; // @[executor.scala 473:84]
  wire [7:0] _GEN_3238 = mask_3[0] ? byte_768 : _GEN_2902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3239 = mask_3[1] ? byte_769 : _GEN_2903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3240 = mask_3[2] ? byte_770 : _GEN_2904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3241 = mask_3[3] ? byte_771 : _GEN_2905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3242 = _GEN_8658 == 8'h14 ? _GEN_3238 : _GEN_2902; // @[executor.scala 473:84]
  wire [7:0] _GEN_3243 = _GEN_8658 == 8'h14 ? _GEN_3239 : _GEN_2903; // @[executor.scala 473:84]
  wire [7:0] _GEN_3244 = _GEN_8658 == 8'h14 ? _GEN_3240 : _GEN_2904; // @[executor.scala 473:84]
  wire [7:0] _GEN_3245 = _GEN_8658 == 8'h14 ? _GEN_3241 : _GEN_2905; // @[executor.scala 473:84]
  wire [7:0] _GEN_3246 = mask_3[0] ? byte_768 : _GEN_2906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3247 = mask_3[1] ? byte_769 : _GEN_2907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3248 = mask_3[2] ? byte_770 : _GEN_2908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3249 = mask_3[3] ? byte_771 : _GEN_2909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3250 = _GEN_8658 == 8'h15 ? _GEN_3246 : _GEN_2906; // @[executor.scala 473:84]
  wire [7:0] _GEN_3251 = _GEN_8658 == 8'h15 ? _GEN_3247 : _GEN_2907; // @[executor.scala 473:84]
  wire [7:0] _GEN_3252 = _GEN_8658 == 8'h15 ? _GEN_3248 : _GEN_2908; // @[executor.scala 473:84]
  wire [7:0] _GEN_3253 = _GEN_8658 == 8'h15 ? _GEN_3249 : _GEN_2909; // @[executor.scala 473:84]
  wire [7:0] _GEN_3254 = mask_3[0] ? byte_768 : _GEN_2910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3255 = mask_3[1] ? byte_769 : _GEN_2911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3256 = mask_3[2] ? byte_770 : _GEN_2912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3257 = mask_3[3] ? byte_771 : _GEN_2913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3258 = _GEN_8658 == 8'h16 ? _GEN_3254 : _GEN_2910; // @[executor.scala 473:84]
  wire [7:0] _GEN_3259 = _GEN_8658 == 8'h16 ? _GEN_3255 : _GEN_2911; // @[executor.scala 473:84]
  wire [7:0] _GEN_3260 = _GEN_8658 == 8'h16 ? _GEN_3256 : _GEN_2912; // @[executor.scala 473:84]
  wire [7:0] _GEN_3261 = _GEN_8658 == 8'h16 ? _GEN_3257 : _GEN_2913; // @[executor.scala 473:84]
  wire [7:0] _GEN_3262 = mask_3[0] ? byte_768 : _GEN_2914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3263 = mask_3[1] ? byte_769 : _GEN_2915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3264 = mask_3[2] ? byte_770 : _GEN_2916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3265 = mask_3[3] ? byte_771 : _GEN_2917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3266 = _GEN_8658 == 8'h17 ? _GEN_3262 : _GEN_2914; // @[executor.scala 473:84]
  wire [7:0] _GEN_3267 = _GEN_8658 == 8'h17 ? _GEN_3263 : _GEN_2915; // @[executor.scala 473:84]
  wire [7:0] _GEN_3268 = _GEN_8658 == 8'h17 ? _GEN_3264 : _GEN_2916; // @[executor.scala 473:84]
  wire [7:0] _GEN_3269 = _GEN_8658 == 8'h17 ? _GEN_3265 : _GEN_2917; // @[executor.scala 473:84]
  wire [7:0] _GEN_3270 = mask_3[0] ? byte_768 : _GEN_2918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3271 = mask_3[1] ? byte_769 : _GEN_2919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3272 = mask_3[2] ? byte_770 : _GEN_2920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3273 = mask_3[3] ? byte_771 : _GEN_2921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3274 = _GEN_8658 == 8'h18 ? _GEN_3270 : _GEN_2918; // @[executor.scala 473:84]
  wire [7:0] _GEN_3275 = _GEN_8658 == 8'h18 ? _GEN_3271 : _GEN_2919; // @[executor.scala 473:84]
  wire [7:0] _GEN_3276 = _GEN_8658 == 8'h18 ? _GEN_3272 : _GEN_2920; // @[executor.scala 473:84]
  wire [7:0] _GEN_3277 = _GEN_8658 == 8'h18 ? _GEN_3273 : _GEN_2921; // @[executor.scala 473:84]
  wire [7:0] _GEN_3278 = mask_3[0] ? byte_768 : _GEN_2922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3279 = mask_3[1] ? byte_769 : _GEN_2923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3280 = mask_3[2] ? byte_770 : _GEN_2924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3281 = mask_3[3] ? byte_771 : _GEN_2925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3282 = _GEN_8658 == 8'h19 ? _GEN_3278 : _GEN_2922; // @[executor.scala 473:84]
  wire [7:0] _GEN_3283 = _GEN_8658 == 8'h19 ? _GEN_3279 : _GEN_2923; // @[executor.scala 473:84]
  wire [7:0] _GEN_3284 = _GEN_8658 == 8'h19 ? _GEN_3280 : _GEN_2924; // @[executor.scala 473:84]
  wire [7:0] _GEN_3285 = _GEN_8658 == 8'h19 ? _GEN_3281 : _GEN_2925; // @[executor.scala 473:84]
  wire [7:0] _GEN_3286 = mask_3[0] ? byte_768 : _GEN_2926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3287 = mask_3[1] ? byte_769 : _GEN_2927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3288 = mask_3[2] ? byte_770 : _GEN_2928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3289 = mask_3[3] ? byte_771 : _GEN_2929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3290 = _GEN_8658 == 8'h1a ? _GEN_3286 : _GEN_2926; // @[executor.scala 473:84]
  wire [7:0] _GEN_3291 = _GEN_8658 == 8'h1a ? _GEN_3287 : _GEN_2927; // @[executor.scala 473:84]
  wire [7:0] _GEN_3292 = _GEN_8658 == 8'h1a ? _GEN_3288 : _GEN_2928; // @[executor.scala 473:84]
  wire [7:0] _GEN_3293 = _GEN_8658 == 8'h1a ? _GEN_3289 : _GEN_2929; // @[executor.scala 473:84]
  wire [7:0] _GEN_3294 = mask_3[0] ? byte_768 : _GEN_2930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3295 = mask_3[1] ? byte_769 : _GEN_2931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3296 = mask_3[2] ? byte_770 : _GEN_2932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3297 = mask_3[3] ? byte_771 : _GEN_2933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3298 = _GEN_8658 == 8'h1b ? _GEN_3294 : _GEN_2930; // @[executor.scala 473:84]
  wire [7:0] _GEN_3299 = _GEN_8658 == 8'h1b ? _GEN_3295 : _GEN_2931; // @[executor.scala 473:84]
  wire [7:0] _GEN_3300 = _GEN_8658 == 8'h1b ? _GEN_3296 : _GEN_2932; // @[executor.scala 473:84]
  wire [7:0] _GEN_3301 = _GEN_8658 == 8'h1b ? _GEN_3297 : _GEN_2933; // @[executor.scala 473:84]
  wire [7:0] _GEN_3302 = mask_3[0] ? byte_768 : _GEN_2934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3303 = mask_3[1] ? byte_769 : _GEN_2935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3304 = mask_3[2] ? byte_770 : _GEN_2936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3305 = mask_3[3] ? byte_771 : _GEN_2937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3306 = _GEN_8658 == 8'h1c ? _GEN_3302 : _GEN_2934; // @[executor.scala 473:84]
  wire [7:0] _GEN_3307 = _GEN_8658 == 8'h1c ? _GEN_3303 : _GEN_2935; // @[executor.scala 473:84]
  wire [7:0] _GEN_3308 = _GEN_8658 == 8'h1c ? _GEN_3304 : _GEN_2936; // @[executor.scala 473:84]
  wire [7:0] _GEN_3309 = _GEN_8658 == 8'h1c ? _GEN_3305 : _GEN_2937; // @[executor.scala 473:84]
  wire [7:0] _GEN_3310 = mask_3[0] ? byte_768 : _GEN_2938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3311 = mask_3[1] ? byte_769 : _GEN_2939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3312 = mask_3[2] ? byte_770 : _GEN_2940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3313 = mask_3[3] ? byte_771 : _GEN_2941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3314 = _GEN_8658 == 8'h1d ? _GEN_3310 : _GEN_2938; // @[executor.scala 473:84]
  wire [7:0] _GEN_3315 = _GEN_8658 == 8'h1d ? _GEN_3311 : _GEN_2939; // @[executor.scala 473:84]
  wire [7:0] _GEN_3316 = _GEN_8658 == 8'h1d ? _GEN_3312 : _GEN_2940; // @[executor.scala 473:84]
  wire [7:0] _GEN_3317 = _GEN_8658 == 8'h1d ? _GEN_3313 : _GEN_2941; // @[executor.scala 473:84]
  wire [7:0] _GEN_3318 = mask_3[0] ? byte_768 : _GEN_2942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3319 = mask_3[1] ? byte_769 : _GEN_2943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3320 = mask_3[2] ? byte_770 : _GEN_2944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3321 = mask_3[3] ? byte_771 : _GEN_2945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3322 = _GEN_8658 == 8'h1e ? _GEN_3318 : _GEN_2942; // @[executor.scala 473:84]
  wire [7:0] _GEN_3323 = _GEN_8658 == 8'h1e ? _GEN_3319 : _GEN_2943; // @[executor.scala 473:84]
  wire [7:0] _GEN_3324 = _GEN_8658 == 8'h1e ? _GEN_3320 : _GEN_2944; // @[executor.scala 473:84]
  wire [7:0] _GEN_3325 = _GEN_8658 == 8'h1e ? _GEN_3321 : _GEN_2945; // @[executor.scala 473:84]
  wire [7:0] _GEN_3326 = mask_3[0] ? byte_768 : _GEN_2946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3327 = mask_3[1] ? byte_769 : _GEN_2947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3328 = mask_3[2] ? byte_770 : _GEN_2948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3329 = mask_3[3] ? byte_771 : _GEN_2949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3330 = _GEN_8658 == 8'h1f ? _GEN_3326 : _GEN_2946; // @[executor.scala 473:84]
  wire [7:0] _GEN_3331 = _GEN_8658 == 8'h1f ? _GEN_3327 : _GEN_2947; // @[executor.scala 473:84]
  wire [7:0] _GEN_3332 = _GEN_8658 == 8'h1f ? _GEN_3328 : _GEN_2948; // @[executor.scala 473:84]
  wire [7:0] _GEN_3333 = _GEN_8658 == 8'h1f ? _GEN_3329 : _GEN_2949; // @[executor.scala 473:84]
  wire [7:0] _GEN_3334 = mask_3[0] ? byte_768 : _GEN_2950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3335 = mask_3[1] ? byte_769 : _GEN_2951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3336 = mask_3[2] ? byte_770 : _GEN_2952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3337 = mask_3[3] ? byte_771 : _GEN_2953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3338 = _GEN_8658 == 8'h20 ? _GEN_3334 : _GEN_2950; // @[executor.scala 473:84]
  wire [7:0] _GEN_3339 = _GEN_8658 == 8'h20 ? _GEN_3335 : _GEN_2951; // @[executor.scala 473:84]
  wire [7:0] _GEN_3340 = _GEN_8658 == 8'h20 ? _GEN_3336 : _GEN_2952; // @[executor.scala 473:84]
  wire [7:0] _GEN_3341 = _GEN_8658 == 8'h20 ? _GEN_3337 : _GEN_2953; // @[executor.scala 473:84]
  wire [7:0] _GEN_3342 = mask_3[0] ? byte_768 : _GEN_2954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3343 = mask_3[1] ? byte_769 : _GEN_2955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3344 = mask_3[2] ? byte_770 : _GEN_2956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3345 = mask_3[3] ? byte_771 : _GEN_2957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3346 = _GEN_8658 == 8'h21 ? _GEN_3342 : _GEN_2954; // @[executor.scala 473:84]
  wire [7:0] _GEN_3347 = _GEN_8658 == 8'h21 ? _GEN_3343 : _GEN_2955; // @[executor.scala 473:84]
  wire [7:0] _GEN_3348 = _GEN_8658 == 8'h21 ? _GEN_3344 : _GEN_2956; // @[executor.scala 473:84]
  wire [7:0] _GEN_3349 = _GEN_8658 == 8'h21 ? _GEN_3345 : _GEN_2957; // @[executor.scala 473:84]
  wire [7:0] _GEN_3350 = mask_3[0] ? byte_768 : _GEN_2958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3351 = mask_3[1] ? byte_769 : _GEN_2959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3352 = mask_3[2] ? byte_770 : _GEN_2960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3353 = mask_3[3] ? byte_771 : _GEN_2961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3354 = _GEN_8658 == 8'h22 ? _GEN_3350 : _GEN_2958; // @[executor.scala 473:84]
  wire [7:0] _GEN_3355 = _GEN_8658 == 8'h22 ? _GEN_3351 : _GEN_2959; // @[executor.scala 473:84]
  wire [7:0] _GEN_3356 = _GEN_8658 == 8'h22 ? _GEN_3352 : _GEN_2960; // @[executor.scala 473:84]
  wire [7:0] _GEN_3357 = _GEN_8658 == 8'h22 ? _GEN_3353 : _GEN_2961; // @[executor.scala 473:84]
  wire [7:0] _GEN_3358 = mask_3[0] ? byte_768 : _GEN_2962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3359 = mask_3[1] ? byte_769 : _GEN_2963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3360 = mask_3[2] ? byte_770 : _GEN_2964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3361 = mask_3[3] ? byte_771 : _GEN_2965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3362 = _GEN_8658 == 8'h23 ? _GEN_3358 : _GEN_2962; // @[executor.scala 473:84]
  wire [7:0] _GEN_3363 = _GEN_8658 == 8'h23 ? _GEN_3359 : _GEN_2963; // @[executor.scala 473:84]
  wire [7:0] _GEN_3364 = _GEN_8658 == 8'h23 ? _GEN_3360 : _GEN_2964; // @[executor.scala 473:84]
  wire [7:0] _GEN_3365 = _GEN_8658 == 8'h23 ? _GEN_3361 : _GEN_2965; // @[executor.scala 473:84]
  wire [7:0] _GEN_3366 = mask_3[0] ? byte_768 : _GEN_2966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3367 = mask_3[1] ? byte_769 : _GEN_2967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3368 = mask_3[2] ? byte_770 : _GEN_2968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3369 = mask_3[3] ? byte_771 : _GEN_2969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3370 = _GEN_8658 == 8'h24 ? _GEN_3366 : _GEN_2966; // @[executor.scala 473:84]
  wire [7:0] _GEN_3371 = _GEN_8658 == 8'h24 ? _GEN_3367 : _GEN_2967; // @[executor.scala 473:84]
  wire [7:0] _GEN_3372 = _GEN_8658 == 8'h24 ? _GEN_3368 : _GEN_2968; // @[executor.scala 473:84]
  wire [7:0] _GEN_3373 = _GEN_8658 == 8'h24 ? _GEN_3369 : _GEN_2969; // @[executor.scala 473:84]
  wire [7:0] _GEN_3374 = mask_3[0] ? byte_768 : _GEN_2970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3375 = mask_3[1] ? byte_769 : _GEN_2971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3376 = mask_3[2] ? byte_770 : _GEN_2972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3377 = mask_3[3] ? byte_771 : _GEN_2973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3378 = _GEN_8658 == 8'h25 ? _GEN_3374 : _GEN_2970; // @[executor.scala 473:84]
  wire [7:0] _GEN_3379 = _GEN_8658 == 8'h25 ? _GEN_3375 : _GEN_2971; // @[executor.scala 473:84]
  wire [7:0] _GEN_3380 = _GEN_8658 == 8'h25 ? _GEN_3376 : _GEN_2972; // @[executor.scala 473:84]
  wire [7:0] _GEN_3381 = _GEN_8658 == 8'h25 ? _GEN_3377 : _GEN_2973; // @[executor.scala 473:84]
  wire [7:0] _GEN_3382 = mask_3[0] ? byte_768 : _GEN_2974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3383 = mask_3[1] ? byte_769 : _GEN_2975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3384 = mask_3[2] ? byte_770 : _GEN_2976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3385 = mask_3[3] ? byte_771 : _GEN_2977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3386 = _GEN_8658 == 8'h26 ? _GEN_3382 : _GEN_2974; // @[executor.scala 473:84]
  wire [7:0] _GEN_3387 = _GEN_8658 == 8'h26 ? _GEN_3383 : _GEN_2975; // @[executor.scala 473:84]
  wire [7:0] _GEN_3388 = _GEN_8658 == 8'h26 ? _GEN_3384 : _GEN_2976; // @[executor.scala 473:84]
  wire [7:0] _GEN_3389 = _GEN_8658 == 8'h26 ? _GEN_3385 : _GEN_2977; // @[executor.scala 473:84]
  wire [7:0] _GEN_3390 = mask_3[0] ? byte_768 : _GEN_2978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3391 = mask_3[1] ? byte_769 : _GEN_2979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3392 = mask_3[2] ? byte_770 : _GEN_2980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3393 = mask_3[3] ? byte_771 : _GEN_2981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3394 = _GEN_8658 == 8'h27 ? _GEN_3390 : _GEN_2978; // @[executor.scala 473:84]
  wire [7:0] _GEN_3395 = _GEN_8658 == 8'h27 ? _GEN_3391 : _GEN_2979; // @[executor.scala 473:84]
  wire [7:0] _GEN_3396 = _GEN_8658 == 8'h27 ? _GEN_3392 : _GEN_2980; // @[executor.scala 473:84]
  wire [7:0] _GEN_3397 = _GEN_8658 == 8'h27 ? _GEN_3393 : _GEN_2981; // @[executor.scala 473:84]
  wire [7:0] _GEN_3398 = mask_3[0] ? byte_768 : _GEN_2982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3399 = mask_3[1] ? byte_769 : _GEN_2983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3400 = mask_3[2] ? byte_770 : _GEN_2984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3401 = mask_3[3] ? byte_771 : _GEN_2985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3402 = _GEN_8658 == 8'h28 ? _GEN_3398 : _GEN_2982; // @[executor.scala 473:84]
  wire [7:0] _GEN_3403 = _GEN_8658 == 8'h28 ? _GEN_3399 : _GEN_2983; // @[executor.scala 473:84]
  wire [7:0] _GEN_3404 = _GEN_8658 == 8'h28 ? _GEN_3400 : _GEN_2984; // @[executor.scala 473:84]
  wire [7:0] _GEN_3405 = _GEN_8658 == 8'h28 ? _GEN_3401 : _GEN_2985; // @[executor.scala 473:84]
  wire [7:0] _GEN_3406 = mask_3[0] ? byte_768 : _GEN_2986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3407 = mask_3[1] ? byte_769 : _GEN_2987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3408 = mask_3[2] ? byte_770 : _GEN_2988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3409 = mask_3[3] ? byte_771 : _GEN_2989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3410 = _GEN_8658 == 8'h29 ? _GEN_3406 : _GEN_2986; // @[executor.scala 473:84]
  wire [7:0] _GEN_3411 = _GEN_8658 == 8'h29 ? _GEN_3407 : _GEN_2987; // @[executor.scala 473:84]
  wire [7:0] _GEN_3412 = _GEN_8658 == 8'h29 ? _GEN_3408 : _GEN_2988; // @[executor.scala 473:84]
  wire [7:0] _GEN_3413 = _GEN_8658 == 8'h29 ? _GEN_3409 : _GEN_2989; // @[executor.scala 473:84]
  wire [7:0] _GEN_3414 = mask_3[0] ? byte_768 : _GEN_2990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3415 = mask_3[1] ? byte_769 : _GEN_2991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3416 = mask_3[2] ? byte_770 : _GEN_2992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3417 = mask_3[3] ? byte_771 : _GEN_2993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3418 = _GEN_8658 == 8'h2a ? _GEN_3414 : _GEN_2990; // @[executor.scala 473:84]
  wire [7:0] _GEN_3419 = _GEN_8658 == 8'h2a ? _GEN_3415 : _GEN_2991; // @[executor.scala 473:84]
  wire [7:0] _GEN_3420 = _GEN_8658 == 8'h2a ? _GEN_3416 : _GEN_2992; // @[executor.scala 473:84]
  wire [7:0] _GEN_3421 = _GEN_8658 == 8'h2a ? _GEN_3417 : _GEN_2993; // @[executor.scala 473:84]
  wire [7:0] _GEN_3422 = mask_3[0] ? byte_768 : _GEN_2994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3423 = mask_3[1] ? byte_769 : _GEN_2995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3424 = mask_3[2] ? byte_770 : _GEN_2996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3425 = mask_3[3] ? byte_771 : _GEN_2997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3426 = _GEN_8658 == 8'h2b ? _GEN_3422 : _GEN_2994; // @[executor.scala 473:84]
  wire [7:0] _GEN_3427 = _GEN_8658 == 8'h2b ? _GEN_3423 : _GEN_2995; // @[executor.scala 473:84]
  wire [7:0] _GEN_3428 = _GEN_8658 == 8'h2b ? _GEN_3424 : _GEN_2996; // @[executor.scala 473:84]
  wire [7:0] _GEN_3429 = _GEN_8658 == 8'h2b ? _GEN_3425 : _GEN_2997; // @[executor.scala 473:84]
  wire [7:0] _GEN_3430 = mask_3[0] ? byte_768 : _GEN_2998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3431 = mask_3[1] ? byte_769 : _GEN_2999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3432 = mask_3[2] ? byte_770 : _GEN_3000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3433 = mask_3[3] ? byte_771 : _GEN_3001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3434 = _GEN_8658 == 8'h2c ? _GEN_3430 : _GEN_2998; // @[executor.scala 473:84]
  wire [7:0] _GEN_3435 = _GEN_8658 == 8'h2c ? _GEN_3431 : _GEN_2999; // @[executor.scala 473:84]
  wire [7:0] _GEN_3436 = _GEN_8658 == 8'h2c ? _GEN_3432 : _GEN_3000; // @[executor.scala 473:84]
  wire [7:0] _GEN_3437 = _GEN_8658 == 8'h2c ? _GEN_3433 : _GEN_3001; // @[executor.scala 473:84]
  wire [7:0] _GEN_3438 = mask_3[0] ? byte_768 : _GEN_3002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3439 = mask_3[1] ? byte_769 : _GEN_3003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3440 = mask_3[2] ? byte_770 : _GEN_3004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3441 = mask_3[3] ? byte_771 : _GEN_3005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3442 = _GEN_8658 == 8'h2d ? _GEN_3438 : _GEN_3002; // @[executor.scala 473:84]
  wire [7:0] _GEN_3443 = _GEN_8658 == 8'h2d ? _GEN_3439 : _GEN_3003; // @[executor.scala 473:84]
  wire [7:0] _GEN_3444 = _GEN_8658 == 8'h2d ? _GEN_3440 : _GEN_3004; // @[executor.scala 473:84]
  wire [7:0] _GEN_3445 = _GEN_8658 == 8'h2d ? _GEN_3441 : _GEN_3005; // @[executor.scala 473:84]
  wire [7:0] _GEN_3446 = mask_3[0] ? byte_768 : _GEN_3006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3447 = mask_3[1] ? byte_769 : _GEN_3007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3448 = mask_3[2] ? byte_770 : _GEN_3008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3449 = mask_3[3] ? byte_771 : _GEN_3009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3450 = _GEN_8658 == 8'h2e ? _GEN_3446 : _GEN_3006; // @[executor.scala 473:84]
  wire [7:0] _GEN_3451 = _GEN_8658 == 8'h2e ? _GEN_3447 : _GEN_3007; // @[executor.scala 473:84]
  wire [7:0] _GEN_3452 = _GEN_8658 == 8'h2e ? _GEN_3448 : _GEN_3008; // @[executor.scala 473:84]
  wire [7:0] _GEN_3453 = _GEN_8658 == 8'h2e ? _GEN_3449 : _GEN_3009; // @[executor.scala 473:84]
  wire [7:0] _GEN_3454 = mask_3[0] ? byte_768 : _GEN_3010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3455 = mask_3[1] ? byte_769 : _GEN_3011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3456 = mask_3[2] ? byte_770 : _GEN_3012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3457 = mask_3[3] ? byte_771 : _GEN_3013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3458 = _GEN_8658 == 8'h2f ? _GEN_3454 : _GEN_3010; // @[executor.scala 473:84]
  wire [7:0] _GEN_3459 = _GEN_8658 == 8'h2f ? _GEN_3455 : _GEN_3011; // @[executor.scala 473:84]
  wire [7:0] _GEN_3460 = _GEN_8658 == 8'h2f ? _GEN_3456 : _GEN_3012; // @[executor.scala 473:84]
  wire [7:0] _GEN_3461 = _GEN_8658 == 8'h2f ? _GEN_3457 : _GEN_3013; // @[executor.scala 473:84]
  wire [7:0] _GEN_3462 = mask_3[0] ? byte_768 : _GEN_3014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3463 = mask_3[1] ? byte_769 : _GEN_3015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3464 = mask_3[2] ? byte_770 : _GEN_3016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3465 = mask_3[3] ? byte_771 : _GEN_3017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3466 = _GEN_8658 == 8'h30 ? _GEN_3462 : _GEN_3014; // @[executor.scala 473:84]
  wire [7:0] _GEN_3467 = _GEN_8658 == 8'h30 ? _GEN_3463 : _GEN_3015; // @[executor.scala 473:84]
  wire [7:0] _GEN_3468 = _GEN_8658 == 8'h30 ? _GEN_3464 : _GEN_3016; // @[executor.scala 473:84]
  wire [7:0] _GEN_3469 = _GEN_8658 == 8'h30 ? _GEN_3465 : _GEN_3017; // @[executor.scala 473:84]
  wire [7:0] _GEN_3470 = mask_3[0] ? byte_768 : _GEN_3018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3471 = mask_3[1] ? byte_769 : _GEN_3019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3472 = mask_3[2] ? byte_770 : _GEN_3020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3473 = mask_3[3] ? byte_771 : _GEN_3021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3474 = _GEN_8658 == 8'h31 ? _GEN_3470 : _GEN_3018; // @[executor.scala 473:84]
  wire [7:0] _GEN_3475 = _GEN_8658 == 8'h31 ? _GEN_3471 : _GEN_3019; // @[executor.scala 473:84]
  wire [7:0] _GEN_3476 = _GEN_8658 == 8'h31 ? _GEN_3472 : _GEN_3020; // @[executor.scala 473:84]
  wire [7:0] _GEN_3477 = _GEN_8658 == 8'h31 ? _GEN_3473 : _GEN_3021; // @[executor.scala 473:84]
  wire [7:0] _GEN_3478 = mask_3[0] ? byte_768 : _GEN_3022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3479 = mask_3[1] ? byte_769 : _GEN_3023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3480 = mask_3[2] ? byte_770 : _GEN_3024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3481 = mask_3[3] ? byte_771 : _GEN_3025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3482 = _GEN_8658 == 8'h32 ? _GEN_3478 : _GEN_3022; // @[executor.scala 473:84]
  wire [7:0] _GEN_3483 = _GEN_8658 == 8'h32 ? _GEN_3479 : _GEN_3023; // @[executor.scala 473:84]
  wire [7:0] _GEN_3484 = _GEN_8658 == 8'h32 ? _GEN_3480 : _GEN_3024; // @[executor.scala 473:84]
  wire [7:0] _GEN_3485 = _GEN_8658 == 8'h32 ? _GEN_3481 : _GEN_3025; // @[executor.scala 473:84]
  wire [7:0] _GEN_3486 = mask_3[0] ? byte_768 : _GEN_3026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3487 = mask_3[1] ? byte_769 : _GEN_3027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3488 = mask_3[2] ? byte_770 : _GEN_3028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3489 = mask_3[3] ? byte_771 : _GEN_3029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3490 = _GEN_8658 == 8'h33 ? _GEN_3486 : _GEN_3026; // @[executor.scala 473:84]
  wire [7:0] _GEN_3491 = _GEN_8658 == 8'h33 ? _GEN_3487 : _GEN_3027; // @[executor.scala 473:84]
  wire [7:0] _GEN_3492 = _GEN_8658 == 8'h33 ? _GEN_3488 : _GEN_3028; // @[executor.scala 473:84]
  wire [7:0] _GEN_3493 = _GEN_8658 == 8'h33 ? _GEN_3489 : _GEN_3029; // @[executor.scala 473:84]
  wire [7:0] _GEN_3494 = mask_3[0] ? byte_768 : _GEN_3030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3495 = mask_3[1] ? byte_769 : _GEN_3031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3496 = mask_3[2] ? byte_770 : _GEN_3032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3497 = mask_3[3] ? byte_771 : _GEN_3033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3498 = _GEN_8658 == 8'h34 ? _GEN_3494 : _GEN_3030; // @[executor.scala 473:84]
  wire [7:0] _GEN_3499 = _GEN_8658 == 8'h34 ? _GEN_3495 : _GEN_3031; // @[executor.scala 473:84]
  wire [7:0] _GEN_3500 = _GEN_8658 == 8'h34 ? _GEN_3496 : _GEN_3032; // @[executor.scala 473:84]
  wire [7:0] _GEN_3501 = _GEN_8658 == 8'h34 ? _GEN_3497 : _GEN_3033; // @[executor.scala 473:84]
  wire [7:0] _GEN_3502 = mask_3[0] ? byte_768 : _GEN_3034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3503 = mask_3[1] ? byte_769 : _GEN_3035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3504 = mask_3[2] ? byte_770 : _GEN_3036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3505 = mask_3[3] ? byte_771 : _GEN_3037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3506 = _GEN_8658 == 8'h35 ? _GEN_3502 : _GEN_3034; // @[executor.scala 473:84]
  wire [7:0] _GEN_3507 = _GEN_8658 == 8'h35 ? _GEN_3503 : _GEN_3035; // @[executor.scala 473:84]
  wire [7:0] _GEN_3508 = _GEN_8658 == 8'h35 ? _GEN_3504 : _GEN_3036; // @[executor.scala 473:84]
  wire [7:0] _GEN_3509 = _GEN_8658 == 8'h35 ? _GEN_3505 : _GEN_3037; // @[executor.scala 473:84]
  wire [7:0] _GEN_3510 = mask_3[0] ? byte_768 : _GEN_3038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3511 = mask_3[1] ? byte_769 : _GEN_3039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3512 = mask_3[2] ? byte_770 : _GEN_3040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3513 = mask_3[3] ? byte_771 : _GEN_3041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3514 = _GEN_8658 == 8'h36 ? _GEN_3510 : _GEN_3038; // @[executor.scala 473:84]
  wire [7:0] _GEN_3515 = _GEN_8658 == 8'h36 ? _GEN_3511 : _GEN_3039; // @[executor.scala 473:84]
  wire [7:0] _GEN_3516 = _GEN_8658 == 8'h36 ? _GEN_3512 : _GEN_3040; // @[executor.scala 473:84]
  wire [7:0] _GEN_3517 = _GEN_8658 == 8'h36 ? _GEN_3513 : _GEN_3041; // @[executor.scala 473:84]
  wire [7:0] _GEN_3518 = mask_3[0] ? byte_768 : _GEN_3042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3519 = mask_3[1] ? byte_769 : _GEN_3043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3520 = mask_3[2] ? byte_770 : _GEN_3044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3521 = mask_3[3] ? byte_771 : _GEN_3045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3522 = _GEN_8658 == 8'h37 ? _GEN_3518 : _GEN_3042; // @[executor.scala 473:84]
  wire [7:0] _GEN_3523 = _GEN_8658 == 8'h37 ? _GEN_3519 : _GEN_3043; // @[executor.scala 473:84]
  wire [7:0] _GEN_3524 = _GEN_8658 == 8'h37 ? _GEN_3520 : _GEN_3044; // @[executor.scala 473:84]
  wire [7:0] _GEN_3525 = _GEN_8658 == 8'h37 ? _GEN_3521 : _GEN_3045; // @[executor.scala 473:84]
  wire [7:0] _GEN_3526 = mask_3[0] ? byte_768 : _GEN_3046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3527 = mask_3[1] ? byte_769 : _GEN_3047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3528 = mask_3[2] ? byte_770 : _GEN_3048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3529 = mask_3[3] ? byte_771 : _GEN_3049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3530 = _GEN_8658 == 8'h38 ? _GEN_3526 : _GEN_3046; // @[executor.scala 473:84]
  wire [7:0] _GEN_3531 = _GEN_8658 == 8'h38 ? _GEN_3527 : _GEN_3047; // @[executor.scala 473:84]
  wire [7:0] _GEN_3532 = _GEN_8658 == 8'h38 ? _GEN_3528 : _GEN_3048; // @[executor.scala 473:84]
  wire [7:0] _GEN_3533 = _GEN_8658 == 8'h38 ? _GEN_3529 : _GEN_3049; // @[executor.scala 473:84]
  wire [7:0] _GEN_3534 = mask_3[0] ? byte_768 : _GEN_3050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3535 = mask_3[1] ? byte_769 : _GEN_3051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3536 = mask_3[2] ? byte_770 : _GEN_3052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3537 = mask_3[3] ? byte_771 : _GEN_3053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3538 = _GEN_8658 == 8'h39 ? _GEN_3534 : _GEN_3050; // @[executor.scala 473:84]
  wire [7:0] _GEN_3539 = _GEN_8658 == 8'h39 ? _GEN_3535 : _GEN_3051; // @[executor.scala 473:84]
  wire [7:0] _GEN_3540 = _GEN_8658 == 8'h39 ? _GEN_3536 : _GEN_3052; // @[executor.scala 473:84]
  wire [7:0] _GEN_3541 = _GEN_8658 == 8'h39 ? _GEN_3537 : _GEN_3053; // @[executor.scala 473:84]
  wire [7:0] _GEN_3542 = mask_3[0] ? byte_768 : _GEN_3054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3543 = mask_3[1] ? byte_769 : _GEN_3055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3544 = mask_3[2] ? byte_770 : _GEN_3056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3545 = mask_3[3] ? byte_771 : _GEN_3057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3546 = _GEN_8658 == 8'h3a ? _GEN_3542 : _GEN_3054; // @[executor.scala 473:84]
  wire [7:0] _GEN_3547 = _GEN_8658 == 8'h3a ? _GEN_3543 : _GEN_3055; // @[executor.scala 473:84]
  wire [7:0] _GEN_3548 = _GEN_8658 == 8'h3a ? _GEN_3544 : _GEN_3056; // @[executor.scala 473:84]
  wire [7:0] _GEN_3549 = _GEN_8658 == 8'h3a ? _GEN_3545 : _GEN_3057; // @[executor.scala 473:84]
  wire [7:0] _GEN_3550 = mask_3[0] ? byte_768 : _GEN_3058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3551 = mask_3[1] ? byte_769 : _GEN_3059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3552 = mask_3[2] ? byte_770 : _GEN_3060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3553 = mask_3[3] ? byte_771 : _GEN_3061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3554 = _GEN_8658 == 8'h3b ? _GEN_3550 : _GEN_3058; // @[executor.scala 473:84]
  wire [7:0] _GEN_3555 = _GEN_8658 == 8'h3b ? _GEN_3551 : _GEN_3059; // @[executor.scala 473:84]
  wire [7:0] _GEN_3556 = _GEN_8658 == 8'h3b ? _GEN_3552 : _GEN_3060; // @[executor.scala 473:84]
  wire [7:0] _GEN_3557 = _GEN_8658 == 8'h3b ? _GEN_3553 : _GEN_3061; // @[executor.scala 473:84]
  wire [7:0] _GEN_3558 = mask_3[0] ? byte_768 : _GEN_3062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3559 = mask_3[1] ? byte_769 : _GEN_3063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3560 = mask_3[2] ? byte_770 : _GEN_3064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3561 = mask_3[3] ? byte_771 : _GEN_3065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3562 = _GEN_8658 == 8'h3c ? _GEN_3558 : _GEN_3062; // @[executor.scala 473:84]
  wire [7:0] _GEN_3563 = _GEN_8658 == 8'h3c ? _GEN_3559 : _GEN_3063; // @[executor.scala 473:84]
  wire [7:0] _GEN_3564 = _GEN_8658 == 8'h3c ? _GEN_3560 : _GEN_3064; // @[executor.scala 473:84]
  wire [7:0] _GEN_3565 = _GEN_8658 == 8'h3c ? _GEN_3561 : _GEN_3065; // @[executor.scala 473:84]
  wire [7:0] _GEN_3566 = mask_3[0] ? byte_768 : _GEN_3066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3567 = mask_3[1] ? byte_769 : _GEN_3067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3568 = mask_3[2] ? byte_770 : _GEN_3068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3569 = mask_3[3] ? byte_771 : _GEN_3069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3570 = _GEN_8658 == 8'h3d ? _GEN_3566 : _GEN_3066; // @[executor.scala 473:84]
  wire [7:0] _GEN_3571 = _GEN_8658 == 8'h3d ? _GEN_3567 : _GEN_3067; // @[executor.scala 473:84]
  wire [7:0] _GEN_3572 = _GEN_8658 == 8'h3d ? _GEN_3568 : _GEN_3068; // @[executor.scala 473:84]
  wire [7:0] _GEN_3573 = _GEN_8658 == 8'h3d ? _GEN_3569 : _GEN_3069; // @[executor.scala 473:84]
  wire [7:0] _GEN_3574 = mask_3[0] ? byte_768 : _GEN_3070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3575 = mask_3[1] ? byte_769 : _GEN_3071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3576 = mask_3[2] ? byte_770 : _GEN_3072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3577 = mask_3[3] ? byte_771 : _GEN_3073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3578 = _GEN_8658 == 8'h3e ? _GEN_3574 : _GEN_3070; // @[executor.scala 473:84]
  wire [7:0] _GEN_3579 = _GEN_8658 == 8'h3e ? _GEN_3575 : _GEN_3071; // @[executor.scala 473:84]
  wire [7:0] _GEN_3580 = _GEN_8658 == 8'h3e ? _GEN_3576 : _GEN_3072; // @[executor.scala 473:84]
  wire [7:0] _GEN_3581 = _GEN_8658 == 8'h3e ? _GEN_3577 : _GEN_3073; // @[executor.scala 473:84]
  wire [7:0] _GEN_3582 = mask_3[0] ? byte_768 : _GEN_3074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3583 = mask_3[1] ? byte_769 : _GEN_3075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3584 = mask_3[2] ? byte_770 : _GEN_3076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3585 = mask_3[3] ? byte_771 : _GEN_3077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3586 = _GEN_8658 == 8'h3f ? _GEN_3582 : _GEN_3074; // @[executor.scala 473:84]
  wire [7:0] _GEN_3587 = _GEN_8658 == 8'h3f ? _GEN_3583 : _GEN_3075; // @[executor.scala 473:84]
  wire [7:0] _GEN_3588 = _GEN_8658 == 8'h3f ? _GEN_3584 : _GEN_3076; // @[executor.scala 473:84]
  wire [7:0] _GEN_3589 = _GEN_8658 == 8'h3f ? _GEN_3585 : _GEN_3077; // @[executor.scala 473:84]
  wire [7:0] _GEN_3590 = opcode_3 != 4'h0 ? _GEN_3082 : _GEN_2822; // @[executor.scala 470:55]
  wire [7:0] _GEN_3591 = opcode_3 != 4'h0 ? _GEN_3083 : _GEN_2823; // @[executor.scala 470:55]
  wire [7:0] _GEN_3592 = opcode_3 != 4'h0 ? _GEN_3084 : _GEN_2824; // @[executor.scala 470:55]
  wire [7:0] _GEN_3593 = opcode_3 != 4'h0 ? _GEN_3085 : _GEN_2825; // @[executor.scala 470:55]
  wire [7:0] _GEN_3594 = opcode_3 != 4'h0 ? _GEN_3090 : _GEN_2826; // @[executor.scala 470:55]
  wire [7:0] _GEN_3595 = opcode_3 != 4'h0 ? _GEN_3091 : _GEN_2827; // @[executor.scala 470:55]
  wire [7:0] _GEN_3596 = opcode_3 != 4'h0 ? _GEN_3092 : _GEN_2828; // @[executor.scala 470:55]
  wire [7:0] _GEN_3597 = opcode_3 != 4'h0 ? _GEN_3093 : _GEN_2829; // @[executor.scala 470:55]
  wire [7:0] _GEN_3598 = opcode_3 != 4'h0 ? _GEN_3098 : _GEN_2830; // @[executor.scala 470:55]
  wire [7:0] _GEN_3599 = opcode_3 != 4'h0 ? _GEN_3099 : _GEN_2831; // @[executor.scala 470:55]
  wire [7:0] _GEN_3600 = opcode_3 != 4'h0 ? _GEN_3100 : _GEN_2832; // @[executor.scala 470:55]
  wire [7:0] _GEN_3601 = opcode_3 != 4'h0 ? _GEN_3101 : _GEN_2833; // @[executor.scala 470:55]
  wire [7:0] _GEN_3602 = opcode_3 != 4'h0 ? _GEN_3106 : _GEN_2834; // @[executor.scala 470:55]
  wire [7:0] _GEN_3603 = opcode_3 != 4'h0 ? _GEN_3107 : _GEN_2835; // @[executor.scala 470:55]
  wire [7:0] _GEN_3604 = opcode_3 != 4'h0 ? _GEN_3108 : _GEN_2836; // @[executor.scala 470:55]
  wire [7:0] _GEN_3605 = opcode_3 != 4'h0 ? _GEN_3109 : _GEN_2837; // @[executor.scala 470:55]
  wire [7:0] _GEN_3606 = opcode_3 != 4'h0 ? _GEN_3114 : _GEN_2838; // @[executor.scala 470:55]
  wire [7:0] _GEN_3607 = opcode_3 != 4'h0 ? _GEN_3115 : _GEN_2839; // @[executor.scala 470:55]
  wire [7:0] _GEN_3608 = opcode_3 != 4'h0 ? _GEN_3116 : _GEN_2840; // @[executor.scala 470:55]
  wire [7:0] _GEN_3609 = opcode_3 != 4'h0 ? _GEN_3117 : _GEN_2841; // @[executor.scala 470:55]
  wire [7:0] _GEN_3610 = opcode_3 != 4'h0 ? _GEN_3122 : _GEN_2842; // @[executor.scala 470:55]
  wire [7:0] _GEN_3611 = opcode_3 != 4'h0 ? _GEN_3123 : _GEN_2843; // @[executor.scala 470:55]
  wire [7:0] _GEN_3612 = opcode_3 != 4'h0 ? _GEN_3124 : _GEN_2844; // @[executor.scala 470:55]
  wire [7:0] _GEN_3613 = opcode_3 != 4'h0 ? _GEN_3125 : _GEN_2845; // @[executor.scala 470:55]
  wire [7:0] _GEN_3614 = opcode_3 != 4'h0 ? _GEN_3130 : _GEN_2846; // @[executor.scala 470:55]
  wire [7:0] _GEN_3615 = opcode_3 != 4'h0 ? _GEN_3131 : _GEN_2847; // @[executor.scala 470:55]
  wire [7:0] _GEN_3616 = opcode_3 != 4'h0 ? _GEN_3132 : _GEN_2848; // @[executor.scala 470:55]
  wire [7:0] _GEN_3617 = opcode_3 != 4'h0 ? _GEN_3133 : _GEN_2849; // @[executor.scala 470:55]
  wire [7:0] _GEN_3618 = opcode_3 != 4'h0 ? _GEN_3138 : _GEN_2850; // @[executor.scala 470:55]
  wire [7:0] _GEN_3619 = opcode_3 != 4'h0 ? _GEN_3139 : _GEN_2851; // @[executor.scala 470:55]
  wire [7:0] _GEN_3620 = opcode_3 != 4'h0 ? _GEN_3140 : _GEN_2852; // @[executor.scala 470:55]
  wire [7:0] _GEN_3621 = opcode_3 != 4'h0 ? _GEN_3141 : _GEN_2853; // @[executor.scala 470:55]
  wire [7:0] _GEN_3622 = opcode_3 != 4'h0 ? _GEN_3146 : _GEN_2854; // @[executor.scala 470:55]
  wire [7:0] _GEN_3623 = opcode_3 != 4'h0 ? _GEN_3147 : _GEN_2855; // @[executor.scala 470:55]
  wire [7:0] _GEN_3624 = opcode_3 != 4'h0 ? _GEN_3148 : _GEN_2856; // @[executor.scala 470:55]
  wire [7:0] _GEN_3625 = opcode_3 != 4'h0 ? _GEN_3149 : _GEN_2857; // @[executor.scala 470:55]
  wire [7:0] _GEN_3626 = opcode_3 != 4'h0 ? _GEN_3154 : _GEN_2858; // @[executor.scala 470:55]
  wire [7:0] _GEN_3627 = opcode_3 != 4'h0 ? _GEN_3155 : _GEN_2859; // @[executor.scala 470:55]
  wire [7:0] _GEN_3628 = opcode_3 != 4'h0 ? _GEN_3156 : _GEN_2860; // @[executor.scala 470:55]
  wire [7:0] _GEN_3629 = opcode_3 != 4'h0 ? _GEN_3157 : _GEN_2861; // @[executor.scala 470:55]
  wire [7:0] _GEN_3630 = opcode_3 != 4'h0 ? _GEN_3162 : _GEN_2862; // @[executor.scala 470:55]
  wire [7:0] _GEN_3631 = opcode_3 != 4'h0 ? _GEN_3163 : _GEN_2863; // @[executor.scala 470:55]
  wire [7:0] _GEN_3632 = opcode_3 != 4'h0 ? _GEN_3164 : _GEN_2864; // @[executor.scala 470:55]
  wire [7:0] _GEN_3633 = opcode_3 != 4'h0 ? _GEN_3165 : _GEN_2865; // @[executor.scala 470:55]
  wire [7:0] _GEN_3634 = opcode_3 != 4'h0 ? _GEN_3170 : _GEN_2866; // @[executor.scala 470:55]
  wire [7:0] _GEN_3635 = opcode_3 != 4'h0 ? _GEN_3171 : _GEN_2867; // @[executor.scala 470:55]
  wire [7:0] _GEN_3636 = opcode_3 != 4'h0 ? _GEN_3172 : _GEN_2868; // @[executor.scala 470:55]
  wire [7:0] _GEN_3637 = opcode_3 != 4'h0 ? _GEN_3173 : _GEN_2869; // @[executor.scala 470:55]
  wire [7:0] _GEN_3638 = opcode_3 != 4'h0 ? _GEN_3178 : _GEN_2870; // @[executor.scala 470:55]
  wire [7:0] _GEN_3639 = opcode_3 != 4'h0 ? _GEN_3179 : _GEN_2871; // @[executor.scala 470:55]
  wire [7:0] _GEN_3640 = opcode_3 != 4'h0 ? _GEN_3180 : _GEN_2872; // @[executor.scala 470:55]
  wire [7:0] _GEN_3641 = opcode_3 != 4'h0 ? _GEN_3181 : _GEN_2873; // @[executor.scala 470:55]
  wire [7:0] _GEN_3642 = opcode_3 != 4'h0 ? _GEN_3186 : _GEN_2874; // @[executor.scala 470:55]
  wire [7:0] _GEN_3643 = opcode_3 != 4'h0 ? _GEN_3187 : _GEN_2875; // @[executor.scala 470:55]
  wire [7:0] _GEN_3644 = opcode_3 != 4'h0 ? _GEN_3188 : _GEN_2876; // @[executor.scala 470:55]
  wire [7:0] _GEN_3645 = opcode_3 != 4'h0 ? _GEN_3189 : _GEN_2877; // @[executor.scala 470:55]
  wire [7:0] _GEN_3646 = opcode_3 != 4'h0 ? _GEN_3194 : _GEN_2878; // @[executor.scala 470:55]
  wire [7:0] _GEN_3647 = opcode_3 != 4'h0 ? _GEN_3195 : _GEN_2879; // @[executor.scala 470:55]
  wire [7:0] _GEN_3648 = opcode_3 != 4'h0 ? _GEN_3196 : _GEN_2880; // @[executor.scala 470:55]
  wire [7:0] _GEN_3649 = opcode_3 != 4'h0 ? _GEN_3197 : _GEN_2881; // @[executor.scala 470:55]
  wire [7:0] _GEN_3650 = opcode_3 != 4'h0 ? _GEN_3202 : _GEN_2882; // @[executor.scala 470:55]
  wire [7:0] _GEN_3651 = opcode_3 != 4'h0 ? _GEN_3203 : _GEN_2883; // @[executor.scala 470:55]
  wire [7:0] _GEN_3652 = opcode_3 != 4'h0 ? _GEN_3204 : _GEN_2884; // @[executor.scala 470:55]
  wire [7:0] _GEN_3653 = opcode_3 != 4'h0 ? _GEN_3205 : _GEN_2885; // @[executor.scala 470:55]
  wire [7:0] _GEN_3654 = opcode_3 != 4'h0 ? _GEN_3210 : _GEN_2886; // @[executor.scala 470:55]
  wire [7:0] _GEN_3655 = opcode_3 != 4'h0 ? _GEN_3211 : _GEN_2887; // @[executor.scala 470:55]
  wire [7:0] _GEN_3656 = opcode_3 != 4'h0 ? _GEN_3212 : _GEN_2888; // @[executor.scala 470:55]
  wire [7:0] _GEN_3657 = opcode_3 != 4'h0 ? _GEN_3213 : _GEN_2889; // @[executor.scala 470:55]
  wire [7:0] _GEN_3658 = opcode_3 != 4'h0 ? _GEN_3218 : _GEN_2890; // @[executor.scala 470:55]
  wire [7:0] _GEN_3659 = opcode_3 != 4'h0 ? _GEN_3219 : _GEN_2891; // @[executor.scala 470:55]
  wire [7:0] _GEN_3660 = opcode_3 != 4'h0 ? _GEN_3220 : _GEN_2892; // @[executor.scala 470:55]
  wire [7:0] _GEN_3661 = opcode_3 != 4'h0 ? _GEN_3221 : _GEN_2893; // @[executor.scala 470:55]
  wire [7:0] _GEN_3662 = opcode_3 != 4'h0 ? _GEN_3226 : _GEN_2894; // @[executor.scala 470:55]
  wire [7:0] _GEN_3663 = opcode_3 != 4'h0 ? _GEN_3227 : _GEN_2895; // @[executor.scala 470:55]
  wire [7:0] _GEN_3664 = opcode_3 != 4'h0 ? _GEN_3228 : _GEN_2896; // @[executor.scala 470:55]
  wire [7:0] _GEN_3665 = opcode_3 != 4'h0 ? _GEN_3229 : _GEN_2897; // @[executor.scala 470:55]
  wire [7:0] _GEN_3666 = opcode_3 != 4'h0 ? _GEN_3234 : _GEN_2898; // @[executor.scala 470:55]
  wire [7:0] _GEN_3667 = opcode_3 != 4'h0 ? _GEN_3235 : _GEN_2899; // @[executor.scala 470:55]
  wire [7:0] _GEN_3668 = opcode_3 != 4'h0 ? _GEN_3236 : _GEN_2900; // @[executor.scala 470:55]
  wire [7:0] _GEN_3669 = opcode_3 != 4'h0 ? _GEN_3237 : _GEN_2901; // @[executor.scala 470:55]
  wire [7:0] _GEN_3670 = opcode_3 != 4'h0 ? _GEN_3242 : _GEN_2902; // @[executor.scala 470:55]
  wire [7:0] _GEN_3671 = opcode_3 != 4'h0 ? _GEN_3243 : _GEN_2903; // @[executor.scala 470:55]
  wire [7:0] _GEN_3672 = opcode_3 != 4'h0 ? _GEN_3244 : _GEN_2904; // @[executor.scala 470:55]
  wire [7:0] _GEN_3673 = opcode_3 != 4'h0 ? _GEN_3245 : _GEN_2905; // @[executor.scala 470:55]
  wire [7:0] _GEN_3674 = opcode_3 != 4'h0 ? _GEN_3250 : _GEN_2906; // @[executor.scala 470:55]
  wire [7:0] _GEN_3675 = opcode_3 != 4'h0 ? _GEN_3251 : _GEN_2907; // @[executor.scala 470:55]
  wire [7:0] _GEN_3676 = opcode_3 != 4'h0 ? _GEN_3252 : _GEN_2908; // @[executor.scala 470:55]
  wire [7:0] _GEN_3677 = opcode_3 != 4'h0 ? _GEN_3253 : _GEN_2909; // @[executor.scala 470:55]
  wire [7:0] _GEN_3678 = opcode_3 != 4'h0 ? _GEN_3258 : _GEN_2910; // @[executor.scala 470:55]
  wire [7:0] _GEN_3679 = opcode_3 != 4'h0 ? _GEN_3259 : _GEN_2911; // @[executor.scala 470:55]
  wire [7:0] _GEN_3680 = opcode_3 != 4'h0 ? _GEN_3260 : _GEN_2912; // @[executor.scala 470:55]
  wire [7:0] _GEN_3681 = opcode_3 != 4'h0 ? _GEN_3261 : _GEN_2913; // @[executor.scala 470:55]
  wire [7:0] _GEN_3682 = opcode_3 != 4'h0 ? _GEN_3266 : _GEN_2914; // @[executor.scala 470:55]
  wire [7:0] _GEN_3683 = opcode_3 != 4'h0 ? _GEN_3267 : _GEN_2915; // @[executor.scala 470:55]
  wire [7:0] _GEN_3684 = opcode_3 != 4'h0 ? _GEN_3268 : _GEN_2916; // @[executor.scala 470:55]
  wire [7:0] _GEN_3685 = opcode_3 != 4'h0 ? _GEN_3269 : _GEN_2917; // @[executor.scala 470:55]
  wire [7:0] _GEN_3686 = opcode_3 != 4'h0 ? _GEN_3274 : _GEN_2918; // @[executor.scala 470:55]
  wire [7:0] _GEN_3687 = opcode_3 != 4'h0 ? _GEN_3275 : _GEN_2919; // @[executor.scala 470:55]
  wire [7:0] _GEN_3688 = opcode_3 != 4'h0 ? _GEN_3276 : _GEN_2920; // @[executor.scala 470:55]
  wire [7:0] _GEN_3689 = opcode_3 != 4'h0 ? _GEN_3277 : _GEN_2921; // @[executor.scala 470:55]
  wire [7:0] _GEN_3690 = opcode_3 != 4'h0 ? _GEN_3282 : _GEN_2922; // @[executor.scala 470:55]
  wire [7:0] _GEN_3691 = opcode_3 != 4'h0 ? _GEN_3283 : _GEN_2923; // @[executor.scala 470:55]
  wire [7:0] _GEN_3692 = opcode_3 != 4'h0 ? _GEN_3284 : _GEN_2924; // @[executor.scala 470:55]
  wire [7:0] _GEN_3693 = opcode_3 != 4'h0 ? _GEN_3285 : _GEN_2925; // @[executor.scala 470:55]
  wire [7:0] _GEN_3694 = opcode_3 != 4'h0 ? _GEN_3290 : _GEN_2926; // @[executor.scala 470:55]
  wire [7:0] _GEN_3695 = opcode_3 != 4'h0 ? _GEN_3291 : _GEN_2927; // @[executor.scala 470:55]
  wire [7:0] _GEN_3696 = opcode_3 != 4'h0 ? _GEN_3292 : _GEN_2928; // @[executor.scala 470:55]
  wire [7:0] _GEN_3697 = opcode_3 != 4'h0 ? _GEN_3293 : _GEN_2929; // @[executor.scala 470:55]
  wire [7:0] _GEN_3698 = opcode_3 != 4'h0 ? _GEN_3298 : _GEN_2930; // @[executor.scala 470:55]
  wire [7:0] _GEN_3699 = opcode_3 != 4'h0 ? _GEN_3299 : _GEN_2931; // @[executor.scala 470:55]
  wire [7:0] _GEN_3700 = opcode_3 != 4'h0 ? _GEN_3300 : _GEN_2932; // @[executor.scala 470:55]
  wire [7:0] _GEN_3701 = opcode_3 != 4'h0 ? _GEN_3301 : _GEN_2933; // @[executor.scala 470:55]
  wire [7:0] _GEN_3702 = opcode_3 != 4'h0 ? _GEN_3306 : _GEN_2934; // @[executor.scala 470:55]
  wire [7:0] _GEN_3703 = opcode_3 != 4'h0 ? _GEN_3307 : _GEN_2935; // @[executor.scala 470:55]
  wire [7:0] _GEN_3704 = opcode_3 != 4'h0 ? _GEN_3308 : _GEN_2936; // @[executor.scala 470:55]
  wire [7:0] _GEN_3705 = opcode_3 != 4'h0 ? _GEN_3309 : _GEN_2937; // @[executor.scala 470:55]
  wire [7:0] _GEN_3706 = opcode_3 != 4'h0 ? _GEN_3314 : _GEN_2938; // @[executor.scala 470:55]
  wire [7:0] _GEN_3707 = opcode_3 != 4'h0 ? _GEN_3315 : _GEN_2939; // @[executor.scala 470:55]
  wire [7:0] _GEN_3708 = opcode_3 != 4'h0 ? _GEN_3316 : _GEN_2940; // @[executor.scala 470:55]
  wire [7:0] _GEN_3709 = opcode_3 != 4'h0 ? _GEN_3317 : _GEN_2941; // @[executor.scala 470:55]
  wire [7:0] _GEN_3710 = opcode_3 != 4'h0 ? _GEN_3322 : _GEN_2942; // @[executor.scala 470:55]
  wire [7:0] _GEN_3711 = opcode_3 != 4'h0 ? _GEN_3323 : _GEN_2943; // @[executor.scala 470:55]
  wire [7:0] _GEN_3712 = opcode_3 != 4'h0 ? _GEN_3324 : _GEN_2944; // @[executor.scala 470:55]
  wire [7:0] _GEN_3713 = opcode_3 != 4'h0 ? _GEN_3325 : _GEN_2945; // @[executor.scala 470:55]
  wire [7:0] _GEN_3714 = opcode_3 != 4'h0 ? _GEN_3330 : _GEN_2946; // @[executor.scala 470:55]
  wire [7:0] _GEN_3715 = opcode_3 != 4'h0 ? _GEN_3331 : _GEN_2947; // @[executor.scala 470:55]
  wire [7:0] _GEN_3716 = opcode_3 != 4'h0 ? _GEN_3332 : _GEN_2948; // @[executor.scala 470:55]
  wire [7:0] _GEN_3717 = opcode_3 != 4'h0 ? _GEN_3333 : _GEN_2949; // @[executor.scala 470:55]
  wire [7:0] _GEN_3718 = opcode_3 != 4'h0 ? _GEN_3338 : _GEN_2950; // @[executor.scala 470:55]
  wire [7:0] _GEN_3719 = opcode_3 != 4'h0 ? _GEN_3339 : _GEN_2951; // @[executor.scala 470:55]
  wire [7:0] _GEN_3720 = opcode_3 != 4'h0 ? _GEN_3340 : _GEN_2952; // @[executor.scala 470:55]
  wire [7:0] _GEN_3721 = opcode_3 != 4'h0 ? _GEN_3341 : _GEN_2953; // @[executor.scala 470:55]
  wire [7:0] _GEN_3722 = opcode_3 != 4'h0 ? _GEN_3346 : _GEN_2954; // @[executor.scala 470:55]
  wire [7:0] _GEN_3723 = opcode_3 != 4'h0 ? _GEN_3347 : _GEN_2955; // @[executor.scala 470:55]
  wire [7:0] _GEN_3724 = opcode_3 != 4'h0 ? _GEN_3348 : _GEN_2956; // @[executor.scala 470:55]
  wire [7:0] _GEN_3725 = opcode_3 != 4'h0 ? _GEN_3349 : _GEN_2957; // @[executor.scala 470:55]
  wire [7:0] _GEN_3726 = opcode_3 != 4'h0 ? _GEN_3354 : _GEN_2958; // @[executor.scala 470:55]
  wire [7:0] _GEN_3727 = opcode_3 != 4'h0 ? _GEN_3355 : _GEN_2959; // @[executor.scala 470:55]
  wire [7:0] _GEN_3728 = opcode_3 != 4'h0 ? _GEN_3356 : _GEN_2960; // @[executor.scala 470:55]
  wire [7:0] _GEN_3729 = opcode_3 != 4'h0 ? _GEN_3357 : _GEN_2961; // @[executor.scala 470:55]
  wire [7:0] _GEN_3730 = opcode_3 != 4'h0 ? _GEN_3362 : _GEN_2962; // @[executor.scala 470:55]
  wire [7:0] _GEN_3731 = opcode_3 != 4'h0 ? _GEN_3363 : _GEN_2963; // @[executor.scala 470:55]
  wire [7:0] _GEN_3732 = opcode_3 != 4'h0 ? _GEN_3364 : _GEN_2964; // @[executor.scala 470:55]
  wire [7:0] _GEN_3733 = opcode_3 != 4'h0 ? _GEN_3365 : _GEN_2965; // @[executor.scala 470:55]
  wire [7:0] _GEN_3734 = opcode_3 != 4'h0 ? _GEN_3370 : _GEN_2966; // @[executor.scala 470:55]
  wire [7:0] _GEN_3735 = opcode_3 != 4'h0 ? _GEN_3371 : _GEN_2967; // @[executor.scala 470:55]
  wire [7:0] _GEN_3736 = opcode_3 != 4'h0 ? _GEN_3372 : _GEN_2968; // @[executor.scala 470:55]
  wire [7:0] _GEN_3737 = opcode_3 != 4'h0 ? _GEN_3373 : _GEN_2969; // @[executor.scala 470:55]
  wire [7:0] _GEN_3738 = opcode_3 != 4'h0 ? _GEN_3378 : _GEN_2970; // @[executor.scala 470:55]
  wire [7:0] _GEN_3739 = opcode_3 != 4'h0 ? _GEN_3379 : _GEN_2971; // @[executor.scala 470:55]
  wire [7:0] _GEN_3740 = opcode_3 != 4'h0 ? _GEN_3380 : _GEN_2972; // @[executor.scala 470:55]
  wire [7:0] _GEN_3741 = opcode_3 != 4'h0 ? _GEN_3381 : _GEN_2973; // @[executor.scala 470:55]
  wire [7:0] _GEN_3742 = opcode_3 != 4'h0 ? _GEN_3386 : _GEN_2974; // @[executor.scala 470:55]
  wire [7:0] _GEN_3743 = opcode_3 != 4'h0 ? _GEN_3387 : _GEN_2975; // @[executor.scala 470:55]
  wire [7:0] _GEN_3744 = opcode_3 != 4'h0 ? _GEN_3388 : _GEN_2976; // @[executor.scala 470:55]
  wire [7:0] _GEN_3745 = opcode_3 != 4'h0 ? _GEN_3389 : _GEN_2977; // @[executor.scala 470:55]
  wire [7:0] _GEN_3746 = opcode_3 != 4'h0 ? _GEN_3394 : _GEN_2978; // @[executor.scala 470:55]
  wire [7:0] _GEN_3747 = opcode_3 != 4'h0 ? _GEN_3395 : _GEN_2979; // @[executor.scala 470:55]
  wire [7:0] _GEN_3748 = opcode_3 != 4'h0 ? _GEN_3396 : _GEN_2980; // @[executor.scala 470:55]
  wire [7:0] _GEN_3749 = opcode_3 != 4'h0 ? _GEN_3397 : _GEN_2981; // @[executor.scala 470:55]
  wire [7:0] _GEN_3750 = opcode_3 != 4'h0 ? _GEN_3402 : _GEN_2982; // @[executor.scala 470:55]
  wire [7:0] _GEN_3751 = opcode_3 != 4'h0 ? _GEN_3403 : _GEN_2983; // @[executor.scala 470:55]
  wire [7:0] _GEN_3752 = opcode_3 != 4'h0 ? _GEN_3404 : _GEN_2984; // @[executor.scala 470:55]
  wire [7:0] _GEN_3753 = opcode_3 != 4'h0 ? _GEN_3405 : _GEN_2985; // @[executor.scala 470:55]
  wire [7:0] _GEN_3754 = opcode_3 != 4'h0 ? _GEN_3410 : _GEN_2986; // @[executor.scala 470:55]
  wire [7:0] _GEN_3755 = opcode_3 != 4'h0 ? _GEN_3411 : _GEN_2987; // @[executor.scala 470:55]
  wire [7:0] _GEN_3756 = opcode_3 != 4'h0 ? _GEN_3412 : _GEN_2988; // @[executor.scala 470:55]
  wire [7:0] _GEN_3757 = opcode_3 != 4'h0 ? _GEN_3413 : _GEN_2989; // @[executor.scala 470:55]
  wire [7:0] _GEN_3758 = opcode_3 != 4'h0 ? _GEN_3418 : _GEN_2990; // @[executor.scala 470:55]
  wire [7:0] _GEN_3759 = opcode_3 != 4'h0 ? _GEN_3419 : _GEN_2991; // @[executor.scala 470:55]
  wire [7:0] _GEN_3760 = opcode_3 != 4'h0 ? _GEN_3420 : _GEN_2992; // @[executor.scala 470:55]
  wire [7:0] _GEN_3761 = opcode_3 != 4'h0 ? _GEN_3421 : _GEN_2993; // @[executor.scala 470:55]
  wire [7:0] _GEN_3762 = opcode_3 != 4'h0 ? _GEN_3426 : _GEN_2994; // @[executor.scala 470:55]
  wire [7:0] _GEN_3763 = opcode_3 != 4'h0 ? _GEN_3427 : _GEN_2995; // @[executor.scala 470:55]
  wire [7:0] _GEN_3764 = opcode_3 != 4'h0 ? _GEN_3428 : _GEN_2996; // @[executor.scala 470:55]
  wire [7:0] _GEN_3765 = opcode_3 != 4'h0 ? _GEN_3429 : _GEN_2997; // @[executor.scala 470:55]
  wire [7:0] _GEN_3766 = opcode_3 != 4'h0 ? _GEN_3434 : _GEN_2998; // @[executor.scala 470:55]
  wire [7:0] _GEN_3767 = opcode_3 != 4'h0 ? _GEN_3435 : _GEN_2999; // @[executor.scala 470:55]
  wire [7:0] _GEN_3768 = opcode_3 != 4'h0 ? _GEN_3436 : _GEN_3000; // @[executor.scala 470:55]
  wire [7:0] _GEN_3769 = opcode_3 != 4'h0 ? _GEN_3437 : _GEN_3001; // @[executor.scala 470:55]
  wire [7:0] _GEN_3770 = opcode_3 != 4'h0 ? _GEN_3442 : _GEN_3002; // @[executor.scala 470:55]
  wire [7:0] _GEN_3771 = opcode_3 != 4'h0 ? _GEN_3443 : _GEN_3003; // @[executor.scala 470:55]
  wire [7:0] _GEN_3772 = opcode_3 != 4'h0 ? _GEN_3444 : _GEN_3004; // @[executor.scala 470:55]
  wire [7:0] _GEN_3773 = opcode_3 != 4'h0 ? _GEN_3445 : _GEN_3005; // @[executor.scala 470:55]
  wire [7:0] _GEN_3774 = opcode_3 != 4'h0 ? _GEN_3450 : _GEN_3006; // @[executor.scala 470:55]
  wire [7:0] _GEN_3775 = opcode_3 != 4'h0 ? _GEN_3451 : _GEN_3007; // @[executor.scala 470:55]
  wire [7:0] _GEN_3776 = opcode_3 != 4'h0 ? _GEN_3452 : _GEN_3008; // @[executor.scala 470:55]
  wire [7:0] _GEN_3777 = opcode_3 != 4'h0 ? _GEN_3453 : _GEN_3009; // @[executor.scala 470:55]
  wire [7:0] _GEN_3778 = opcode_3 != 4'h0 ? _GEN_3458 : _GEN_3010; // @[executor.scala 470:55]
  wire [7:0] _GEN_3779 = opcode_3 != 4'h0 ? _GEN_3459 : _GEN_3011; // @[executor.scala 470:55]
  wire [7:0] _GEN_3780 = opcode_3 != 4'h0 ? _GEN_3460 : _GEN_3012; // @[executor.scala 470:55]
  wire [7:0] _GEN_3781 = opcode_3 != 4'h0 ? _GEN_3461 : _GEN_3013; // @[executor.scala 470:55]
  wire [7:0] _GEN_3782 = opcode_3 != 4'h0 ? _GEN_3466 : _GEN_3014; // @[executor.scala 470:55]
  wire [7:0] _GEN_3783 = opcode_3 != 4'h0 ? _GEN_3467 : _GEN_3015; // @[executor.scala 470:55]
  wire [7:0] _GEN_3784 = opcode_3 != 4'h0 ? _GEN_3468 : _GEN_3016; // @[executor.scala 470:55]
  wire [7:0] _GEN_3785 = opcode_3 != 4'h0 ? _GEN_3469 : _GEN_3017; // @[executor.scala 470:55]
  wire [7:0] _GEN_3786 = opcode_3 != 4'h0 ? _GEN_3474 : _GEN_3018; // @[executor.scala 470:55]
  wire [7:0] _GEN_3787 = opcode_3 != 4'h0 ? _GEN_3475 : _GEN_3019; // @[executor.scala 470:55]
  wire [7:0] _GEN_3788 = opcode_3 != 4'h0 ? _GEN_3476 : _GEN_3020; // @[executor.scala 470:55]
  wire [7:0] _GEN_3789 = opcode_3 != 4'h0 ? _GEN_3477 : _GEN_3021; // @[executor.scala 470:55]
  wire [7:0] _GEN_3790 = opcode_3 != 4'h0 ? _GEN_3482 : _GEN_3022; // @[executor.scala 470:55]
  wire [7:0] _GEN_3791 = opcode_3 != 4'h0 ? _GEN_3483 : _GEN_3023; // @[executor.scala 470:55]
  wire [7:0] _GEN_3792 = opcode_3 != 4'h0 ? _GEN_3484 : _GEN_3024; // @[executor.scala 470:55]
  wire [7:0] _GEN_3793 = opcode_3 != 4'h0 ? _GEN_3485 : _GEN_3025; // @[executor.scala 470:55]
  wire [7:0] _GEN_3794 = opcode_3 != 4'h0 ? _GEN_3490 : _GEN_3026; // @[executor.scala 470:55]
  wire [7:0] _GEN_3795 = opcode_3 != 4'h0 ? _GEN_3491 : _GEN_3027; // @[executor.scala 470:55]
  wire [7:0] _GEN_3796 = opcode_3 != 4'h0 ? _GEN_3492 : _GEN_3028; // @[executor.scala 470:55]
  wire [7:0] _GEN_3797 = opcode_3 != 4'h0 ? _GEN_3493 : _GEN_3029; // @[executor.scala 470:55]
  wire [7:0] _GEN_3798 = opcode_3 != 4'h0 ? _GEN_3498 : _GEN_3030; // @[executor.scala 470:55]
  wire [7:0] _GEN_3799 = opcode_3 != 4'h0 ? _GEN_3499 : _GEN_3031; // @[executor.scala 470:55]
  wire [7:0] _GEN_3800 = opcode_3 != 4'h0 ? _GEN_3500 : _GEN_3032; // @[executor.scala 470:55]
  wire [7:0] _GEN_3801 = opcode_3 != 4'h0 ? _GEN_3501 : _GEN_3033; // @[executor.scala 470:55]
  wire [7:0] _GEN_3802 = opcode_3 != 4'h0 ? _GEN_3506 : _GEN_3034; // @[executor.scala 470:55]
  wire [7:0] _GEN_3803 = opcode_3 != 4'h0 ? _GEN_3507 : _GEN_3035; // @[executor.scala 470:55]
  wire [7:0] _GEN_3804 = opcode_3 != 4'h0 ? _GEN_3508 : _GEN_3036; // @[executor.scala 470:55]
  wire [7:0] _GEN_3805 = opcode_3 != 4'h0 ? _GEN_3509 : _GEN_3037; // @[executor.scala 470:55]
  wire [7:0] _GEN_3806 = opcode_3 != 4'h0 ? _GEN_3514 : _GEN_3038; // @[executor.scala 470:55]
  wire [7:0] _GEN_3807 = opcode_3 != 4'h0 ? _GEN_3515 : _GEN_3039; // @[executor.scala 470:55]
  wire [7:0] _GEN_3808 = opcode_3 != 4'h0 ? _GEN_3516 : _GEN_3040; // @[executor.scala 470:55]
  wire [7:0] _GEN_3809 = opcode_3 != 4'h0 ? _GEN_3517 : _GEN_3041; // @[executor.scala 470:55]
  wire [7:0] _GEN_3810 = opcode_3 != 4'h0 ? _GEN_3522 : _GEN_3042; // @[executor.scala 470:55]
  wire [7:0] _GEN_3811 = opcode_3 != 4'h0 ? _GEN_3523 : _GEN_3043; // @[executor.scala 470:55]
  wire [7:0] _GEN_3812 = opcode_3 != 4'h0 ? _GEN_3524 : _GEN_3044; // @[executor.scala 470:55]
  wire [7:0] _GEN_3813 = opcode_3 != 4'h0 ? _GEN_3525 : _GEN_3045; // @[executor.scala 470:55]
  wire [7:0] _GEN_3814 = opcode_3 != 4'h0 ? _GEN_3530 : _GEN_3046; // @[executor.scala 470:55]
  wire [7:0] _GEN_3815 = opcode_3 != 4'h0 ? _GEN_3531 : _GEN_3047; // @[executor.scala 470:55]
  wire [7:0] _GEN_3816 = opcode_3 != 4'h0 ? _GEN_3532 : _GEN_3048; // @[executor.scala 470:55]
  wire [7:0] _GEN_3817 = opcode_3 != 4'h0 ? _GEN_3533 : _GEN_3049; // @[executor.scala 470:55]
  wire [7:0] _GEN_3818 = opcode_3 != 4'h0 ? _GEN_3538 : _GEN_3050; // @[executor.scala 470:55]
  wire [7:0] _GEN_3819 = opcode_3 != 4'h0 ? _GEN_3539 : _GEN_3051; // @[executor.scala 470:55]
  wire [7:0] _GEN_3820 = opcode_3 != 4'h0 ? _GEN_3540 : _GEN_3052; // @[executor.scala 470:55]
  wire [7:0] _GEN_3821 = opcode_3 != 4'h0 ? _GEN_3541 : _GEN_3053; // @[executor.scala 470:55]
  wire [7:0] _GEN_3822 = opcode_3 != 4'h0 ? _GEN_3546 : _GEN_3054; // @[executor.scala 470:55]
  wire [7:0] _GEN_3823 = opcode_3 != 4'h0 ? _GEN_3547 : _GEN_3055; // @[executor.scala 470:55]
  wire [7:0] _GEN_3824 = opcode_3 != 4'h0 ? _GEN_3548 : _GEN_3056; // @[executor.scala 470:55]
  wire [7:0] _GEN_3825 = opcode_3 != 4'h0 ? _GEN_3549 : _GEN_3057; // @[executor.scala 470:55]
  wire [7:0] _GEN_3826 = opcode_3 != 4'h0 ? _GEN_3554 : _GEN_3058; // @[executor.scala 470:55]
  wire [7:0] _GEN_3827 = opcode_3 != 4'h0 ? _GEN_3555 : _GEN_3059; // @[executor.scala 470:55]
  wire [7:0] _GEN_3828 = opcode_3 != 4'h0 ? _GEN_3556 : _GEN_3060; // @[executor.scala 470:55]
  wire [7:0] _GEN_3829 = opcode_3 != 4'h0 ? _GEN_3557 : _GEN_3061; // @[executor.scala 470:55]
  wire [7:0] _GEN_3830 = opcode_3 != 4'h0 ? _GEN_3562 : _GEN_3062; // @[executor.scala 470:55]
  wire [7:0] _GEN_3831 = opcode_3 != 4'h0 ? _GEN_3563 : _GEN_3063; // @[executor.scala 470:55]
  wire [7:0] _GEN_3832 = opcode_3 != 4'h0 ? _GEN_3564 : _GEN_3064; // @[executor.scala 470:55]
  wire [7:0] _GEN_3833 = opcode_3 != 4'h0 ? _GEN_3565 : _GEN_3065; // @[executor.scala 470:55]
  wire [7:0] _GEN_3834 = opcode_3 != 4'h0 ? _GEN_3570 : _GEN_3066; // @[executor.scala 470:55]
  wire [7:0] _GEN_3835 = opcode_3 != 4'h0 ? _GEN_3571 : _GEN_3067; // @[executor.scala 470:55]
  wire [7:0] _GEN_3836 = opcode_3 != 4'h0 ? _GEN_3572 : _GEN_3068; // @[executor.scala 470:55]
  wire [7:0] _GEN_3837 = opcode_3 != 4'h0 ? _GEN_3573 : _GEN_3069; // @[executor.scala 470:55]
  wire [7:0] _GEN_3838 = opcode_3 != 4'h0 ? _GEN_3578 : _GEN_3070; // @[executor.scala 470:55]
  wire [7:0] _GEN_3839 = opcode_3 != 4'h0 ? _GEN_3579 : _GEN_3071; // @[executor.scala 470:55]
  wire [7:0] _GEN_3840 = opcode_3 != 4'h0 ? _GEN_3580 : _GEN_3072; // @[executor.scala 470:55]
  wire [7:0] _GEN_3841 = opcode_3 != 4'h0 ? _GEN_3581 : _GEN_3073; // @[executor.scala 470:55]
  wire [7:0] _GEN_3842 = opcode_3 != 4'h0 ? _GEN_3586 : _GEN_3074; // @[executor.scala 470:55]
  wire [7:0] _GEN_3843 = opcode_3 != 4'h0 ? _GEN_3587 : _GEN_3075; // @[executor.scala 470:55]
  wire [7:0] _GEN_3844 = opcode_3 != 4'h0 ? _GEN_3588 : _GEN_3076; // @[executor.scala 470:55]
  wire [7:0] _GEN_3845 = opcode_3 != 4'h0 ? _GEN_3589 : _GEN_3077; // @[executor.scala 470:55]
  wire [3:0] _GEN_3846 = opcode_3 == 4'hf ? parameter_2_3[13:10] : _GEN_2820; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_3847 = opcode_3 == 4'hf ? parameter_2_3[0] : _GEN_2821; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_3848 = opcode_3 == 4'hf ? _GEN_2822 : _GEN_3590; // @[executor.scala 466:52]
  wire [7:0] _GEN_3849 = opcode_3 == 4'hf ? _GEN_2823 : _GEN_3591; // @[executor.scala 466:52]
  wire [7:0] _GEN_3850 = opcode_3 == 4'hf ? _GEN_2824 : _GEN_3592; // @[executor.scala 466:52]
  wire [7:0] _GEN_3851 = opcode_3 == 4'hf ? _GEN_2825 : _GEN_3593; // @[executor.scala 466:52]
  wire [7:0] _GEN_3852 = opcode_3 == 4'hf ? _GEN_2826 : _GEN_3594; // @[executor.scala 466:52]
  wire [7:0] _GEN_3853 = opcode_3 == 4'hf ? _GEN_2827 : _GEN_3595; // @[executor.scala 466:52]
  wire [7:0] _GEN_3854 = opcode_3 == 4'hf ? _GEN_2828 : _GEN_3596; // @[executor.scala 466:52]
  wire [7:0] _GEN_3855 = opcode_3 == 4'hf ? _GEN_2829 : _GEN_3597; // @[executor.scala 466:52]
  wire [7:0] _GEN_3856 = opcode_3 == 4'hf ? _GEN_2830 : _GEN_3598; // @[executor.scala 466:52]
  wire [7:0] _GEN_3857 = opcode_3 == 4'hf ? _GEN_2831 : _GEN_3599; // @[executor.scala 466:52]
  wire [7:0] _GEN_3858 = opcode_3 == 4'hf ? _GEN_2832 : _GEN_3600; // @[executor.scala 466:52]
  wire [7:0] _GEN_3859 = opcode_3 == 4'hf ? _GEN_2833 : _GEN_3601; // @[executor.scala 466:52]
  wire [7:0] _GEN_3860 = opcode_3 == 4'hf ? _GEN_2834 : _GEN_3602; // @[executor.scala 466:52]
  wire [7:0] _GEN_3861 = opcode_3 == 4'hf ? _GEN_2835 : _GEN_3603; // @[executor.scala 466:52]
  wire [7:0] _GEN_3862 = opcode_3 == 4'hf ? _GEN_2836 : _GEN_3604; // @[executor.scala 466:52]
  wire [7:0] _GEN_3863 = opcode_3 == 4'hf ? _GEN_2837 : _GEN_3605; // @[executor.scala 466:52]
  wire [7:0] _GEN_3864 = opcode_3 == 4'hf ? _GEN_2838 : _GEN_3606; // @[executor.scala 466:52]
  wire [7:0] _GEN_3865 = opcode_3 == 4'hf ? _GEN_2839 : _GEN_3607; // @[executor.scala 466:52]
  wire [7:0] _GEN_3866 = opcode_3 == 4'hf ? _GEN_2840 : _GEN_3608; // @[executor.scala 466:52]
  wire [7:0] _GEN_3867 = opcode_3 == 4'hf ? _GEN_2841 : _GEN_3609; // @[executor.scala 466:52]
  wire [7:0] _GEN_3868 = opcode_3 == 4'hf ? _GEN_2842 : _GEN_3610; // @[executor.scala 466:52]
  wire [7:0] _GEN_3869 = opcode_3 == 4'hf ? _GEN_2843 : _GEN_3611; // @[executor.scala 466:52]
  wire [7:0] _GEN_3870 = opcode_3 == 4'hf ? _GEN_2844 : _GEN_3612; // @[executor.scala 466:52]
  wire [7:0] _GEN_3871 = opcode_3 == 4'hf ? _GEN_2845 : _GEN_3613; // @[executor.scala 466:52]
  wire [7:0] _GEN_3872 = opcode_3 == 4'hf ? _GEN_2846 : _GEN_3614; // @[executor.scala 466:52]
  wire [7:0] _GEN_3873 = opcode_3 == 4'hf ? _GEN_2847 : _GEN_3615; // @[executor.scala 466:52]
  wire [7:0] _GEN_3874 = opcode_3 == 4'hf ? _GEN_2848 : _GEN_3616; // @[executor.scala 466:52]
  wire [7:0] _GEN_3875 = opcode_3 == 4'hf ? _GEN_2849 : _GEN_3617; // @[executor.scala 466:52]
  wire [7:0] _GEN_3876 = opcode_3 == 4'hf ? _GEN_2850 : _GEN_3618; // @[executor.scala 466:52]
  wire [7:0] _GEN_3877 = opcode_3 == 4'hf ? _GEN_2851 : _GEN_3619; // @[executor.scala 466:52]
  wire [7:0] _GEN_3878 = opcode_3 == 4'hf ? _GEN_2852 : _GEN_3620; // @[executor.scala 466:52]
  wire [7:0] _GEN_3879 = opcode_3 == 4'hf ? _GEN_2853 : _GEN_3621; // @[executor.scala 466:52]
  wire [7:0] _GEN_3880 = opcode_3 == 4'hf ? _GEN_2854 : _GEN_3622; // @[executor.scala 466:52]
  wire [7:0] _GEN_3881 = opcode_3 == 4'hf ? _GEN_2855 : _GEN_3623; // @[executor.scala 466:52]
  wire [7:0] _GEN_3882 = opcode_3 == 4'hf ? _GEN_2856 : _GEN_3624; // @[executor.scala 466:52]
  wire [7:0] _GEN_3883 = opcode_3 == 4'hf ? _GEN_2857 : _GEN_3625; // @[executor.scala 466:52]
  wire [7:0] _GEN_3884 = opcode_3 == 4'hf ? _GEN_2858 : _GEN_3626; // @[executor.scala 466:52]
  wire [7:0] _GEN_3885 = opcode_3 == 4'hf ? _GEN_2859 : _GEN_3627; // @[executor.scala 466:52]
  wire [7:0] _GEN_3886 = opcode_3 == 4'hf ? _GEN_2860 : _GEN_3628; // @[executor.scala 466:52]
  wire [7:0] _GEN_3887 = opcode_3 == 4'hf ? _GEN_2861 : _GEN_3629; // @[executor.scala 466:52]
  wire [7:0] _GEN_3888 = opcode_3 == 4'hf ? _GEN_2862 : _GEN_3630; // @[executor.scala 466:52]
  wire [7:0] _GEN_3889 = opcode_3 == 4'hf ? _GEN_2863 : _GEN_3631; // @[executor.scala 466:52]
  wire [7:0] _GEN_3890 = opcode_3 == 4'hf ? _GEN_2864 : _GEN_3632; // @[executor.scala 466:52]
  wire [7:0] _GEN_3891 = opcode_3 == 4'hf ? _GEN_2865 : _GEN_3633; // @[executor.scala 466:52]
  wire [7:0] _GEN_3892 = opcode_3 == 4'hf ? _GEN_2866 : _GEN_3634; // @[executor.scala 466:52]
  wire [7:0] _GEN_3893 = opcode_3 == 4'hf ? _GEN_2867 : _GEN_3635; // @[executor.scala 466:52]
  wire [7:0] _GEN_3894 = opcode_3 == 4'hf ? _GEN_2868 : _GEN_3636; // @[executor.scala 466:52]
  wire [7:0] _GEN_3895 = opcode_3 == 4'hf ? _GEN_2869 : _GEN_3637; // @[executor.scala 466:52]
  wire [7:0] _GEN_3896 = opcode_3 == 4'hf ? _GEN_2870 : _GEN_3638; // @[executor.scala 466:52]
  wire [7:0] _GEN_3897 = opcode_3 == 4'hf ? _GEN_2871 : _GEN_3639; // @[executor.scala 466:52]
  wire [7:0] _GEN_3898 = opcode_3 == 4'hf ? _GEN_2872 : _GEN_3640; // @[executor.scala 466:52]
  wire [7:0] _GEN_3899 = opcode_3 == 4'hf ? _GEN_2873 : _GEN_3641; // @[executor.scala 466:52]
  wire [7:0] _GEN_3900 = opcode_3 == 4'hf ? _GEN_2874 : _GEN_3642; // @[executor.scala 466:52]
  wire [7:0] _GEN_3901 = opcode_3 == 4'hf ? _GEN_2875 : _GEN_3643; // @[executor.scala 466:52]
  wire [7:0] _GEN_3902 = opcode_3 == 4'hf ? _GEN_2876 : _GEN_3644; // @[executor.scala 466:52]
  wire [7:0] _GEN_3903 = opcode_3 == 4'hf ? _GEN_2877 : _GEN_3645; // @[executor.scala 466:52]
  wire [7:0] _GEN_3904 = opcode_3 == 4'hf ? _GEN_2878 : _GEN_3646; // @[executor.scala 466:52]
  wire [7:0] _GEN_3905 = opcode_3 == 4'hf ? _GEN_2879 : _GEN_3647; // @[executor.scala 466:52]
  wire [7:0] _GEN_3906 = opcode_3 == 4'hf ? _GEN_2880 : _GEN_3648; // @[executor.scala 466:52]
  wire [7:0] _GEN_3907 = opcode_3 == 4'hf ? _GEN_2881 : _GEN_3649; // @[executor.scala 466:52]
  wire [7:0] _GEN_3908 = opcode_3 == 4'hf ? _GEN_2882 : _GEN_3650; // @[executor.scala 466:52]
  wire [7:0] _GEN_3909 = opcode_3 == 4'hf ? _GEN_2883 : _GEN_3651; // @[executor.scala 466:52]
  wire [7:0] _GEN_3910 = opcode_3 == 4'hf ? _GEN_2884 : _GEN_3652; // @[executor.scala 466:52]
  wire [7:0] _GEN_3911 = opcode_3 == 4'hf ? _GEN_2885 : _GEN_3653; // @[executor.scala 466:52]
  wire [7:0] _GEN_3912 = opcode_3 == 4'hf ? _GEN_2886 : _GEN_3654; // @[executor.scala 466:52]
  wire [7:0] _GEN_3913 = opcode_3 == 4'hf ? _GEN_2887 : _GEN_3655; // @[executor.scala 466:52]
  wire [7:0] _GEN_3914 = opcode_3 == 4'hf ? _GEN_2888 : _GEN_3656; // @[executor.scala 466:52]
  wire [7:0] _GEN_3915 = opcode_3 == 4'hf ? _GEN_2889 : _GEN_3657; // @[executor.scala 466:52]
  wire [7:0] _GEN_3916 = opcode_3 == 4'hf ? _GEN_2890 : _GEN_3658; // @[executor.scala 466:52]
  wire [7:0] _GEN_3917 = opcode_3 == 4'hf ? _GEN_2891 : _GEN_3659; // @[executor.scala 466:52]
  wire [7:0] _GEN_3918 = opcode_3 == 4'hf ? _GEN_2892 : _GEN_3660; // @[executor.scala 466:52]
  wire [7:0] _GEN_3919 = opcode_3 == 4'hf ? _GEN_2893 : _GEN_3661; // @[executor.scala 466:52]
  wire [7:0] _GEN_3920 = opcode_3 == 4'hf ? _GEN_2894 : _GEN_3662; // @[executor.scala 466:52]
  wire [7:0] _GEN_3921 = opcode_3 == 4'hf ? _GEN_2895 : _GEN_3663; // @[executor.scala 466:52]
  wire [7:0] _GEN_3922 = opcode_3 == 4'hf ? _GEN_2896 : _GEN_3664; // @[executor.scala 466:52]
  wire [7:0] _GEN_3923 = opcode_3 == 4'hf ? _GEN_2897 : _GEN_3665; // @[executor.scala 466:52]
  wire [7:0] _GEN_3924 = opcode_3 == 4'hf ? _GEN_2898 : _GEN_3666; // @[executor.scala 466:52]
  wire [7:0] _GEN_3925 = opcode_3 == 4'hf ? _GEN_2899 : _GEN_3667; // @[executor.scala 466:52]
  wire [7:0] _GEN_3926 = opcode_3 == 4'hf ? _GEN_2900 : _GEN_3668; // @[executor.scala 466:52]
  wire [7:0] _GEN_3927 = opcode_3 == 4'hf ? _GEN_2901 : _GEN_3669; // @[executor.scala 466:52]
  wire [7:0] _GEN_3928 = opcode_3 == 4'hf ? _GEN_2902 : _GEN_3670; // @[executor.scala 466:52]
  wire [7:0] _GEN_3929 = opcode_3 == 4'hf ? _GEN_2903 : _GEN_3671; // @[executor.scala 466:52]
  wire [7:0] _GEN_3930 = opcode_3 == 4'hf ? _GEN_2904 : _GEN_3672; // @[executor.scala 466:52]
  wire [7:0] _GEN_3931 = opcode_3 == 4'hf ? _GEN_2905 : _GEN_3673; // @[executor.scala 466:52]
  wire [7:0] _GEN_3932 = opcode_3 == 4'hf ? _GEN_2906 : _GEN_3674; // @[executor.scala 466:52]
  wire [7:0] _GEN_3933 = opcode_3 == 4'hf ? _GEN_2907 : _GEN_3675; // @[executor.scala 466:52]
  wire [7:0] _GEN_3934 = opcode_3 == 4'hf ? _GEN_2908 : _GEN_3676; // @[executor.scala 466:52]
  wire [7:0] _GEN_3935 = opcode_3 == 4'hf ? _GEN_2909 : _GEN_3677; // @[executor.scala 466:52]
  wire [7:0] _GEN_3936 = opcode_3 == 4'hf ? _GEN_2910 : _GEN_3678; // @[executor.scala 466:52]
  wire [7:0] _GEN_3937 = opcode_3 == 4'hf ? _GEN_2911 : _GEN_3679; // @[executor.scala 466:52]
  wire [7:0] _GEN_3938 = opcode_3 == 4'hf ? _GEN_2912 : _GEN_3680; // @[executor.scala 466:52]
  wire [7:0] _GEN_3939 = opcode_3 == 4'hf ? _GEN_2913 : _GEN_3681; // @[executor.scala 466:52]
  wire [7:0] _GEN_3940 = opcode_3 == 4'hf ? _GEN_2914 : _GEN_3682; // @[executor.scala 466:52]
  wire [7:0] _GEN_3941 = opcode_3 == 4'hf ? _GEN_2915 : _GEN_3683; // @[executor.scala 466:52]
  wire [7:0] _GEN_3942 = opcode_3 == 4'hf ? _GEN_2916 : _GEN_3684; // @[executor.scala 466:52]
  wire [7:0] _GEN_3943 = opcode_3 == 4'hf ? _GEN_2917 : _GEN_3685; // @[executor.scala 466:52]
  wire [7:0] _GEN_3944 = opcode_3 == 4'hf ? _GEN_2918 : _GEN_3686; // @[executor.scala 466:52]
  wire [7:0] _GEN_3945 = opcode_3 == 4'hf ? _GEN_2919 : _GEN_3687; // @[executor.scala 466:52]
  wire [7:0] _GEN_3946 = opcode_3 == 4'hf ? _GEN_2920 : _GEN_3688; // @[executor.scala 466:52]
  wire [7:0] _GEN_3947 = opcode_3 == 4'hf ? _GEN_2921 : _GEN_3689; // @[executor.scala 466:52]
  wire [7:0] _GEN_3948 = opcode_3 == 4'hf ? _GEN_2922 : _GEN_3690; // @[executor.scala 466:52]
  wire [7:0] _GEN_3949 = opcode_3 == 4'hf ? _GEN_2923 : _GEN_3691; // @[executor.scala 466:52]
  wire [7:0] _GEN_3950 = opcode_3 == 4'hf ? _GEN_2924 : _GEN_3692; // @[executor.scala 466:52]
  wire [7:0] _GEN_3951 = opcode_3 == 4'hf ? _GEN_2925 : _GEN_3693; // @[executor.scala 466:52]
  wire [7:0] _GEN_3952 = opcode_3 == 4'hf ? _GEN_2926 : _GEN_3694; // @[executor.scala 466:52]
  wire [7:0] _GEN_3953 = opcode_3 == 4'hf ? _GEN_2927 : _GEN_3695; // @[executor.scala 466:52]
  wire [7:0] _GEN_3954 = opcode_3 == 4'hf ? _GEN_2928 : _GEN_3696; // @[executor.scala 466:52]
  wire [7:0] _GEN_3955 = opcode_3 == 4'hf ? _GEN_2929 : _GEN_3697; // @[executor.scala 466:52]
  wire [7:0] _GEN_3956 = opcode_3 == 4'hf ? _GEN_2930 : _GEN_3698; // @[executor.scala 466:52]
  wire [7:0] _GEN_3957 = opcode_3 == 4'hf ? _GEN_2931 : _GEN_3699; // @[executor.scala 466:52]
  wire [7:0] _GEN_3958 = opcode_3 == 4'hf ? _GEN_2932 : _GEN_3700; // @[executor.scala 466:52]
  wire [7:0] _GEN_3959 = opcode_3 == 4'hf ? _GEN_2933 : _GEN_3701; // @[executor.scala 466:52]
  wire [7:0] _GEN_3960 = opcode_3 == 4'hf ? _GEN_2934 : _GEN_3702; // @[executor.scala 466:52]
  wire [7:0] _GEN_3961 = opcode_3 == 4'hf ? _GEN_2935 : _GEN_3703; // @[executor.scala 466:52]
  wire [7:0] _GEN_3962 = opcode_3 == 4'hf ? _GEN_2936 : _GEN_3704; // @[executor.scala 466:52]
  wire [7:0] _GEN_3963 = opcode_3 == 4'hf ? _GEN_2937 : _GEN_3705; // @[executor.scala 466:52]
  wire [7:0] _GEN_3964 = opcode_3 == 4'hf ? _GEN_2938 : _GEN_3706; // @[executor.scala 466:52]
  wire [7:0] _GEN_3965 = opcode_3 == 4'hf ? _GEN_2939 : _GEN_3707; // @[executor.scala 466:52]
  wire [7:0] _GEN_3966 = opcode_3 == 4'hf ? _GEN_2940 : _GEN_3708; // @[executor.scala 466:52]
  wire [7:0] _GEN_3967 = opcode_3 == 4'hf ? _GEN_2941 : _GEN_3709; // @[executor.scala 466:52]
  wire [7:0] _GEN_3968 = opcode_3 == 4'hf ? _GEN_2942 : _GEN_3710; // @[executor.scala 466:52]
  wire [7:0] _GEN_3969 = opcode_3 == 4'hf ? _GEN_2943 : _GEN_3711; // @[executor.scala 466:52]
  wire [7:0] _GEN_3970 = opcode_3 == 4'hf ? _GEN_2944 : _GEN_3712; // @[executor.scala 466:52]
  wire [7:0] _GEN_3971 = opcode_3 == 4'hf ? _GEN_2945 : _GEN_3713; // @[executor.scala 466:52]
  wire [7:0] _GEN_3972 = opcode_3 == 4'hf ? _GEN_2946 : _GEN_3714; // @[executor.scala 466:52]
  wire [7:0] _GEN_3973 = opcode_3 == 4'hf ? _GEN_2947 : _GEN_3715; // @[executor.scala 466:52]
  wire [7:0] _GEN_3974 = opcode_3 == 4'hf ? _GEN_2948 : _GEN_3716; // @[executor.scala 466:52]
  wire [7:0] _GEN_3975 = opcode_3 == 4'hf ? _GEN_2949 : _GEN_3717; // @[executor.scala 466:52]
  wire [7:0] _GEN_3976 = opcode_3 == 4'hf ? _GEN_2950 : _GEN_3718; // @[executor.scala 466:52]
  wire [7:0] _GEN_3977 = opcode_3 == 4'hf ? _GEN_2951 : _GEN_3719; // @[executor.scala 466:52]
  wire [7:0] _GEN_3978 = opcode_3 == 4'hf ? _GEN_2952 : _GEN_3720; // @[executor.scala 466:52]
  wire [7:0] _GEN_3979 = opcode_3 == 4'hf ? _GEN_2953 : _GEN_3721; // @[executor.scala 466:52]
  wire [7:0] _GEN_3980 = opcode_3 == 4'hf ? _GEN_2954 : _GEN_3722; // @[executor.scala 466:52]
  wire [7:0] _GEN_3981 = opcode_3 == 4'hf ? _GEN_2955 : _GEN_3723; // @[executor.scala 466:52]
  wire [7:0] _GEN_3982 = opcode_3 == 4'hf ? _GEN_2956 : _GEN_3724; // @[executor.scala 466:52]
  wire [7:0] _GEN_3983 = opcode_3 == 4'hf ? _GEN_2957 : _GEN_3725; // @[executor.scala 466:52]
  wire [7:0] _GEN_3984 = opcode_3 == 4'hf ? _GEN_2958 : _GEN_3726; // @[executor.scala 466:52]
  wire [7:0] _GEN_3985 = opcode_3 == 4'hf ? _GEN_2959 : _GEN_3727; // @[executor.scala 466:52]
  wire [7:0] _GEN_3986 = opcode_3 == 4'hf ? _GEN_2960 : _GEN_3728; // @[executor.scala 466:52]
  wire [7:0] _GEN_3987 = opcode_3 == 4'hf ? _GEN_2961 : _GEN_3729; // @[executor.scala 466:52]
  wire [7:0] _GEN_3988 = opcode_3 == 4'hf ? _GEN_2962 : _GEN_3730; // @[executor.scala 466:52]
  wire [7:0] _GEN_3989 = opcode_3 == 4'hf ? _GEN_2963 : _GEN_3731; // @[executor.scala 466:52]
  wire [7:0] _GEN_3990 = opcode_3 == 4'hf ? _GEN_2964 : _GEN_3732; // @[executor.scala 466:52]
  wire [7:0] _GEN_3991 = opcode_3 == 4'hf ? _GEN_2965 : _GEN_3733; // @[executor.scala 466:52]
  wire [7:0] _GEN_3992 = opcode_3 == 4'hf ? _GEN_2966 : _GEN_3734; // @[executor.scala 466:52]
  wire [7:0] _GEN_3993 = opcode_3 == 4'hf ? _GEN_2967 : _GEN_3735; // @[executor.scala 466:52]
  wire [7:0] _GEN_3994 = opcode_3 == 4'hf ? _GEN_2968 : _GEN_3736; // @[executor.scala 466:52]
  wire [7:0] _GEN_3995 = opcode_3 == 4'hf ? _GEN_2969 : _GEN_3737; // @[executor.scala 466:52]
  wire [7:0] _GEN_3996 = opcode_3 == 4'hf ? _GEN_2970 : _GEN_3738; // @[executor.scala 466:52]
  wire [7:0] _GEN_3997 = opcode_3 == 4'hf ? _GEN_2971 : _GEN_3739; // @[executor.scala 466:52]
  wire [7:0] _GEN_3998 = opcode_3 == 4'hf ? _GEN_2972 : _GEN_3740; // @[executor.scala 466:52]
  wire [7:0] _GEN_3999 = opcode_3 == 4'hf ? _GEN_2973 : _GEN_3741; // @[executor.scala 466:52]
  wire [7:0] _GEN_4000 = opcode_3 == 4'hf ? _GEN_2974 : _GEN_3742; // @[executor.scala 466:52]
  wire [7:0] _GEN_4001 = opcode_3 == 4'hf ? _GEN_2975 : _GEN_3743; // @[executor.scala 466:52]
  wire [7:0] _GEN_4002 = opcode_3 == 4'hf ? _GEN_2976 : _GEN_3744; // @[executor.scala 466:52]
  wire [7:0] _GEN_4003 = opcode_3 == 4'hf ? _GEN_2977 : _GEN_3745; // @[executor.scala 466:52]
  wire [7:0] _GEN_4004 = opcode_3 == 4'hf ? _GEN_2978 : _GEN_3746; // @[executor.scala 466:52]
  wire [7:0] _GEN_4005 = opcode_3 == 4'hf ? _GEN_2979 : _GEN_3747; // @[executor.scala 466:52]
  wire [7:0] _GEN_4006 = opcode_3 == 4'hf ? _GEN_2980 : _GEN_3748; // @[executor.scala 466:52]
  wire [7:0] _GEN_4007 = opcode_3 == 4'hf ? _GEN_2981 : _GEN_3749; // @[executor.scala 466:52]
  wire [7:0] _GEN_4008 = opcode_3 == 4'hf ? _GEN_2982 : _GEN_3750; // @[executor.scala 466:52]
  wire [7:0] _GEN_4009 = opcode_3 == 4'hf ? _GEN_2983 : _GEN_3751; // @[executor.scala 466:52]
  wire [7:0] _GEN_4010 = opcode_3 == 4'hf ? _GEN_2984 : _GEN_3752; // @[executor.scala 466:52]
  wire [7:0] _GEN_4011 = opcode_3 == 4'hf ? _GEN_2985 : _GEN_3753; // @[executor.scala 466:52]
  wire [7:0] _GEN_4012 = opcode_3 == 4'hf ? _GEN_2986 : _GEN_3754; // @[executor.scala 466:52]
  wire [7:0] _GEN_4013 = opcode_3 == 4'hf ? _GEN_2987 : _GEN_3755; // @[executor.scala 466:52]
  wire [7:0] _GEN_4014 = opcode_3 == 4'hf ? _GEN_2988 : _GEN_3756; // @[executor.scala 466:52]
  wire [7:0] _GEN_4015 = opcode_3 == 4'hf ? _GEN_2989 : _GEN_3757; // @[executor.scala 466:52]
  wire [7:0] _GEN_4016 = opcode_3 == 4'hf ? _GEN_2990 : _GEN_3758; // @[executor.scala 466:52]
  wire [7:0] _GEN_4017 = opcode_3 == 4'hf ? _GEN_2991 : _GEN_3759; // @[executor.scala 466:52]
  wire [7:0] _GEN_4018 = opcode_3 == 4'hf ? _GEN_2992 : _GEN_3760; // @[executor.scala 466:52]
  wire [7:0] _GEN_4019 = opcode_3 == 4'hf ? _GEN_2993 : _GEN_3761; // @[executor.scala 466:52]
  wire [7:0] _GEN_4020 = opcode_3 == 4'hf ? _GEN_2994 : _GEN_3762; // @[executor.scala 466:52]
  wire [7:0] _GEN_4021 = opcode_3 == 4'hf ? _GEN_2995 : _GEN_3763; // @[executor.scala 466:52]
  wire [7:0] _GEN_4022 = opcode_3 == 4'hf ? _GEN_2996 : _GEN_3764; // @[executor.scala 466:52]
  wire [7:0] _GEN_4023 = opcode_3 == 4'hf ? _GEN_2997 : _GEN_3765; // @[executor.scala 466:52]
  wire [7:0] _GEN_4024 = opcode_3 == 4'hf ? _GEN_2998 : _GEN_3766; // @[executor.scala 466:52]
  wire [7:0] _GEN_4025 = opcode_3 == 4'hf ? _GEN_2999 : _GEN_3767; // @[executor.scala 466:52]
  wire [7:0] _GEN_4026 = opcode_3 == 4'hf ? _GEN_3000 : _GEN_3768; // @[executor.scala 466:52]
  wire [7:0] _GEN_4027 = opcode_3 == 4'hf ? _GEN_3001 : _GEN_3769; // @[executor.scala 466:52]
  wire [7:0] _GEN_4028 = opcode_3 == 4'hf ? _GEN_3002 : _GEN_3770; // @[executor.scala 466:52]
  wire [7:0] _GEN_4029 = opcode_3 == 4'hf ? _GEN_3003 : _GEN_3771; // @[executor.scala 466:52]
  wire [7:0] _GEN_4030 = opcode_3 == 4'hf ? _GEN_3004 : _GEN_3772; // @[executor.scala 466:52]
  wire [7:0] _GEN_4031 = opcode_3 == 4'hf ? _GEN_3005 : _GEN_3773; // @[executor.scala 466:52]
  wire [7:0] _GEN_4032 = opcode_3 == 4'hf ? _GEN_3006 : _GEN_3774; // @[executor.scala 466:52]
  wire [7:0] _GEN_4033 = opcode_3 == 4'hf ? _GEN_3007 : _GEN_3775; // @[executor.scala 466:52]
  wire [7:0] _GEN_4034 = opcode_3 == 4'hf ? _GEN_3008 : _GEN_3776; // @[executor.scala 466:52]
  wire [7:0] _GEN_4035 = opcode_3 == 4'hf ? _GEN_3009 : _GEN_3777; // @[executor.scala 466:52]
  wire [7:0] _GEN_4036 = opcode_3 == 4'hf ? _GEN_3010 : _GEN_3778; // @[executor.scala 466:52]
  wire [7:0] _GEN_4037 = opcode_3 == 4'hf ? _GEN_3011 : _GEN_3779; // @[executor.scala 466:52]
  wire [7:0] _GEN_4038 = opcode_3 == 4'hf ? _GEN_3012 : _GEN_3780; // @[executor.scala 466:52]
  wire [7:0] _GEN_4039 = opcode_3 == 4'hf ? _GEN_3013 : _GEN_3781; // @[executor.scala 466:52]
  wire [7:0] _GEN_4040 = opcode_3 == 4'hf ? _GEN_3014 : _GEN_3782; // @[executor.scala 466:52]
  wire [7:0] _GEN_4041 = opcode_3 == 4'hf ? _GEN_3015 : _GEN_3783; // @[executor.scala 466:52]
  wire [7:0] _GEN_4042 = opcode_3 == 4'hf ? _GEN_3016 : _GEN_3784; // @[executor.scala 466:52]
  wire [7:0] _GEN_4043 = opcode_3 == 4'hf ? _GEN_3017 : _GEN_3785; // @[executor.scala 466:52]
  wire [7:0] _GEN_4044 = opcode_3 == 4'hf ? _GEN_3018 : _GEN_3786; // @[executor.scala 466:52]
  wire [7:0] _GEN_4045 = opcode_3 == 4'hf ? _GEN_3019 : _GEN_3787; // @[executor.scala 466:52]
  wire [7:0] _GEN_4046 = opcode_3 == 4'hf ? _GEN_3020 : _GEN_3788; // @[executor.scala 466:52]
  wire [7:0] _GEN_4047 = opcode_3 == 4'hf ? _GEN_3021 : _GEN_3789; // @[executor.scala 466:52]
  wire [7:0] _GEN_4048 = opcode_3 == 4'hf ? _GEN_3022 : _GEN_3790; // @[executor.scala 466:52]
  wire [7:0] _GEN_4049 = opcode_3 == 4'hf ? _GEN_3023 : _GEN_3791; // @[executor.scala 466:52]
  wire [7:0] _GEN_4050 = opcode_3 == 4'hf ? _GEN_3024 : _GEN_3792; // @[executor.scala 466:52]
  wire [7:0] _GEN_4051 = opcode_3 == 4'hf ? _GEN_3025 : _GEN_3793; // @[executor.scala 466:52]
  wire [7:0] _GEN_4052 = opcode_3 == 4'hf ? _GEN_3026 : _GEN_3794; // @[executor.scala 466:52]
  wire [7:0] _GEN_4053 = opcode_3 == 4'hf ? _GEN_3027 : _GEN_3795; // @[executor.scala 466:52]
  wire [7:0] _GEN_4054 = opcode_3 == 4'hf ? _GEN_3028 : _GEN_3796; // @[executor.scala 466:52]
  wire [7:0] _GEN_4055 = opcode_3 == 4'hf ? _GEN_3029 : _GEN_3797; // @[executor.scala 466:52]
  wire [7:0] _GEN_4056 = opcode_3 == 4'hf ? _GEN_3030 : _GEN_3798; // @[executor.scala 466:52]
  wire [7:0] _GEN_4057 = opcode_3 == 4'hf ? _GEN_3031 : _GEN_3799; // @[executor.scala 466:52]
  wire [7:0] _GEN_4058 = opcode_3 == 4'hf ? _GEN_3032 : _GEN_3800; // @[executor.scala 466:52]
  wire [7:0] _GEN_4059 = opcode_3 == 4'hf ? _GEN_3033 : _GEN_3801; // @[executor.scala 466:52]
  wire [7:0] _GEN_4060 = opcode_3 == 4'hf ? _GEN_3034 : _GEN_3802; // @[executor.scala 466:52]
  wire [7:0] _GEN_4061 = opcode_3 == 4'hf ? _GEN_3035 : _GEN_3803; // @[executor.scala 466:52]
  wire [7:0] _GEN_4062 = opcode_3 == 4'hf ? _GEN_3036 : _GEN_3804; // @[executor.scala 466:52]
  wire [7:0] _GEN_4063 = opcode_3 == 4'hf ? _GEN_3037 : _GEN_3805; // @[executor.scala 466:52]
  wire [7:0] _GEN_4064 = opcode_3 == 4'hf ? _GEN_3038 : _GEN_3806; // @[executor.scala 466:52]
  wire [7:0] _GEN_4065 = opcode_3 == 4'hf ? _GEN_3039 : _GEN_3807; // @[executor.scala 466:52]
  wire [7:0] _GEN_4066 = opcode_3 == 4'hf ? _GEN_3040 : _GEN_3808; // @[executor.scala 466:52]
  wire [7:0] _GEN_4067 = opcode_3 == 4'hf ? _GEN_3041 : _GEN_3809; // @[executor.scala 466:52]
  wire [7:0] _GEN_4068 = opcode_3 == 4'hf ? _GEN_3042 : _GEN_3810; // @[executor.scala 466:52]
  wire [7:0] _GEN_4069 = opcode_3 == 4'hf ? _GEN_3043 : _GEN_3811; // @[executor.scala 466:52]
  wire [7:0] _GEN_4070 = opcode_3 == 4'hf ? _GEN_3044 : _GEN_3812; // @[executor.scala 466:52]
  wire [7:0] _GEN_4071 = opcode_3 == 4'hf ? _GEN_3045 : _GEN_3813; // @[executor.scala 466:52]
  wire [7:0] _GEN_4072 = opcode_3 == 4'hf ? _GEN_3046 : _GEN_3814; // @[executor.scala 466:52]
  wire [7:0] _GEN_4073 = opcode_3 == 4'hf ? _GEN_3047 : _GEN_3815; // @[executor.scala 466:52]
  wire [7:0] _GEN_4074 = opcode_3 == 4'hf ? _GEN_3048 : _GEN_3816; // @[executor.scala 466:52]
  wire [7:0] _GEN_4075 = opcode_3 == 4'hf ? _GEN_3049 : _GEN_3817; // @[executor.scala 466:52]
  wire [7:0] _GEN_4076 = opcode_3 == 4'hf ? _GEN_3050 : _GEN_3818; // @[executor.scala 466:52]
  wire [7:0] _GEN_4077 = opcode_3 == 4'hf ? _GEN_3051 : _GEN_3819; // @[executor.scala 466:52]
  wire [7:0] _GEN_4078 = opcode_3 == 4'hf ? _GEN_3052 : _GEN_3820; // @[executor.scala 466:52]
  wire [7:0] _GEN_4079 = opcode_3 == 4'hf ? _GEN_3053 : _GEN_3821; // @[executor.scala 466:52]
  wire [7:0] _GEN_4080 = opcode_3 == 4'hf ? _GEN_3054 : _GEN_3822; // @[executor.scala 466:52]
  wire [7:0] _GEN_4081 = opcode_3 == 4'hf ? _GEN_3055 : _GEN_3823; // @[executor.scala 466:52]
  wire [7:0] _GEN_4082 = opcode_3 == 4'hf ? _GEN_3056 : _GEN_3824; // @[executor.scala 466:52]
  wire [7:0] _GEN_4083 = opcode_3 == 4'hf ? _GEN_3057 : _GEN_3825; // @[executor.scala 466:52]
  wire [7:0] _GEN_4084 = opcode_3 == 4'hf ? _GEN_3058 : _GEN_3826; // @[executor.scala 466:52]
  wire [7:0] _GEN_4085 = opcode_3 == 4'hf ? _GEN_3059 : _GEN_3827; // @[executor.scala 466:52]
  wire [7:0] _GEN_4086 = opcode_3 == 4'hf ? _GEN_3060 : _GEN_3828; // @[executor.scala 466:52]
  wire [7:0] _GEN_4087 = opcode_3 == 4'hf ? _GEN_3061 : _GEN_3829; // @[executor.scala 466:52]
  wire [7:0] _GEN_4088 = opcode_3 == 4'hf ? _GEN_3062 : _GEN_3830; // @[executor.scala 466:52]
  wire [7:0] _GEN_4089 = opcode_3 == 4'hf ? _GEN_3063 : _GEN_3831; // @[executor.scala 466:52]
  wire [7:0] _GEN_4090 = opcode_3 == 4'hf ? _GEN_3064 : _GEN_3832; // @[executor.scala 466:52]
  wire [7:0] _GEN_4091 = opcode_3 == 4'hf ? _GEN_3065 : _GEN_3833; // @[executor.scala 466:52]
  wire [7:0] _GEN_4092 = opcode_3 == 4'hf ? _GEN_3066 : _GEN_3834; // @[executor.scala 466:52]
  wire [7:0] _GEN_4093 = opcode_3 == 4'hf ? _GEN_3067 : _GEN_3835; // @[executor.scala 466:52]
  wire [7:0] _GEN_4094 = opcode_3 == 4'hf ? _GEN_3068 : _GEN_3836; // @[executor.scala 466:52]
  wire [7:0] _GEN_4095 = opcode_3 == 4'hf ? _GEN_3069 : _GEN_3837; // @[executor.scala 466:52]
  wire [7:0] _GEN_4096 = opcode_3 == 4'hf ? _GEN_3070 : _GEN_3838; // @[executor.scala 466:52]
  wire [7:0] _GEN_4097 = opcode_3 == 4'hf ? _GEN_3071 : _GEN_3839; // @[executor.scala 466:52]
  wire [7:0] _GEN_4098 = opcode_3 == 4'hf ? _GEN_3072 : _GEN_3840; // @[executor.scala 466:52]
  wire [7:0] _GEN_4099 = opcode_3 == 4'hf ? _GEN_3073 : _GEN_3841; // @[executor.scala 466:52]
  wire [7:0] _GEN_4100 = opcode_3 == 4'hf ? _GEN_3074 : _GEN_3842; // @[executor.scala 466:52]
  wire [7:0] _GEN_4101 = opcode_3 == 4'hf ? _GEN_3075 : _GEN_3843; // @[executor.scala 466:52]
  wire [7:0] _GEN_4102 = opcode_3 == 4'hf ? _GEN_3076 : _GEN_3844; // @[executor.scala 466:52]
  wire [7:0] _GEN_4103 = opcode_3 == 4'hf ? _GEN_3077 : _GEN_3845; // @[executor.scala 466:52]
  wire [3:0] opcode_4 = vliw_4[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_4 = vliw_4[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8722 = {{2'd0}, dst_offset_4}; // @[executor.scala 473:49]
  wire [7:0] byte_1024 = field_4[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4104 = mask_4[0] ? byte_1024 : _GEN_3848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1025 = field_4[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4105 = mask_4[1] ? byte_1025 : _GEN_3849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1026 = field_4[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4106 = mask_4[2] ? byte_1026 : _GEN_3850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1027 = field_4[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4107 = mask_4[3] ? byte_1027 : _GEN_3851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4108 = _GEN_8722 == 8'h0 ? _GEN_4104 : _GEN_3848; // @[executor.scala 473:84]
  wire [7:0] _GEN_4109 = _GEN_8722 == 8'h0 ? _GEN_4105 : _GEN_3849; // @[executor.scala 473:84]
  wire [7:0] _GEN_4110 = _GEN_8722 == 8'h0 ? _GEN_4106 : _GEN_3850; // @[executor.scala 473:84]
  wire [7:0] _GEN_4111 = _GEN_8722 == 8'h0 ? _GEN_4107 : _GEN_3851; // @[executor.scala 473:84]
  wire [7:0] _GEN_4112 = mask_4[0] ? byte_1024 : _GEN_3852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4113 = mask_4[1] ? byte_1025 : _GEN_3853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4114 = mask_4[2] ? byte_1026 : _GEN_3854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4115 = mask_4[3] ? byte_1027 : _GEN_3855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4116 = _GEN_8722 == 8'h1 ? _GEN_4112 : _GEN_3852; // @[executor.scala 473:84]
  wire [7:0] _GEN_4117 = _GEN_8722 == 8'h1 ? _GEN_4113 : _GEN_3853; // @[executor.scala 473:84]
  wire [7:0] _GEN_4118 = _GEN_8722 == 8'h1 ? _GEN_4114 : _GEN_3854; // @[executor.scala 473:84]
  wire [7:0] _GEN_4119 = _GEN_8722 == 8'h1 ? _GEN_4115 : _GEN_3855; // @[executor.scala 473:84]
  wire [7:0] _GEN_4120 = mask_4[0] ? byte_1024 : _GEN_3856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4121 = mask_4[1] ? byte_1025 : _GEN_3857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4122 = mask_4[2] ? byte_1026 : _GEN_3858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4123 = mask_4[3] ? byte_1027 : _GEN_3859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4124 = _GEN_8722 == 8'h2 ? _GEN_4120 : _GEN_3856; // @[executor.scala 473:84]
  wire [7:0] _GEN_4125 = _GEN_8722 == 8'h2 ? _GEN_4121 : _GEN_3857; // @[executor.scala 473:84]
  wire [7:0] _GEN_4126 = _GEN_8722 == 8'h2 ? _GEN_4122 : _GEN_3858; // @[executor.scala 473:84]
  wire [7:0] _GEN_4127 = _GEN_8722 == 8'h2 ? _GEN_4123 : _GEN_3859; // @[executor.scala 473:84]
  wire [7:0] _GEN_4128 = mask_4[0] ? byte_1024 : _GEN_3860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4129 = mask_4[1] ? byte_1025 : _GEN_3861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4130 = mask_4[2] ? byte_1026 : _GEN_3862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4131 = mask_4[3] ? byte_1027 : _GEN_3863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4132 = _GEN_8722 == 8'h3 ? _GEN_4128 : _GEN_3860; // @[executor.scala 473:84]
  wire [7:0] _GEN_4133 = _GEN_8722 == 8'h3 ? _GEN_4129 : _GEN_3861; // @[executor.scala 473:84]
  wire [7:0] _GEN_4134 = _GEN_8722 == 8'h3 ? _GEN_4130 : _GEN_3862; // @[executor.scala 473:84]
  wire [7:0] _GEN_4135 = _GEN_8722 == 8'h3 ? _GEN_4131 : _GEN_3863; // @[executor.scala 473:84]
  wire [7:0] _GEN_4136 = mask_4[0] ? byte_1024 : _GEN_3864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4137 = mask_4[1] ? byte_1025 : _GEN_3865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4138 = mask_4[2] ? byte_1026 : _GEN_3866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4139 = mask_4[3] ? byte_1027 : _GEN_3867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4140 = _GEN_8722 == 8'h4 ? _GEN_4136 : _GEN_3864; // @[executor.scala 473:84]
  wire [7:0] _GEN_4141 = _GEN_8722 == 8'h4 ? _GEN_4137 : _GEN_3865; // @[executor.scala 473:84]
  wire [7:0] _GEN_4142 = _GEN_8722 == 8'h4 ? _GEN_4138 : _GEN_3866; // @[executor.scala 473:84]
  wire [7:0] _GEN_4143 = _GEN_8722 == 8'h4 ? _GEN_4139 : _GEN_3867; // @[executor.scala 473:84]
  wire [7:0] _GEN_4144 = mask_4[0] ? byte_1024 : _GEN_3868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4145 = mask_4[1] ? byte_1025 : _GEN_3869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4146 = mask_4[2] ? byte_1026 : _GEN_3870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4147 = mask_4[3] ? byte_1027 : _GEN_3871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4148 = _GEN_8722 == 8'h5 ? _GEN_4144 : _GEN_3868; // @[executor.scala 473:84]
  wire [7:0] _GEN_4149 = _GEN_8722 == 8'h5 ? _GEN_4145 : _GEN_3869; // @[executor.scala 473:84]
  wire [7:0] _GEN_4150 = _GEN_8722 == 8'h5 ? _GEN_4146 : _GEN_3870; // @[executor.scala 473:84]
  wire [7:0] _GEN_4151 = _GEN_8722 == 8'h5 ? _GEN_4147 : _GEN_3871; // @[executor.scala 473:84]
  wire [7:0] _GEN_4152 = mask_4[0] ? byte_1024 : _GEN_3872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4153 = mask_4[1] ? byte_1025 : _GEN_3873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4154 = mask_4[2] ? byte_1026 : _GEN_3874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4155 = mask_4[3] ? byte_1027 : _GEN_3875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4156 = _GEN_8722 == 8'h6 ? _GEN_4152 : _GEN_3872; // @[executor.scala 473:84]
  wire [7:0] _GEN_4157 = _GEN_8722 == 8'h6 ? _GEN_4153 : _GEN_3873; // @[executor.scala 473:84]
  wire [7:0] _GEN_4158 = _GEN_8722 == 8'h6 ? _GEN_4154 : _GEN_3874; // @[executor.scala 473:84]
  wire [7:0] _GEN_4159 = _GEN_8722 == 8'h6 ? _GEN_4155 : _GEN_3875; // @[executor.scala 473:84]
  wire [7:0] _GEN_4160 = mask_4[0] ? byte_1024 : _GEN_3876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4161 = mask_4[1] ? byte_1025 : _GEN_3877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4162 = mask_4[2] ? byte_1026 : _GEN_3878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4163 = mask_4[3] ? byte_1027 : _GEN_3879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4164 = _GEN_8722 == 8'h7 ? _GEN_4160 : _GEN_3876; // @[executor.scala 473:84]
  wire [7:0] _GEN_4165 = _GEN_8722 == 8'h7 ? _GEN_4161 : _GEN_3877; // @[executor.scala 473:84]
  wire [7:0] _GEN_4166 = _GEN_8722 == 8'h7 ? _GEN_4162 : _GEN_3878; // @[executor.scala 473:84]
  wire [7:0] _GEN_4167 = _GEN_8722 == 8'h7 ? _GEN_4163 : _GEN_3879; // @[executor.scala 473:84]
  wire [7:0] _GEN_4168 = mask_4[0] ? byte_1024 : _GEN_3880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4169 = mask_4[1] ? byte_1025 : _GEN_3881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4170 = mask_4[2] ? byte_1026 : _GEN_3882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4171 = mask_4[3] ? byte_1027 : _GEN_3883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4172 = _GEN_8722 == 8'h8 ? _GEN_4168 : _GEN_3880; // @[executor.scala 473:84]
  wire [7:0] _GEN_4173 = _GEN_8722 == 8'h8 ? _GEN_4169 : _GEN_3881; // @[executor.scala 473:84]
  wire [7:0] _GEN_4174 = _GEN_8722 == 8'h8 ? _GEN_4170 : _GEN_3882; // @[executor.scala 473:84]
  wire [7:0] _GEN_4175 = _GEN_8722 == 8'h8 ? _GEN_4171 : _GEN_3883; // @[executor.scala 473:84]
  wire [7:0] _GEN_4176 = mask_4[0] ? byte_1024 : _GEN_3884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4177 = mask_4[1] ? byte_1025 : _GEN_3885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4178 = mask_4[2] ? byte_1026 : _GEN_3886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4179 = mask_4[3] ? byte_1027 : _GEN_3887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4180 = _GEN_8722 == 8'h9 ? _GEN_4176 : _GEN_3884; // @[executor.scala 473:84]
  wire [7:0] _GEN_4181 = _GEN_8722 == 8'h9 ? _GEN_4177 : _GEN_3885; // @[executor.scala 473:84]
  wire [7:0] _GEN_4182 = _GEN_8722 == 8'h9 ? _GEN_4178 : _GEN_3886; // @[executor.scala 473:84]
  wire [7:0] _GEN_4183 = _GEN_8722 == 8'h9 ? _GEN_4179 : _GEN_3887; // @[executor.scala 473:84]
  wire [7:0] _GEN_4184 = mask_4[0] ? byte_1024 : _GEN_3888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4185 = mask_4[1] ? byte_1025 : _GEN_3889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4186 = mask_4[2] ? byte_1026 : _GEN_3890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4187 = mask_4[3] ? byte_1027 : _GEN_3891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4188 = _GEN_8722 == 8'ha ? _GEN_4184 : _GEN_3888; // @[executor.scala 473:84]
  wire [7:0] _GEN_4189 = _GEN_8722 == 8'ha ? _GEN_4185 : _GEN_3889; // @[executor.scala 473:84]
  wire [7:0] _GEN_4190 = _GEN_8722 == 8'ha ? _GEN_4186 : _GEN_3890; // @[executor.scala 473:84]
  wire [7:0] _GEN_4191 = _GEN_8722 == 8'ha ? _GEN_4187 : _GEN_3891; // @[executor.scala 473:84]
  wire [7:0] _GEN_4192 = mask_4[0] ? byte_1024 : _GEN_3892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4193 = mask_4[1] ? byte_1025 : _GEN_3893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4194 = mask_4[2] ? byte_1026 : _GEN_3894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4195 = mask_4[3] ? byte_1027 : _GEN_3895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4196 = _GEN_8722 == 8'hb ? _GEN_4192 : _GEN_3892; // @[executor.scala 473:84]
  wire [7:0] _GEN_4197 = _GEN_8722 == 8'hb ? _GEN_4193 : _GEN_3893; // @[executor.scala 473:84]
  wire [7:0] _GEN_4198 = _GEN_8722 == 8'hb ? _GEN_4194 : _GEN_3894; // @[executor.scala 473:84]
  wire [7:0] _GEN_4199 = _GEN_8722 == 8'hb ? _GEN_4195 : _GEN_3895; // @[executor.scala 473:84]
  wire [7:0] _GEN_4200 = mask_4[0] ? byte_1024 : _GEN_3896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4201 = mask_4[1] ? byte_1025 : _GEN_3897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4202 = mask_4[2] ? byte_1026 : _GEN_3898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4203 = mask_4[3] ? byte_1027 : _GEN_3899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4204 = _GEN_8722 == 8'hc ? _GEN_4200 : _GEN_3896; // @[executor.scala 473:84]
  wire [7:0] _GEN_4205 = _GEN_8722 == 8'hc ? _GEN_4201 : _GEN_3897; // @[executor.scala 473:84]
  wire [7:0] _GEN_4206 = _GEN_8722 == 8'hc ? _GEN_4202 : _GEN_3898; // @[executor.scala 473:84]
  wire [7:0] _GEN_4207 = _GEN_8722 == 8'hc ? _GEN_4203 : _GEN_3899; // @[executor.scala 473:84]
  wire [7:0] _GEN_4208 = mask_4[0] ? byte_1024 : _GEN_3900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4209 = mask_4[1] ? byte_1025 : _GEN_3901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4210 = mask_4[2] ? byte_1026 : _GEN_3902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4211 = mask_4[3] ? byte_1027 : _GEN_3903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4212 = _GEN_8722 == 8'hd ? _GEN_4208 : _GEN_3900; // @[executor.scala 473:84]
  wire [7:0] _GEN_4213 = _GEN_8722 == 8'hd ? _GEN_4209 : _GEN_3901; // @[executor.scala 473:84]
  wire [7:0] _GEN_4214 = _GEN_8722 == 8'hd ? _GEN_4210 : _GEN_3902; // @[executor.scala 473:84]
  wire [7:0] _GEN_4215 = _GEN_8722 == 8'hd ? _GEN_4211 : _GEN_3903; // @[executor.scala 473:84]
  wire [7:0] _GEN_4216 = mask_4[0] ? byte_1024 : _GEN_3904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4217 = mask_4[1] ? byte_1025 : _GEN_3905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4218 = mask_4[2] ? byte_1026 : _GEN_3906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4219 = mask_4[3] ? byte_1027 : _GEN_3907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4220 = _GEN_8722 == 8'he ? _GEN_4216 : _GEN_3904; // @[executor.scala 473:84]
  wire [7:0] _GEN_4221 = _GEN_8722 == 8'he ? _GEN_4217 : _GEN_3905; // @[executor.scala 473:84]
  wire [7:0] _GEN_4222 = _GEN_8722 == 8'he ? _GEN_4218 : _GEN_3906; // @[executor.scala 473:84]
  wire [7:0] _GEN_4223 = _GEN_8722 == 8'he ? _GEN_4219 : _GEN_3907; // @[executor.scala 473:84]
  wire [7:0] _GEN_4224 = mask_4[0] ? byte_1024 : _GEN_3908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4225 = mask_4[1] ? byte_1025 : _GEN_3909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4226 = mask_4[2] ? byte_1026 : _GEN_3910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4227 = mask_4[3] ? byte_1027 : _GEN_3911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4228 = _GEN_8722 == 8'hf ? _GEN_4224 : _GEN_3908; // @[executor.scala 473:84]
  wire [7:0] _GEN_4229 = _GEN_8722 == 8'hf ? _GEN_4225 : _GEN_3909; // @[executor.scala 473:84]
  wire [7:0] _GEN_4230 = _GEN_8722 == 8'hf ? _GEN_4226 : _GEN_3910; // @[executor.scala 473:84]
  wire [7:0] _GEN_4231 = _GEN_8722 == 8'hf ? _GEN_4227 : _GEN_3911; // @[executor.scala 473:84]
  wire [7:0] _GEN_4232 = mask_4[0] ? byte_1024 : _GEN_3912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4233 = mask_4[1] ? byte_1025 : _GEN_3913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4234 = mask_4[2] ? byte_1026 : _GEN_3914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4235 = mask_4[3] ? byte_1027 : _GEN_3915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4236 = _GEN_8722 == 8'h10 ? _GEN_4232 : _GEN_3912; // @[executor.scala 473:84]
  wire [7:0] _GEN_4237 = _GEN_8722 == 8'h10 ? _GEN_4233 : _GEN_3913; // @[executor.scala 473:84]
  wire [7:0] _GEN_4238 = _GEN_8722 == 8'h10 ? _GEN_4234 : _GEN_3914; // @[executor.scala 473:84]
  wire [7:0] _GEN_4239 = _GEN_8722 == 8'h10 ? _GEN_4235 : _GEN_3915; // @[executor.scala 473:84]
  wire [7:0] _GEN_4240 = mask_4[0] ? byte_1024 : _GEN_3916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4241 = mask_4[1] ? byte_1025 : _GEN_3917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4242 = mask_4[2] ? byte_1026 : _GEN_3918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4243 = mask_4[3] ? byte_1027 : _GEN_3919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4244 = _GEN_8722 == 8'h11 ? _GEN_4240 : _GEN_3916; // @[executor.scala 473:84]
  wire [7:0] _GEN_4245 = _GEN_8722 == 8'h11 ? _GEN_4241 : _GEN_3917; // @[executor.scala 473:84]
  wire [7:0] _GEN_4246 = _GEN_8722 == 8'h11 ? _GEN_4242 : _GEN_3918; // @[executor.scala 473:84]
  wire [7:0] _GEN_4247 = _GEN_8722 == 8'h11 ? _GEN_4243 : _GEN_3919; // @[executor.scala 473:84]
  wire [7:0] _GEN_4248 = mask_4[0] ? byte_1024 : _GEN_3920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4249 = mask_4[1] ? byte_1025 : _GEN_3921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4250 = mask_4[2] ? byte_1026 : _GEN_3922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4251 = mask_4[3] ? byte_1027 : _GEN_3923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4252 = _GEN_8722 == 8'h12 ? _GEN_4248 : _GEN_3920; // @[executor.scala 473:84]
  wire [7:0] _GEN_4253 = _GEN_8722 == 8'h12 ? _GEN_4249 : _GEN_3921; // @[executor.scala 473:84]
  wire [7:0] _GEN_4254 = _GEN_8722 == 8'h12 ? _GEN_4250 : _GEN_3922; // @[executor.scala 473:84]
  wire [7:0] _GEN_4255 = _GEN_8722 == 8'h12 ? _GEN_4251 : _GEN_3923; // @[executor.scala 473:84]
  wire [7:0] _GEN_4256 = mask_4[0] ? byte_1024 : _GEN_3924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4257 = mask_4[1] ? byte_1025 : _GEN_3925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4258 = mask_4[2] ? byte_1026 : _GEN_3926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4259 = mask_4[3] ? byte_1027 : _GEN_3927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4260 = _GEN_8722 == 8'h13 ? _GEN_4256 : _GEN_3924; // @[executor.scala 473:84]
  wire [7:0] _GEN_4261 = _GEN_8722 == 8'h13 ? _GEN_4257 : _GEN_3925; // @[executor.scala 473:84]
  wire [7:0] _GEN_4262 = _GEN_8722 == 8'h13 ? _GEN_4258 : _GEN_3926; // @[executor.scala 473:84]
  wire [7:0] _GEN_4263 = _GEN_8722 == 8'h13 ? _GEN_4259 : _GEN_3927; // @[executor.scala 473:84]
  wire [7:0] _GEN_4264 = mask_4[0] ? byte_1024 : _GEN_3928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4265 = mask_4[1] ? byte_1025 : _GEN_3929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4266 = mask_4[2] ? byte_1026 : _GEN_3930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4267 = mask_4[3] ? byte_1027 : _GEN_3931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4268 = _GEN_8722 == 8'h14 ? _GEN_4264 : _GEN_3928; // @[executor.scala 473:84]
  wire [7:0] _GEN_4269 = _GEN_8722 == 8'h14 ? _GEN_4265 : _GEN_3929; // @[executor.scala 473:84]
  wire [7:0] _GEN_4270 = _GEN_8722 == 8'h14 ? _GEN_4266 : _GEN_3930; // @[executor.scala 473:84]
  wire [7:0] _GEN_4271 = _GEN_8722 == 8'h14 ? _GEN_4267 : _GEN_3931; // @[executor.scala 473:84]
  wire [7:0] _GEN_4272 = mask_4[0] ? byte_1024 : _GEN_3932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4273 = mask_4[1] ? byte_1025 : _GEN_3933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4274 = mask_4[2] ? byte_1026 : _GEN_3934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4275 = mask_4[3] ? byte_1027 : _GEN_3935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4276 = _GEN_8722 == 8'h15 ? _GEN_4272 : _GEN_3932; // @[executor.scala 473:84]
  wire [7:0] _GEN_4277 = _GEN_8722 == 8'h15 ? _GEN_4273 : _GEN_3933; // @[executor.scala 473:84]
  wire [7:0] _GEN_4278 = _GEN_8722 == 8'h15 ? _GEN_4274 : _GEN_3934; // @[executor.scala 473:84]
  wire [7:0] _GEN_4279 = _GEN_8722 == 8'h15 ? _GEN_4275 : _GEN_3935; // @[executor.scala 473:84]
  wire [7:0] _GEN_4280 = mask_4[0] ? byte_1024 : _GEN_3936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4281 = mask_4[1] ? byte_1025 : _GEN_3937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4282 = mask_4[2] ? byte_1026 : _GEN_3938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4283 = mask_4[3] ? byte_1027 : _GEN_3939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4284 = _GEN_8722 == 8'h16 ? _GEN_4280 : _GEN_3936; // @[executor.scala 473:84]
  wire [7:0] _GEN_4285 = _GEN_8722 == 8'h16 ? _GEN_4281 : _GEN_3937; // @[executor.scala 473:84]
  wire [7:0] _GEN_4286 = _GEN_8722 == 8'h16 ? _GEN_4282 : _GEN_3938; // @[executor.scala 473:84]
  wire [7:0] _GEN_4287 = _GEN_8722 == 8'h16 ? _GEN_4283 : _GEN_3939; // @[executor.scala 473:84]
  wire [7:0] _GEN_4288 = mask_4[0] ? byte_1024 : _GEN_3940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4289 = mask_4[1] ? byte_1025 : _GEN_3941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4290 = mask_4[2] ? byte_1026 : _GEN_3942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4291 = mask_4[3] ? byte_1027 : _GEN_3943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4292 = _GEN_8722 == 8'h17 ? _GEN_4288 : _GEN_3940; // @[executor.scala 473:84]
  wire [7:0] _GEN_4293 = _GEN_8722 == 8'h17 ? _GEN_4289 : _GEN_3941; // @[executor.scala 473:84]
  wire [7:0] _GEN_4294 = _GEN_8722 == 8'h17 ? _GEN_4290 : _GEN_3942; // @[executor.scala 473:84]
  wire [7:0] _GEN_4295 = _GEN_8722 == 8'h17 ? _GEN_4291 : _GEN_3943; // @[executor.scala 473:84]
  wire [7:0] _GEN_4296 = mask_4[0] ? byte_1024 : _GEN_3944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4297 = mask_4[1] ? byte_1025 : _GEN_3945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4298 = mask_4[2] ? byte_1026 : _GEN_3946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4299 = mask_4[3] ? byte_1027 : _GEN_3947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4300 = _GEN_8722 == 8'h18 ? _GEN_4296 : _GEN_3944; // @[executor.scala 473:84]
  wire [7:0] _GEN_4301 = _GEN_8722 == 8'h18 ? _GEN_4297 : _GEN_3945; // @[executor.scala 473:84]
  wire [7:0] _GEN_4302 = _GEN_8722 == 8'h18 ? _GEN_4298 : _GEN_3946; // @[executor.scala 473:84]
  wire [7:0] _GEN_4303 = _GEN_8722 == 8'h18 ? _GEN_4299 : _GEN_3947; // @[executor.scala 473:84]
  wire [7:0] _GEN_4304 = mask_4[0] ? byte_1024 : _GEN_3948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4305 = mask_4[1] ? byte_1025 : _GEN_3949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4306 = mask_4[2] ? byte_1026 : _GEN_3950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4307 = mask_4[3] ? byte_1027 : _GEN_3951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4308 = _GEN_8722 == 8'h19 ? _GEN_4304 : _GEN_3948; // @[executor.scala 473:84]
  wire [7:0] _GEN_4309 = _GEN_8722 == 8'h19 ? _GEN_4305 : _GEN_3949; // @[executor.scala 473:84]
  wire [7:0] _GEN_4310 = _GEN_8722 == 8'h19 ? _GEN_4306 : _GEN_3950; // @[executor.scala 473:84]
  wire [7:0] _GEN_4311 = _GEN_8722 == 8'h19 ? _GEN_4307 : _GEN_3951; // @[executor.scala 473:84]
  wire [7:0] _GEN_4312 = mask_4[0] ? byte_1024 : _GEN_3952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4313 = mask_4[1] ? byte_1025 : _GEN_3953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4314 = mask_4[2] ? byte_1026 : _GEN_3954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4315 = mask_4[3] ? byte_1027 : _GEN_3955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4316 = _GEN_8722 == 8'h1a ? _GEN_4312 : _GEN_3952; // @[executor.scala 473:84]
  wire [7:0] _GEN_4317 = _GEN_8722 == 8'h1a ? _GEN_4313 : _GEN_3953; // @[executor.scala 473:84]
  wire [7:0] _GEN_4318 = _GEN_8722 == 8'h1a ? _GEN_4314 : _GEN_3954; // @[executor.scala 473:84]
  wire [7:0] _GEN_4319 = _GEN_8722 == 8'h1a ? _GEN_4315 : _GEN_3955; // @[executor.scala 473:84]
  wire [7:0] _GEN_4320 = mask_4[0] ? byte_1024 : _GEN_3956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4321 = mask_4[1] ? byte_1025 : _GEN_3957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4322 = mask_4[2] ? byte_1026 : _GEN_3958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4323 = mask_4[3] ? byte_1027 : _GEN_3959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4324 = _GEN_8722 == 8'h1b ? _GEN_4320 : _GEN_3956; // @[executor.scala 473:84]
  wire [7:0] _GEN_4325 = _GEN_8722 == 8'h1b ? _GEN_4321 : _GEN_3957; // @[executor.scala 473:84]
  wire [7:0] _GEN_4326 = _GEN_8722 == 8'h1b ? _GEN_4322 : _GEN_3958; // @[executor.scala 473:84]
  wire [7:0] _GEN_4327 = _GEN_8722 == 8'h1b ? _GEN_4323 : _GEN_3959; // @[executor.scala 473:84]
  wire [7:0] _GEN_4328 = mask_4[0] ? byte_1024 : _GEN_3960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4329 = mask_4[1] ? byte_1025 : _GEN_3961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4330 = mask_4[2] ? byte_1026 : _GEN_3962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4331 = mask_4[3] ? byte_1027 : _GEN_3963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4332 = _GEN_8722 == 8'h1c ? _GEN_4328 : _GEN_3960; // @[executor.scala 473:84]
  wire [7:0] _GEN_4333 = _GEN_8722 == 8'h1c ? _GEN_4329 : _GEN_3961; // @[executor.scala 473:84]
  wire [7:0] _GEN_4334 = _GEN_8722 == 8'h1c ? _GEN_4330 : _GEN_3962; // @[executor.scala 473:84]
  wire [7:0] _GEN_4335 = _GEN_8722 == 8'h1c ? _GEN_4331 : _GEN_3963; // @[executor.scala 473:84]
  wire [7:0] _GEN_4336 = mask_4[0] ? byte_1024 : _GEN_3964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4337 = mask_4[1] ? byte_1025 : _GEN_3965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4338 = mask_4[2] ? byte_1026 : _GEN_3966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4339 = mask_4[3] ? byte_1027 : _GEN_3967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4340 = _GEN_8722 == 8'h1d ? _GEN_4336 : _GEN_3964; // @[executor.scala 473:84]
  wire [7:0] _GEN_4341 = _GEN_8722 == 8'h1d ? _GEN_4337 : _GEN_3965; // @[executor.scala 473:84]
  wire [7:0] _GEN_4342 = _GEN_8722 == 8'h1d ? _GEN_4338 : _GEN_3966; // @[executor.scala 473:84]
  wire [7:0] _GEN_4343 = _GEN_8722 == 8'h1d ? _GEN_4339 : _GEN_3967; // @[executor.scala 473:84]
  wire [7:0] _GEN_4344 = mask_4[0] ? byte_1024 : _GEN_3968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4345 = mask_4[1] ? byte_1025 : _GEN_3969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4346 = mask_4[2] ? byte_1026 : _GEN_3970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4347 = mask_4[3] ? byte_1027 : _GEN_3971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4348 = _GEN_8722 == 8'h1e ? _GEN_4344 : _GEN_3968; // @[executor.scala 473:84]
  wire [7:0] _GEN_4349 = _GEN_8722 == 8'h1e ? _GEN_4345 : _GEN_3969; // @[executor.scala 473:84]
  wire [7:0] _GEN_4350 = _GEN_8722 == 8'h1e ? _GEN_4346 : _GEN_3970; // @[executor.scala 473:84]
  wire [7:0] _GEN_4351 = _GEN_8722 == 8'h1e ? _GEN_4347 : _GEN_3971; // @[executor.scala 473:84]
  wire [7:0] _GEN_4352 = mask_4[0] ? byte_1024 : _GEN_3972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4353 = mask_4[1] ? byte_1025 : _GEN_3973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4354 = mask_4[2] ? byte_1026 : _GEN_3974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4355 = mask_4[3] ? byte_1027 : _GEN_3975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4356 = _GEN_8722 == 8'h1f ? _GEN_4352 : _GEN_3972; // @[executor.scala 473:84]
  wire [7:0] _GEN_4357 = _GEN_8722 == 8'h1f ? _GEN_4353 : _GEN_3973; // @[executor.scala 473:84]
  wire [7:0] _GEN_4358 = _GEN_8722 == 8'h1f ? _GEN_4354 : _GEN_3974; // @[executor.scala 473:84]
  wire [7:0] _GEN_4359 = _GEN_8722 == 8'h1f ? _GEN_4355 : _GEN_3975; // @[executor.scala 473:84]
  wire [7:0] _GEN_4360 = mask_4[0] ? byte_1024 : _GEN_3976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4361 = mask_4[1] ? byte_1025 : _GEN_3977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4362 = mask_4[2] ? byte_1026 : _GEN_3978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4363 = mask_4[3] ? byte_1027 : _GEN_3979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4364 = _GEN_8722 == 8'h20 ? _GEN_4360 : _GEN_3976; // @[executor.scala 473:84]
  wire [7:0] _GEN_4365 = _GEN_8722 == 8'h20 ? _GEN_4361 : _GEN_3977; // @[executor.scala 473:84]
  wire [7:0] _GEN_4366 = _GEN_8722 == 8'h20 ? _GEN_4362 : _GEN_3978; // @[executor.scala 473:84]
  wire [7:0] _GEN_4367 = _GEN_8722 == 8'h20 ? _GEN_4363 : _GEN_3979; // @[executor.scala 473:84]
  wire [7:0] _GEN_4368 = mask_4[0] ? byte_1024 : _GEN_3980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4369 = mask_4[1] ? byte_1025 : _GEN_3981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4370 = mask_4[2] ? byte_1026 : _GEN_3982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4371 = mask_4[3] ? byte_1027 : _GEN_3983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4372 = _GEN_8722 == 8'h21 ? _GEN_4368 : _GEN_3980; // @[executor.scala 473:84]
  wire [7:0] _GEN_4373 = _GEN_8722 == 8'h21 ? _GEN_4369 : _GEN_3981; // @[executor.scala 473:84]
  wire [7:0] _GEN_4374 = _GEN_8722 == 8'h21 ? _GEN_4370 : _GEN_3982; // @[executor.scala 473:84]
  wire [7:0] _GEN_4375 = _GEN_8722 == 8'h21 ? _GEN_4371 : _GEN_3983; // @[executor.scala 473:84]
  wire [7:0] _GEN_4376 = mask_4[0] ? byte_1024 : _GEN_3984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4377 = mask_4[1] ? byte_1025 : _GEN_3985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4378 = mask_4[2] ? byte_1026 : _GEN_3986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4379 = mask_4[3] ? byte_1027 : _GEN_3987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4380 = _GEN_8722 == 8'h22 ? _GEN_4376 : _GEN_3984; // @[executor.scala 473:84]
  wire [7:0] _GEN_4381 = _GEN_8722 == 8'h22 ? _GEN_4377 : _GEN_3985; // @[executor.scala 473:84]
  wire [7:0] _GEN_4382 = _GEN_8722 == 8'h22 ? _GEN_4378 : _GEN_3986; // @[executor.scala 473:84]
  wire [7:0] _GEN_4383 = _GEN_8722 == 8'h22 ? _GEN_4379 : _GEN_3987; // @[executor.scala 473:84]
  wire [7:0] _GEN_4384 = mask_4[0] ? byte_1024 : _GEN_3988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4385 = mask_4[1] ? byte_1025 : _GEN_3989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4386 = mask_4[2] ? byte_1026 : _GEN_3990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4387 = mask_4[3] ? byte_1027 : _GEN_3991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4388 = _GEN_8722 == 8'h23 ? _GEN_4384 : _GEN_3988; // @[executor.scala 473:84]
  wire [7:0] _GEN_4389 = _GEN_8722 == 8'h23 ? _GEN_4385 : _GEN_3989; // @[executor.scala 473:84]
  wire [7:0] _GEN_4390 = _GEN_8722 == 8'h23 ? _GEN_4386 : _GEN_3990; // @[executor.scala 473:84]
  wire [7:0] _GEN_4391 = _GEN_8722 == 8'h23 ? _GEN_4387 : _GEN_3991; // @[executor.scala 473:84]
  wire [7:0] _GEN_4392 = mask_4[0] ? byte_1024 : _GEN_3992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4393 = mask_4[1] ? byte_1025 : _GEN_3993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4394 = mask_4[2] ? byte_1026 : _GEN_3994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4395 = mask_4[3] ? byte_1027 : _GEN_3995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4396 = _GEN_8722 == 8'h24 ? _GEN_4392 : _GEN_3992; // @[executor.scala 473:84]
  wire [7:0] _GEN_4397 = _GEN_8722 == 8'h24 ? _GEN_4393 : _GEN_3993; // @[executor.scala 473:84]
  wire [7:0] _GEN_4398 = _GEN_8722 == 8'h24 ? _GEN_4394 : _GEN_3994; // @[executor.scala 473:84]
  wire [7:0] _GEN_4399 = _GEN_8722 == 8'h24 ? _GEN_4395 : _GEN_3995; // @[executor.scala 473:84]
  wire [7:0] _GEN_4400 = mask_4[0] ? byte_1024 : _GEN_3996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4401 = mask_4[1] ? byte_1025 : _GEN_3997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4402 = mask_4[2] ? byte_1026 : _GEN_3998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4403 = mask_4[3] ? byte_1027 : _GEN_3999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4404 = _GEN_8722 == 8'h25 ? _GEN_4400 : _GEN_3996; // @[executor.scala 473:84]
  wire [7:0] _GEN_4405 = _GEN_8722 == 8'h25 ? _GEN_4401 : _GEN_3997; // @[executor.scala 473:84]
  wire [7:0] _GEN_4406 = _GEN_8722 == 8'h25 ? _GEN_4402 : _GEN_3998; // @[executor.scala 473:84]
  wire [7:0] _GEN_4407 = _GEN_8722 == 8'h25 ? _GEN_4403 : _GEN_3999; // @[executor.scala 473:84]
  wire [7:0] _GEN_4408 = mask_4[0] ? byte_1024 : _GEN_4000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4409 = mask_4[1] ? byte_1025 : _GEN_4001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4410 = mask_4[2] ? byte_1026 : _GEN_4002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4411 = mask_4[3] ? byte_1027 : _GEN_4003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4412 = _GEN_8722 == 8'h26 ? _GEN_4408 : _GEN_4000; // @[executor.scala 473:84]
  wire [7:0] _GEN_4413 = _GEN_8722 == 8'h26 ? _GEN_4409 : _GEN_4001; // @[executor.scala 473:84]
  wire [7:0] _GEN_4414 = _GEN_8722 == 8'h26 ? _GEN_4410 : _GEN_4002; // @[executor.scala 473:84]
  wire [7:0] _GEN_4415 = _GEN_8722 == 8'h26 ? _GEN_4411 : _GEN_4003; // @[executor.scala 473:84]
  wire [7:0] _GEN_4416 = mask_4[0] ? byte_1024 : _GEN_4004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4417 = mask_4[1] ? byte_1025 : _GEN_4005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4418 = mask_4[2] ? byte_1026 : _GEN_4006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4419 = mask_4[3] ? byte_1027 : _GEN_4007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4420 = _GEN_8722 == 8'h27 ? _GEN_4416 : _GEN_4004; // @[executor.scala 473:84]
  wire [7:0] _GEN_4421 = _GEN_8722 == 8'h27 ? _GEN_4417 : _GEN_4005; // @[executor.scala 473:84]
  wire [7:0] _GEN_4422 = _GEN_8722 == 8'h27 ? _GEN_4418 : _GEN_4006; // @[executor.scala 473:84]
  wire [7:0] _GEN_4423 = _GEN_8722 == 8'h27 ? _GEN_4419 : _GEN_4007; // @[executor.scala 473:84]
  wire [7:0] _GEN_4424 = mask_4[0] ? byte_1024 : _GEN_4008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4425 = mask_4[1] ? byte_1025 : _GEN_4009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4426 = mask_4[2] ? byte_1026 : _GEN_4010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4427 = mask_4[3] ? byte_1027 : _GEN_4011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4428 = _GEN_8722 == 8'h28 ? _GEN_4424 : _GEN_4008; // @[executor.scala 473:84]
  wire [7:0] _GEN_4429 = _GEN_8722 == 8'h28 ? _GEN_4425 : _GEN_4009; // @[executor.scala 473:84]
  wire [7:0] _GEN_4430 = _GEN_8722 == 8'h28 ? _GEN_4426 : _GEN_4010; // @[executor.scala 473:84]
  wire [7:0] _GEN_4431 = _GEN_8722 == 8'h28 ? _GEN_4427 : _GEN_4011; // @[executor.scala 473:84]
  wire [7:0] _GEN_4432 = mask_4[0] ? byte_1024 : _GEN_4012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4433 = mask_4[1] ? byte_1025 : _GEN_4013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4434 = mask_4[2] ? byte_1026 : _GEN_4014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4435 = mask_4[3] ? byte_1027 : _GEN_4015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4436 = _GEN_8722 == 8'h29 ? _GEN_4432 : _GEN_4012; // @[executor.scala 473:84]
  wire [7:0] _GEN_4437 = _GEN_8722 == 8'h29 ? _GEN_4433 : _GEN_4013; // @[executor.scala 473:84]
  wire [7:0] _GEN_4438 = _GEN_8722 == 8'h29 ? _GEN_4434 : _GEN_4014; // @[executor.scala 473:84]
  wire [7:0] _GEN_4439 = _GEN_8722 == 8'h29 ? _GEN_4435 : _GEN_4015; // @[executor.scala 473:84]
  wire [7:0] _GEN_4440 = mask_4[0] ? byte_1024 : _GEN_4016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4441 = mask_4[1] ? byte_1025 : _GEN_4017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4442 = mask_4[2] ? byte_1026 : _GEN_4018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4443 = mask_4[3] ? byte_1027 : _GEN_4019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4444 = _GEN_8722 == 8'h2a ? _GEN_4440 : _GEN_4016; // @[executor.scala 473:84]
  wire [7:0] _GEN_4445 = _GEN_8722 == 8'h2a ? _GEN_4441 : _GEN_4017; // @[executor.scala 473:84]
  wire [7:0] _GEN_4446 = _GEN_8722 == 8'h2a ? _GEN_4442 : _GEN_4018; // @[executor.scala 473:84]
  wire [7:0] _GEN_4447 = _GEN_8722 == 8'h2a ? _GEN_4443 : _GEN_4019; // @[executor.scala 473:84]
  wire [7:0] _GEN_4448 = mask_4[0] ? byte_1024 : _GEN_4020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4449 = mask_4[1] ? byte_1025 : _GEN_4021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4450 = mask_4[2] ? byte_1026 : _GEN_4022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4451 = mask_4[3] ? byte_1027 : _GEN_4023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4452 = _GEN_8722 == 8'h2b ? _GEN_4448 : _GEN_4020; // @[executor.scala 473:84]
  wire [7:0] _GEN_4453 = _GEN_8722 == 8'h2b ? _GEN_4449 : _GEN_4021; // @[executor.scala 473:84]
  wire [7:0] _GEN_4454 = _GEN_8722 == 8'h2b ? _GEN_4450 : _GEN_4022; // @[executor.scala 473:84]
  wire [7:0] _GEN_4455 = _GEN_8722 == 8'h2b ? _GEN_4451 : _GEN_4023; // @[executor.scala 473:84]
  wire [7:0] _GEN_4456 = mask_4[0] ? byte_1024 : _GEN_4024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4457 = mask_4[1] ? byte_1025 : _GEN_4025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4458 = mask_4[2] ? byte_1026 : _GEN_4026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4459 = mask_4[3] ? byte_1027 : _GEN_4027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4460 = _GEN_8722 == 8'h2c ? _GEN_4456 : _GEN_4024; // @[executor.scala 473:84]
  wire [7:0] _GEN_4461 = _GEN_8722 == 8'h2c ? _GEN_4457 : _GEN_4025; // @[executor.scala 473:84]
  wire [7:0] _GEN_4462 = _GEN_8722 == 8'h2c ? _GEN_4458 : _GEN_4026; // @[executor.scala 473:84]
  wire [7:0] _GEN_4463 = _GEN_8722 == 8'h2c ? _GEN_4459 : _GEN_4027; // @[executor.scala 473:84]
  wire [7:0] _GEN_4464 = mask_4[0] ? byte_1024 : _GEN_4028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4465 = mask_4[1] ? byte_1025 : _GEN_4029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4466 = mask_4[2] ? byte_1026 : _GEN_4030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4467 = mask_4[3] ? byte_1027 : _GEN_4031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4468 = _GEN_8722 == 8'h2d ? _GEN_4464 : _GEN_4028; // @[executor.scala 473:84]
  wire [7:0] _GEN_4469 = _GEN_8722 == 8'h2d ? _GEN_4465 : _GEN_4029; // @[executor.scala 473:84]
  wire [7:0] _GEN_4470 = _GEN_8722 == 8'h2d ? _GEN_4466 : _GEN_4030; // @[executor.scala 473:84]
  wire [7:0] _GEN_4471 = _GEN_8722 == 8'h2d ? _GEN_4467 : _GEN_4031; // @[executor.scala 473:84]
  wire [7:0] _GEN_4472 = mask_4[0] ? byte_1024 : _GEN_4032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4473 = mask_4[1] ? byte_1025 : _GEN_4033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4474 = mask_4[2] ? byte_1026 : _GEN_4034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4475 = mask_4[3] ? byte_1027 : _GEN_4035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4476 = _GEN_8722 == 8'h2e ? _GEN_4472 : _GEN_4032; // @[executor.scala 473:84]
  wire [7:0] _GEN_4477 = _GEN_8722 == 8'h2e ? _GEN_4473 : _GEN_4033; // @[executor.scala 473:84]
  wire [7:0] _GEN_4478 = _GEN_8722 == 8'h2e ? _GEN_4474 : _GEN_4034; // @[executor.scala 473:84]
  wire [7:0] _GEN_4479 = _GEN_8722 == 8'h2e ? _GEN_4475 : _GEN_4035; // @[executor.scala 473:84]
  wire [7:0] _GEN_4480 = mask_4[0] ? byte_1024 : _GEN_4036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4481 = mask_4[1] ? byte_1025 : _GEN_4037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4482 = mask_4[2] ? byte_1026 : _GEN_4038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4483 = mask_4[3] ? byte_1027 : _GEN_4039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4484 = _GEN_8722 == 8'h2f ? _GEN_4480 : _GEN_4036; // @[executor.scala 473:84]
  wire [7:0] _GEN_4485 = _GEN_8722 == 8'h2f ? _GEN_4481 : _GEN_4037; // @[executor.scala 473:84]
  wire [7:0] _GEN_4486 = _GEN_8722 == 8'h2f ? _GEN_4482 : _GEN_4038; // @[executor.scala 473:84]
  wire [7:0] _GEN_4487 = _GEN_8722 == 8'h2f ? _GEN_4483 : _GEN_4039; // @[executor.scala 473:84]
  wire [7:0] _GEN_4488 = mask_4[0] ? byte_1024 : _GEN_4040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4489 = mask_4[1] ? byte_1025 : _GEN_4041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4490 = mask_4[2] ? byte_1026 : _GEN_4042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4491 = mask_4[3] ? byte_1027 : _GEN_4043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4492 = _GEN_8722 == 8'h30 ? _GEN_4488 : _GEN_4040; // @[executor.scala 473:84]
  wire [7:0] _GEN_4493 = _GEN_8722 == 8'h30 ? _GEN_4489 : _GEN_4041; // @[executor.scala 473:84]
  wire [7:0] _GEN_4494 = _GEN_8722 == 8'h30 ? _GEN_4490 : _GEN_4042; // @[executor.scala 473:84]
  wire [7:0] _GEN_4495 = _GEN_8722 == 8'h30 ? _GEN_4491 : _GEN_4043; // @[executor.scala 473:84]
  wire [7:0] _GEN_4496 = mask_4[0] ? byte_1024 : _GEN_4044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4497 = mask_4[1] ? byte_1025 : _GEN_4045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4498 = mask_4[2] ? byte_1026 : _GEN_4046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4499 = mask_4[3] ? byte_1027 : _GEN_4047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4500 = _GEN_8722 == 8'h31 ? _GEN_4496 : _GEN_4044; // @[executor.scala 473:84]
  wire [7:0] _GEN_4501 = _GEN_8722 == 8'h31 ? _GEN_4497 : _GEN_4045; // @[executor.scala 473:84]
  wire [7:0] _GEN_4502 = _GEN_8722 == 8'h31 ? _GEN_4498 : _GEN_4046; // @[executor.scala 473:84]
  wire [7:0] _GEN_4503 = _GEN_8722 == 8'h31 ? _GEN_4499 : _GEN_4047; // @[executor.scala 473:84]
  wire [7:0] _GEN_4504 = mask_4[0] ? byte_1024 : _GEN_4048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4505 = mask_4[1] ? byte_1025 : _GEN_4049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4506 = mask_4[2] ? byte_1026 : _GEN_4050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4507 = mask_4[3] ? byte_1027 : _GEN_4051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4508 = _GEN_8722 == 8'h32 ? _GEN_4504 : _GEN_4048; // @[executor.scala 473:84]
  wire [7:0] _GEN_4509 = _GEN_8722 == 8'h32 ? _GEN_4505 : _GEN_4049; // @[executor.scala 473:84]
  wire [7:0] _GEN_4510 = _GEN_8722 == 8'h32 ? _GEN_4506 : _GEN_4050; // @[executor.scala 473:84]
  wire [7:0] _GEN_4511 = _GEN_8722 == 8'h32 ? _GEN_4507 : _GEN_4051; // @[executor.scala 473:84]
  wire [7:0] _GEN_4512 = mask_4[0] ? byte_1024 : _GEN_4052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4513 = mask_4[1] ? byte_1025 : _GEN_4053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4514 = mask_4[2] ? byte_1026 : _GEN_4054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4515 = mask_4[3] ? byte_1027 : _GEN_4055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4516 = _GEN_8722 == 8'h33 ? _GEN_4512 : _GEN_4052; // @[executor.scala 473:84]
  wire [7:0] _GEN_4517 = _GEN_8722 == 8'h33 ? _GEN_4513 : _GEN_4053; // @[executor.scala 473:84]
  wire [7:0] _GEN_4518 = _GEN_8722 == 8'h33 ? _GEN_4514 : _GEN_4054; // @[executor.scala 473:84]
  wire [7:0] _GEN_4519 = _GEN_8722 == 8'h33 ? _GEN_4515 : _GEN_4055; // @[executor.scala 473:84]
  wire [7:0] _GEN_4520 = mask_4[0] ? byte_1024 : _GEN_4056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4521 = mask_4[1] ? byte_1025 : _GEN_4057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4522 = mask_4[2] ? byte_1026 : _GEN_4058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4523 = mask_4[3] ? byte_1027 : _GEN_4059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4524 = _GEN_8722 == 8'h34 ? _GEN_4520 : _GEN_4056; // @[executor.scala 473:84]
  wire [7:0] _GEN_4525 = _GEN_8722 == 8'h34 ? _GEN_4521 : _GEN_4057; // @[executor.scala 473:84]
  wire [7:0] _GEN_4526 = _GEN_8722 == 8'h34 ? _GEN_4522 : _GEN_4058; // @[executor.scala 473:84]
  wire [7:0] _GEN_4527 = _GEN_8722 == 8'h34 ? _GEN_4523 : _GEN_4059; // @[executor.scala 473:84]
  wire [7:0] _GEN_4528 = mask_4[0] ? byte_1024 : _GEN_4060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4529 = mask_4[1] ? byte_1025 : _GEN_4061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4530 = mask_4[2] ? byte_1026 : _GEN_4062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4531 = mask_4[3] ? byte_1027 : _GEN_4063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4532 = _GEN_8722 == 8'h35 ? _GEN_4528 : _GEN_4060; // @[executor.scala 473:84]
  wire [7:0] _GEN_4533 = _GEN_8722 == 8'h35 ? _GEN_4529 : _GEN_4061; // @[executor.scala 473:84]
  wire [7:0] _GEN_4534 = _GEN_8722 == 8'h35 ? _GEN_4530 : _GEN_4062; // @[executor.scala 473:84]
  wire [7:0] _GEN_4535 = _GEN_8722 == 8'h35 ? _GEN_4531 : _GEN_4063; // @[executor.scala 473:84]
  wire [7:0] _GEN_4536 = mask_4[0] ? byte_1024 : _GEN_4064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4537 = mask_4[1] ? byte_1025 : _GEN_4065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4538 = mask_4[2] ? byte_1026 : _GEN_4066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4539 = mask_4[3] ? byte_1027 : _GEN_4067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4540 = _GEN_8722 == 8'h36 ? _GEN_4536 : _GEN_4064; // @[executor.scala 473:84]
  wire [7:0] _GEN_4541 = _GEN_8722 == 8'h36 ? _GEN_4537 : _GEN_4065; // @[executor.scala 473:84]
  wire [7:0] _GEN_4542 = _GEN_8722 == 8'h36 ? _GEN_4538 : _GEN_4066; // @[executor.scala 473:84]
  wire [7:0] _GEN_4543 = _GEN_8722 == 8'h36 ? _GEN_4539 : _GEN_4067; // @[executor.scala 473:84]
  wire [7:0] _GEN_4544 = mask_4[0] ? byte_1024 : _GEN_4068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4545 = mask_4[1] ? byte_1025 : _GEN_4069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4546 = mask_4[2] ? byte_1026 : _GEN_4070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4547 = mask_4[3] ? byte_1027 : _GEN_4071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4548 = _GEN_8722 == 8'h37 ? _GEN_4544 : _GEN_4068; // @[executor.scala 473:84]
  wire [7:0] _GEN_4549 = _GEN_8722 == 8'h37 ? _GEN_4545 : _GEN_4069; // @[executor.scala 473:84]
  wire [7:0] _GEN_4550 = _GEN_8722 == 8'h37 ? _GEN_4546 : _GEN_4070; // @[executor.scala 473:84]
  wire [7:0] _GEN_4551 = _GEN_8722 == 8'h37 ? _GEN_4547 : _GEN_4071; // @[executor.scala 473:84]
  wire [7:0] _GEN_4552 = mask_4[0] ? byte_1024 : _GEN_4072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4553 = mask_4[1] ? byte_1025 : _GEN_4073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4554 = mask_4[2] ? byte_1026 : _GEN_4074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4555 = mask_4[3] ? byte_1027 : _GEN_4075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4556 = _GEN_8722 == 8'h38 ? _GEN_4552 : _GEN_4072; // @[executor.scala 473:84]
  wire [7:0] _GEN_4557 = _GEN_8722 == 8'h38 ? _GEN_4553 : _GEN_4073; // @[executor.scala 473:84]
  wire [7:0] _GEN_4558 = _GEN_8722 == 8'h38 ? _GEN_4554 : _GEN_4074; // @[executor.scala 473:84]
  wire [7:0] _GEN_4559 = _GEN_8722 == 8'h38 ? _GEN_4555 : _GEN_4075; // @[executor.scala 473:84]
  wire [7:0] _GEN_4560 = mask_4[0] ? byte_1024 : _GEN_4076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4561 = mask_4[1] ? byte_1025 : _GEN_4077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4562 = mask_4[2] ? byte_1026 : _GEN_4078; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4563 = mask_4[3] ? byte_1027 : _GEN_4079; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4564 = _GEN_8722 == 8'h39 ? _GEN_4560 : _GEN_4076; // @[executor.scala 473:84]
  wire [7:0] _GEN_4565 = _GEN_8722 == 8'h39 ? _GEN_4561 : _GEN_4077; // @[executor.scala 473:84]
  wire [7:0] _GEN_4566 = _GEN_8722 == 8'h39 ? _GEN_4562 : _GEN_4078; // @[executor.scala 473:84]
  wire [7:0] _GEN_4567 = _GEN_8722 == 8'h39 ? _GEN_4563 : _GEN_4079; // @[executor.scala 473:84]
  wire [7:0] _GEN_4568 = mask_4[0] ? byte_1024 : _GEN_4080; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4569 = mask_4[1] ? byte_1025 : _GEN_4081; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4570 = mask_4[2] ? byte_1026 : _GEN_4082; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4571 = mask_4[3] ? byte_1027 : _GEN_4083; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4572 = _GEN_8722 == 8'h3a ? _GEN_4568 : _GEN_4080; // @[executor.scala 473:84]
  wire [7:0] _GEN_4573 = _GEN_8722 == 8'h3a ? _GEN_4569 : _GEN_4081; // @[executor.scala 473:84]
  wire [7:0] _GEN_4574 = _GEN_8722 == 8'h3a ? _GEN_4570 : _GEN_4082; // @[executor.scala 473:84]
  wire [7:0] _GEN_4575 = _GEN_8722 == 8'h3a ? _GEN_4571 : _GEN_4083; // @[executor.scala 473:84]
  wire [7:0] _GEN_4576 = mask_4[0] ? byte_1024 : _GEN_4084; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4577 = mask_4[1] ? byte_1025 : _GEN_4085; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4578 = mask_4[2] ? byte_1026 : _GEN_4086; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4579 = mask_4[3] ? byte_1027 : _GEN_4087; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4580 = _GEN_8722 == 8'h3b ? _GEN_4576 : _GEN_4084; // @[executor.scala 473:84]
  wire [7:0] _GEN_4581 = _GEN_8722 == 8'h3b ? _GEN_4577 : _GEN_4085; // @[executor.scala 473:84]
  wire [7:0] _GEN_4582 = _GEN_8722 == 8'h3b ? _GEN_4578 : _GEN_4086; // @[executor.scala 473:84]
  wire [7:0] _GEN_4583 = _GEN_8722 == 8'h3b ? _GEN_4579 : _GEN_4087; // @[executor.scala 473:84]
  wire [7:0] _GEN_4584 = mask_4[0] ? byte_1024 : _GEN_4088; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4585 = mask_4[1] ? byte_1025 : _GEN_4089; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4586 = mask_4[2] ? byte_1026 : _GEN_4090; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4587 = mask_4[3] ? byte_1027 : _GEN_4091; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4588 = _GEN_8722 == 8'h3c ? _GEN_4584 : _GEN_4088; // @[executor.scala 473:84]
  wire [7:0] _GEN_4589 = _GEN_8722 == 8'h3c ? _GEN_4585 : _GEN_4089; // @[executor.scala 473:84]
  wire [7:0] _GEN_4590 = _GEN_8722 == 8'h3c ? _GEN_4586 : _GEN_4090; // @[executor.scala 473:84]
  wire [7:0] _GEN_4591 = _GEN_8722 == 8'h3c ? _GEN_4587 : _GEN_4091; // @[executor.scala 473:84]
  wire [7:0] _GEN_4592 = mask_4[0] ? byte_1024 : _GEN_4092; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4593 = mask_4[1] ? byte_1025 : _GEN_4093; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4594 = mask_4[2] ? byte_1026 : _GEN_4094; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4595 = mask_4[3] ? byte_1027 : _GEN_4095; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4596 = _GEN_8722 == 8'h3d ? _GEN_4592 : _GEN_4092; // @[executor.scala 473:84]
  wire [7:0] _GEN_4597 = _GEN_8722 == 8'h3d ? _GEN_4593 : _GEN_4093; // @[executor.scala 473:84]
  wire [7:0] _GEN_4598 = _GEN_8722 == 8'h3d ? _GEN_4594 : _GEN_4094; // @[executor.scala 473:84]
  wire [7:0] _GEN_4599 = _GEN_8722 == 8'h3d ? _GEN_4595 : _GEN_4095; // @[executor.scala 473:84]
  wire [7:0] _GEN_4600 = mask_4[0] ? byte_1024 : _GEN_4096; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4601 = mask_4[1] ? byte_1025 : _GEN_4097; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4602 = mask_4[2] ? byte_1026 : _GEN_4098; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4603 = mask_4[3] ? byte_1027 : _GEN_4099; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4604 = _GEN_8722 == 8'h3e ? _GEN_4600 : _GEN_4096; // @[executor.scala 473:84]
  wire [7:0] _GEN_4605 = _GEN_8722 == 8'h3e ? _GEN_4601 : _GEN_4097; // @[executor.scala 473:84]
  wire [7:0] _GEN_4606 = _GEN_8722 == 8'h3e ? _GEN_4602 : _GEN_4098; // @[executor.scala 473:84]
  wire [7:0] _GEN_4607 = _GEN_8722 == 8'h3e ? _GEN_4603 : _GEN_4099; // @[executor.scala 473:84]
  wire [7:0] _GEN_4608 = mask_4[0] ? byte_1024 : _GEN_4100; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4609 = mask_4[1] ? byte_1025 : _GEN_4101; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4610 = mask_4[2] ? byte_1026 : _GEN_4102; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4611 = mask_4[3] ? byte_1027 : _GEN_4103; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4612 = _GEN_8722 == 8'h3f ? _GEN_4608 : _GEN_4100; // @[executor.scala 473:84]
  wire [7:0] _GEN_4613 = _GEN_8722 == 8'h3f ? _GEN_4609 : _GEN_4101; // @[executor.scala 473:84]
  wire [7:0] _GEN_4614 = _GEN_8722 == 8'h3f ? _GEN_4610 : _GEN_4102; // @[executor.scala 473:84]
  wire [7:0] _GEN_4615 = _GEN_8722 == 8'h3f ? _GEN_4611 : _GEN_4103; // @[executor.scala 473:84]
  wire [7:0] _GEN_4616 = opcode_4 != 4'h0 ? _GEN_4108 : _GEN_3848; // @[executor.scala 470:55]
  wire [7:0] _GEN_4617 = opcode_4 != 4'h0 ? _GEN_4109 : _GEN_3849; // @[executor.scala 470:55]
  wire [7:0] _GEN_4618 = opcode_4 != 4'h0 ? _GEN_4110 : _GEN_3850; // @[executor.scala 470:55]
  wire [7:0] _GEN_4619 = opcode_4 != 4'h0 ? _GEN_4111 : _GEN_3851; // @[executor.scala 470:55]
  wire [7:0] _GEN_4620 = opcode_4 != 4'h0 ? _GEN_4116 : _GEN_3852; // @[executor.scala 470:55]
  wire [7:0] _GEN_4621 = opcode_4 != 4'h0 ? _GEN_4117 : _GEN_3853; // @[executor.scala 470:55]
  wire [7:0] _GEN_4622 = opcode_4 != 4'h0 ? _GEN_4118 : _GEN_3854; // @[executor.scala 470:55]
  wire [7:0] _GEN_4623 = opcode_4 != 4'h0 ? _GEN_4119 : _GEN_3855; // @[executor.scala 470:55]
  wire [7:0] _GEN_4624 = opcode_4 != 4'h0 ? _GEN_4124 : _GEN_3856; // @[executor.scala 470:55]
  wire [7:0] _GEN_4625 = opcode_4 != 4'h0 ? _GEN_4125 : _GEN_3857; // @[executor.scala 470:55]
  wire [7:0] _GEN_4626 = opcode_4 != 4'h0 ? _GEN_4126 : _GEN_3858; // @[executor.scala 470:55]
  wire [7:0] _GEN_4627 = opcode_4 != 4'h0 ? _GEN_4127 : _GEN_3859; // @[executor.scala 470:55]
  wire [7:0] _GEN_4628 = opcode_4 != 4'h0 ? _GEN_4132 : _GEN_3860; // @[executor.scala 470:55]
  wire [7:0] _GEN_4629 = opcode_4 != 4'h0 ? _GEN_4133 : _GEN_3861; // @[executor.scala 470:55]
  wire [7:0] _GEN_4630 = opcode_4 != 4'h0 ? _GEN_4134 : _GEN_3862; // @[executor.scala 470:55]
  wire [7:0] _GEN_4631 = opcode_4 != 4'h0 ? _GEN_4135 : _GEN_3863; // @[executor.scala 470:55]
  wire [7:0] _GEN_4632 = opcode_4 != 4'h0 ? _GEN_4140 : _GEN_3864; // @[executor.scala 470:55]
  wire [7:0] _GEN_4633 = opcode_4 != 4'h0 ? _GEN_4141 : _GEN_3865; // @[executor.scala 470:55]
  wire [7:0] _GEN_4634 = opcode_4 != 4'h0 ? _GEN_4142 : _GEN_3866; // @[executor.scala 470:55]
  wire [7:0] _GEN_4635 = opcode_4 != 4'h0 ? _GEN_4143 : _GEN_3867; // @[executor.scala 470:55]
  wire [7:0] _GEN_4636 = opcode_4 != 4'h0 ? _GEN_4148 : _GEN_3868; // @[executor.scala 470:55]
  wire [7:0] _GEN_4637 = opcode_4 != 4'h0 ? _GEN_4149 : _GEN_3869; // @[executor.scala 470:55]
  wire [7:0] _GEN_4638 = opcode_4 != 4'h0 ? _GEN_4150 : _GEN_3870; // @[executor.scala 470:55]
  wire [7:0] _GEN_4639 = opcode_4 != 4'h0 ? _GEN_4151 : _GEN_3871; // @[executor.scala 470:55]
  wire [7:0] _GEN_4640 = opcode_4 != 4'h0 ? _GEN_4156 : _GEN_3872; // @[executor.scala 470:55]
  wire [7:0] _GEN_4641 = opcode_4 != 4'h0 ? _GEN_4157 : _GEN_3873; // @[executor.scala 470:55]
  wire [7:0] _GEN_4642 = opcode_4 != 4'h0 ? _GEN_4158 : _GEN_3874; // @[executor.scala 470:55]
  wire [7:0] _GEN_4643 = opcode_4 != 4'h0 ? _GEN_4159 : _GEN_3875; // @[executor.scala 470:55]
  wire [7:0] _GEN_4644 = opcode_4 != 4'h0 ? _GEN_4164 : _GEN_3876; // @[executor.scala 470:55]
  wire [7:0] _GEN_4645 = opcode_4 != 4'h0 ? _GEN_4165 : _GEN_3877; // @[executor.scala 470:55]
  wire [7:0] _GEN_4646 = opcode_4 != 4'h0 ? _GEN_4166 : _GEN_3878; // @[executor.scala 470:55]
  wire [7:0] _GEN_4647 = opcode_4 != 4'h0 ? _GEN_4167 : _GEN_3879; // @[executor.scala 470:55]
  wire [7:0] _GEN_4648 = opcode_4 != 4'h0 ? _GEN_4172 : _GEN_3880; // @[executor.scala 470:55]
  wire [7:0] _GEN_4649 = opcode_4 != 4'h0 ? _GEN_4173 : _GEN_3881; // @[executor.scala 470:55]
  wire [7:0] _GEN_4650 = opcode_4 != 4'h0 ? _GEN_4174 : _GEN_3882; // @[executor.scala 470:55]
  wire [7:0] _GEN_4651 = opcode_4 != 4'h0 ? _GEN_4175 : _GEN_3883; // @[executor.scala 470:55]
  wire [7:0] _GEN_4652 = opcode_4 != 4'h0 ? _GEN_4180 : _GEN_3884; // @[executor.scala 470:55]
  wire [7:0] _GEN_4653 = opcode_4 != 4'h0 ? _GEN_4181 : _GEN_3885; // @[executor.scala 470:55]
  wire [7:0] _GEN_4654 = opcode_4 != 4'h0 ? _GEN_4182 : _GEN_3886; // @[executor.scala 470:55]
  wire [7:0] _GEN_4655 = opcode_4 != 4'h0 ? _GEN_4183 : _GEN_3887; // @[executor.scala 470:55]
  wire [7:0] _GEN_4656 = opcode_4 != 4'h0 ? _GEN_4188 : _GEN_3888; // @[executor.scala 470:55]
  wire [7:0] _GEN_4657 = opcode_4 != 4'h0 ? _GEN_4189 : _GEN_3889; // @[executor.scala 470:55]
  wire [7:0] _GEN_4658 = opcode_4 != 4'h0 ? _GEN_4190 : _GEN_3890; // @[executor.scala 470:55]
  wire [7:0] _GEN_4659 = opcode_4 != 4'h0 ? _GEN_4191 : _GEN_3891; // @[executor.scala 470:55]
  wire [7:0] _GEN_4660 = opcode_4 != 4'h0 ? _GEN_4196 : _GEN_3892; // @[executor.scala 470:55]
  wire [7:0] _GEN_4661 = opcode_4 != 4'h0 ? _GEN_4197 : _GEN_3893; // @[executor.scala 470:55]
  wire [7:0] _GEN_4662 = opcode_4 != 4'h0 ? _GEN_4198 : _GEN_3894; // @[executor.scala 470:55]
  wire [7:0] _GEN_4663 = opcode_4 != 4'h0 ? _GEN_4199 : _GEN_3895; // @[executor.scala 470:55]
  wire [7:0] _GEN_4664 = opcode_4 != 4'h0 ? _GEN_4204 : _GEN_3896; // @[executor.scala 470:55]
  wire [7:0] _GEN_4665 = opcode_4 != 4'h0 ? _GEN_4205 : _GEN_3897; // @[executor.scala 470:55]
  wire [7:0] _GEN_4666 = opcode_4 != 4'h0 ? _GEN_4206 : _GEN_3898; // @[executor.scala 470:55]
  wire [7:0] _GEN_4667 = opcode_4 != 4'h0 ? _GEN_4207 : _GEN_3899; // @[executor.scala 470:55]
  wire [7:0] _GEN_4668 = opcode_4 != 4'h0 ? _GEN_4212 : _GEN_3900; // @[executor.scala 470:55]
  wire [7:0] _GEN_4669 = opcode_4 != 4'h0 ? _GEN_4213 : _GEN_3901; // @[executor.scala 470:55]
  wire [7:0] _GEN_4670 = opcode_4 != 4'h0 ? _GEN_4214 : _GEN_3902; // @[executor.scala 470:55]
  wire [7:0] _GEN_4671 = opcode_4 != 4'h0 ? _GEN_4215 : _GEN_3903; // @[executor.scala 470:55]
  wire [7:0] _GEN_4672 = opcode_4 != 4'h0 ? _GEN_4220 : _GEN_3904; // @[executor.scala 470:55]
  wire [7:0] _GEN_4673 = opcode_4 != 4'h0 ? _GEN_4221 : _GEN_3905; // @[executor.scala 470:55]
  wire [7:0] _GEN_4674 = opcode_4 != 4'h0 ? _GEN_4222 : _GEN_3906; // @[executor.scala 470:55]
  wire [7:0] _GEN_4675 = opcode_4 != 4'h0 ? _GEN_4223 : _GEN_3907; // @[executor.scala 470:55]
  wire [7:0] _GEN_4676 = opcode_4 != 4'h0 ? _GEN_4228 : _GEN_3908; // @[executor.scala 470:55]
  wire [7:0] _GEN_4677 = opcode_4 != 4'h0 ? _GEN_4229 : _GEN_3909; // @[executor.scala 470:55]
  wire [7:0] _GEN_4678 = opcode_4 != 4'h0 ? _GEN_4230 : _GEN_3910; // @[executor.scala 470:55]
  wire [7:0] _GEN_4679 = opcode_4 != 4'h0 ? _GEN_4231 : _GEN_3911; // @[executor.scala 470:55]
  wire [7:0] _GEN_4680 = opcode_4 != 4'h0 ? _GEN_4236 : _GEN_3912; // @[executor.scala 470:55]
  wire [7:0] _GEN_4681 = opcode_4 != 4'h0 ? _GEN_4237 : _GEN_3913; // @[executor.scala 470:55]
  wire [7:0] _GEN_4682 = opcode_4 != 4'h0 ? _GEN_4238 : _GEN_3914; // @[executor.scala 470:55]
  wire [7:0] _GEN_4683 = opcode_4 != 4'h0 ? _GEN_4239 : _GEN_3915; // @[executor.scala 470:55]
  wire [7:0] _GEN_4684 = opcode_4 != 4'h0 ? _GEN_4244 : _GEN_3916; // @[executor.scala 470:55]
  wire [7:0] _GEN_4685 = opcode_4 != 4'h0 ? _GEN_4245 : _GEN_3917; // @[executor.scala 470:55]
  wire [7:0] _GEN_4686 = opcode_4 != 4'h0 ? _GEN_4246 : _GEN_3918; // @[executor.scala 470:55]
  wire [7:0] _GEN_4687 = opcode_4 != 4'h0 ? _GEN_4247 : _GEN_3919; // @[executor.scala 470:55]
  wire [7:0] _GEN_4688 = opcode_4 != 4'h0 ? _GEN_4252 : _GEN_3920; // @[executor.scala 470:55]
  wire [7:0] _GEN_4689 = opcode_4 != 4'h0 ? _GEN_4253 : _GEN_3921; // @[executor.scala 470:55]
  wire [7:0] _GEN_4690 = opcode_4 != 4'h0 ? _GEN_4254 : _GEN_3922; // @[executor.scala 470:55]
  wire [7:0] _GEN_4691 = opcode_4 != 4'h0 ? _GEN_4255 : _GEN_3923; // @[executor.scala 470:55]
  wire [7:0] _GEN_4692 = opcode_4 != 4'h0 ? _GEN_4260 : _GEN_3924; // @[executor.scala 470:55]
  wire [7:0] _GEN_4693 = opcode_4 != 4'h0 ? _GEN_4261 : _GEN_3925; // @[executor.scala 470:55]
  wire [7:0] _GEN_4694 = opcode_4 != 4'h0 ? _GEN_4262 : _GEN_3926; // @[executor.scala 470:55]
  wire [7:0] _GEN_4695 = opcode_4 != 4'h0 ? _GEN_4263 : _GEN_3927; // @[executor.scala 470:55]
  wire [7:0] _GEN_4696 = opcode_4 != 4'h0 ? _GEN_4268 : _GEN_3928; // @[executor.scala 470:55]
  wire [7:0] _GEN_4697 = opcode_4 != 4'h0 ? _GEN_4269 : _GEN_3929; // @[executor.scala 470:55]
  wire [7:0] _GEN_4698 = opcode_4 != 4'h0 ? _GEN_4270 : _GEN_3930; // @[executor.scala 470:55]
  wire [7:0] _GEN_4699 = opcode_4 != 4'h0 ? _GEN_4271 : _GEN_3931; // @[executor.scala 470:55]
  wire [7:0] _GEN_4700 = opcode_4 != 4'h0 ? _GEN_4276 : _GEN_3932; // @[executor.scala 470:55]
  wire [7:0] _GEN_4701 = opcode_4 != 4'h0 ? _GEN_4277 : _GEN_3933; // @[executor.scala 470:55]
  wire [7:0] _GEN_4702 = opcode_4 != 4'h0 ? _GEN_4278 : _GEN_3934; // @[executor.scala 470:55]
  wire [7:0] _GEN_4703 = opcode_4 != 4'h0 ? _GEN_4279 : _GEN_3935; // @[executor.scala 470:55]
  wire [7:0] _GEN_4704 = opcode_4 != 4'h0 ? _GEN_4284 : _GEN_3936; // @[executor.scala 470:55]
  wire [7:0] _GEN_4705 = opcode_4 != 4'h0 ? _GEN_4285 : _GEN_3937; // @[executor.scala 470:55]
  wire [7:0] _GEN_4706 = opcode_4 != 4'h0 ? _GEN_4286 : _GEN_3938; // @[executor.scala 470:55]
  wire [7:0] _GEN_4707 = opcode_4 != 4'h0 ? _GEN_4287 : _GEN_3939; // @[executor.scala 470:55]
  wire [7:0] _GEN_4708 = opcode_4 != 4'h0 ? _GEN_4292 : _GEN_3940; // @[executor.scala 470:55]
  wire [7:0] _GEN_4709 = opcode_4 != 4'h0 ? _GEN_4293 : _GEN_3941; // @[executor.scala 470:55]
  wire [7:0] _GEN_4710 = opcode_4 != 4'h0 ? _GEN_4294 : _GEN_3942; // @[executor.scala 470:55]
  wire [7:0] _GEN_4711 = opcode_4 != 4'h0 ? _GEN_4295 : _GEN_3943; // @[executor.scala 470:55]
  wire [7:0] _GEN_4712 = opcode_4 != 4'h0 ? _GEN_4300 : _GEN_3944; // @[executor.scala 470:55]
  wire [7:0] _GEN_4713 = opcode_4 != 4'h0 ? _GEN_4301 : _GEN_3945; // @[executor.scala 470:55]
  wire [7:0] _GEN_4714 = opcode_4 != 4'h0 ? _GEN_4302 : _GEN_3946; // @[executor.scala 470:55]
  wire [7:0] _GEN_4715 = opcode_4 != 4'h0 ? _GEN_4303 : _GEN_3947; // @[executor.scala 470:55]
  wire [7:0] _GEN_4716 = opcode_4 != 4'h0 ? _GEN_4308 : _GEN_3948; // @[executor.scala 470:55]
  wire [7:0] _GEN_4717 = opcode_4 != 4'h0 ? _GEN_4309 : _GEN_3949; // @[executor.scala 470:55]
  wire [7:0] _GEN_4718 = opcode_4 != 4'h0 ? _GEN_4310 : _GEN_3950; // @[executor.scala 470:55]
  wire [7:0] _GEN_4719 = opcode_4 != 4'h0 ? _GEN_4311 : _GEN_3951; // @[executor.scala 470:55]
  wire [7:0] _GEN_4720 = opcode_4 != 4'h0 ? _GEN_4316 : _GEN_3952; // @[executor.scala 470:55]
  wire [7:0] _GEN_4721 = opcode_4 != 4'h0 ? _GEN_4317 : _GEN_3953; // @[executor.scala 470:55]
  wire [7:0] _GEN_4722 = opcode_4 != 4'h0 ? _GEN_4318 : _GEN_3954; // @[executor.scala 470:55]
  wire [7:0] _GEN_4723 = opcode_4 != 4'h0 ? _GEN_4319 : _GEN_3955; // @[executor.scala 470:55]
  wire [7:0] _GEN_4724 = opcode_4 != 4'h0 ? _GEN_4324 : _GEN_3956; // @[executor.scala 470:55]
  wire [7:0] _GEN_4725 = opcode_4 != 4'h0 ? _GEN_4325 : _GEN_3957; // @[executor.scala 470:55]
  wire [7:0] _GEN_4726 = opcode_4 != 4'h0 ? _GEN_4326 : _GEN_3958; // @[executor.scala 470:55]
  wire [7:0] _GEN_4727 = opcode_4 != 4'h0 ? _GEN_4327 : _GEN_3959; // @[executor.scala 470:55]
  wire [7:0] _GEN_4728 = opcode_4 != 4'h0 ? _GEN_4332 : _GEN_3960; // @[executor.scala 470:55]
  wire [7:0] _GEN_4729 = opcode_4 != 4'h0 ? _GEN_4333 : _GEN_3961; // @[executor.scala 470:55]
  wire [7:0] _GEN_4730 = opcode_4 != 4'h0 ? _GEN_4334 : _GEN_3962; // @[executor.scala 470:55]
  wire [7:0] _GEN_4731 = opcode_4 != 4'h0 ? _GEN_4335 : _GEN_3963; // @[executor.scala 470:55]
  wire [7:0] _GEN_4732 = opcode_4 != 4'h0 ? _GEN_4340 : _GEN_3964; // @[executor.scala 470:55]
  wire [7:0] _GEN_4733 = opcode_4 != 4'h0 ? _GEN_4341 : _GEN_3965; // @[executor.scala 470:55]
  wire [7:0] _GEN_4734 = opcode_4 != 4'h0 ? _GEN_4342 : _GEN_3966; // @[executor.scala 470:55]
  wire [7:0] _GEN_4735 = opcode_4 != 4'h0 ? _GEN_4343 : _GEN_3967; // @[executor.scala 470:55]
  wire [7:0] _GEN_4736 = opcode_4 != 4'h0 ? _GEN_4348 : _GEN_3968; // @[executor.scala 470:55]
  wire [7:0] _GEN_4737 = opcode_4 != 4'h0 ? _GEN_4349 : _GEN_3969; // @[executor.scala 470:55]
  wire [7:0] _GEN_4738 = opcode_4 != 4'h0 ? _GEN_4350 : _GEN_3970; // @[executor.scala 470:55]
  wire [7:0] _GEN_4739 = opcode_4 != 4'h0 ? _GEN_4351 : _GEN_3971; // @[executor.scala 470:55]
  wire [7:0] _GEN_4740 = opcode_4 != 4'h0 ? _GEN_4356 : _GEN_3972; // @[executor.scala 470:55]
  wire [7:0] _GEN_4741 = opcode_4 != 4'h0 ? _GEN_4357 : _GEN_3973; // @[executor.scala 470:55]
  wire [7:0] _GEN_4742 = opcode_4 != 4'h0 ? _GEN_4358 : _GEN_3974; // @[executor.scala 470:55]
  wire [7:0] _GEN_4743 = opcode_4 != 4'h0 ? _GEN_4359 : _GEN_3975; // @[executor.scala 470:55]
  wire [7:0] _GEN_4744 = opcode_4 != 4'h0 ? _GEN_4364 : _GEN_3976; // @[executor.scala 470:55]
  wire [7:0] _GEN_4745 = opcode_4 != 4'h0 ? _GEN_4365 : _GEN_3977; // @[executor.scala 470:55]
  wire [7:0] _GEN_4746 = opcode_4 != 4'h0 ? _GEN_4366 : _GEN_3978; // @[executor.scala 470:55]
  wire [7:0] _GEN_4747 = opcode_4 != 4'h0 ? _GEN_4367 : _GEN_3979; // @[executor.scala 470:55]
  wire [7:0] _GEN_4748 = opcode_4 != 4'h0 ? _GEN_4372 : _GEN_3980; // @[executor.scala 470:55]
  wire [7:0] _GEN_4749 = opcode_4 != 4'h0 ? _GEN_4373 : _GEN_3981; // @[executor.scala 470:55]
  wire [7:0] _GEN_4750 = opcode_4 != 4'h0 ? _GEN_4374 : _GEN_3982; // @[executor.scala 470:55]
  wire [7:0] _GEN_4751 = opcode_4 != 4'h0 ? _GEN_4375 : _GEN_3983; // @[executor.scala 470:55]
  wire [7:0] _GEN_4752 = opcode_4 != 4'h0 ? _GEN_4380 : _GEN_3984; // @[executor.scala 470:55]
  wire [7:0] _GEN_4753 = opcode_4 != 4'h0 ? _GEN_4381 : _GEN_3985; // @[executor.scala 470:55]
  wire [7:0] _GEN_4754 = opcode_4 != 4'h0 ? _GEN_4382 : _GEN_3986; // @[executor.scala 470:55]
  wire [7:0] _GEN_4755 = opcode_4 != 4'h0 ? _GEN_4383 : _GEN_3987; // @[executor.scala 470:55]
  wire [7:0] _GEN_4756 = opcode_4 != 4'h0 ? _GEN_4388 : _GEN_3988; // @[executor.scala 470:55]
  wire [7:0] _GEN_4757 = opcode_4 != 4'h0 ? _GEN_4389 : _GEN_3989; // @[executor.scala 470:55]
  wire [7:0] _GEN_4758 = opcode_4 != 4'h0 ? _GEN_4390 : _GEN_3990; // @[executor.scala 470:55]
  wire [7:0] _GEN_4759 = opcode_4 != 4'h0 ? _GEN_4391 : _GEN_3991; // @[executor.scala 470:55]
  wire [7:0] _GEN_4760 = opcode_4 != 4'h0 ? _GEN_4396 : _GEN_3992; // @[executor.scala 470:55]
  wire [7:0] _GEN_4761 = opcode_4 != 4'h0 ? _GEN_4397 : _GEN_3993; // @[executor.scala 470:55]
  wire [7:0] _GEN_4762 = opcode_4 != 4'h0 ? _GEN_4398 : _GEN_3994; // @[executor.scala 470:55]
  wire [7:0] _GEN_4763 = opcode_4 != 4'h0 ? _GEN_4399 : _GEN_3995; // @[executor.scala 470:55]
  wire [7:0] _GEN_4764 = opcode_4 != 4'h0 ? _GEN_4404 : _GEN_3996; // @[executor.scala 470:55]
  wire [7:0] _GEN_4765 = opcode_4 != 4'h0 ? _GEN_4405 : _GEN_3997; // @[executor.scala 470:55]
  wire [7:0] _GEN_4766 = opcode_4 != 4'h0 ? _GEN_4406 : _GEN_3998; // @[executor.scala 470:55]
  wire [7:0] _GEN_4767 = opcode_4 != 4'h0 ? _GEN_4407 : _GEN_3999; // @[executor.scala 470:55]
  wire [7:0] _GEN_4768 = opcode_4 != 4'h0 ? _GEN_4412 : _GEN_4000; // @[executor.scala 470:55]
  wire [7:0] _GEN_4769 = opcode_4 != 4'h0 ? _GEN_4413 : _GEN_4001; // @[executor.scala 470:55]
  wire [7:0] _GEN_4770 = opcode_4 != 4'h0 ? _GEN_4414 : _GEN_4002; // @[executor.scala 470:55]
  wire [7:0] _GEN_4771 = opcode_4 != 4'h0 ? _GEN_4415 : _GEN_4003; // @[executor.scala 470:55]
  wire [7:0] _GEN_4772 = opcode_4 != 4'h0 ? _GEN_4420 : _GEN_4004; // @[executor.scala 470:55]
  wire [7:0] _GEN_4773 = opcode_4 != 4'h0 ? _GEN_4421 : _GEN_4005; // @[executor.scala 470:55]
  wire [7:0] _GEN_4774 = opcode_4 != 4'h0 ? _GEN_4422 : _GEN_4006; // @[executor.scala 470:55]
  wire [7:0] _GEN_4775 = opcode_4 != 4'h0 ? _GEN_4423 : _GEN_4007; // @[executor.scala 470:55]
  wire [7:0] _GEN_4776 = opcode_4 != 4'h0 ? _GEN_4428 : _GEN_4008; // @[executor.scala 470:55]
  wire [7:0] _GEN_4777 = opcode_4 != 4'h0 ? _GEN_4429 : _GEN_4009; // @[executor.scala 470:55]
  wire [7:0] _GEN_4778 = opcode_4 != 4'h0 ? _GEN_4430 : _GEN_4010; // @[executor.scala 470:55]
  wire [7:0] _GEN_4779 = opcode_4 != 4'h0 ? _GEN_4431 : _GEN_4011; // @[executor.scala 470:55]
  wire [7:0] _GEN_4780 = opcode_4 != 4'h0 ? _GEN_4436 : _GEN_4012; // @[executor.scala 470:55]
  wire [7:0] _GEN_4781 = opcode_4 != 4'h0 ? _GEN_4437 : _GEN_4013; // @[executor.scala 470:55]
  wire [7:0] _GEN_4782 = opcode_4 != 4'h0 ? _GEN_4438 : _GEN_4014; // @[executor.scala 470:55]
  wire [7:0] _GEN_4783 = opcode_4 != 4'h0 ? _GEN_4439 : _GEN_4015; // @[executor.scala 470:55]
  wire [7:0] _GEN_4784 = opcode_4 != 4'h0 ? _GEN_4444 : _GEN_4016; // @[executor.scala 470:55]
  wire [7:0] _GEN_4785 = opcode_4 != 4'h0 ? _GEN_4445 : _GEN_4017; // @[executor.scala 470:55]
  wire [7:0] _GEN_4786 = opcode_4 != 4'h0 ? _GEN_4446 : _GEN_4018; // @[executor.scala 470:55]
  wire [7:0] _GEN_4787 = opcode_4 != 4'h0 ? _GEN_4447 : _GEN_4019; // @[executor.scala 470:55]
  wire [7:0] _GEN_4788 = opcode_4 != 4'h0 ? _GEN_4452 : _GEN_4020; // @[executor.scala 470:55]
  wire [7:0] _GEN_4789 = opcode_4 != 4'h0 ? _GEN_4453 : _GEN_4021; // @[executor.scala 470:55]
  wire [7:0] _GEN_4790 = opcode_4 != 4'h0 ? _GEN_4454 : _GEN_4022; // @[executor.scala 470:55]
  wire [7:0] _GEN_4791 = opcode_4 != 4'h0 ? _GEN_4455 : _GEN_4023; // @[executor.scala 470:55]
  wire [7:0] _GEN_4792 = opcode_4 != 4'h0 ? _GEN_4460 : _GEN_4024; // @[executor.scala 470:55]
  wire [7:0] _GEN_4793 = opcode_4 != 4'h0 ? _GEN_4461 : _GEN_4025; // @[executor.scala 470:55]
  wire [7:0] _GEN_4794 = opcode_4 != 4'h0 ? _GEN_4462 : _GEN_4026; // @[executor.scala 470:55]
  wire [7:0] _GEN_4795 = opcode_4 != 4'h0 ? _GEN_4463 : _GEN_4027; // @[executor.scala 470:55]
  wire [7:0] _GEN_4796 = opcode_4 != 4'h0 ? _GEN_4468 : _GEN_4028; // @[executor.scala 470:55]
  wire [7:0] _GEN_4797 = opcode_4 != 4'h0 ? _GEN_4469 : _GEN_4029; // @[executor.scala 470:55]
  wire [7:0] _GEN_4798 = opcode_4 != 4'h0 ? _GEN_4470 : _GEN_4030; // @[executor.scala 470:55]
  wire [7:0] _GEN_4799 = opcode_4 != 4'h0 ? _GEN_4471 : _GEN_4031; // @[executor.scala 470:55]
  wire [7:0] _GEN_4800 = opcode_4 != 4'h0 ? _GEN_4476 : _GEN_4032; // @[executor.scala 470:55]
  wire [7:0] _GEN_4801 = opcode_4 != 4'h0 ? _GEN_4477 : _GEN_4033; // @[executor.scala 470:55]
  wire [7:0] _GEN_4802 = opcode_4 != 4'h0 ? _GEN_4478 : _GEN_4034; // @[executor.scala 470:55]
  wire [7:0] _GEN_4803 = opcode_4 != 4'h0 ? _GEN_4479 : _GEN_4035; // @[executor.scala 470:55]
  wire [7:0] _GEN_4804 = opcode_4 != 4'h0 ? _GEN_4484 : _GEN_4036; // @[executor.scala 470:55]
  wire [7:0] _GEN_4805 = opcode_4 != 4'h0 ? _GEN_4485 : _GEN_4037; // @[executor.scala 470:55]
  wire [7:0] _GEN_4806 = opcode_4 != 4'h0 ? _GEN_4486 : _GEN_4038; // @[executor.scala 470:55]
  wire [7:0] _GEN_4807 = opcode_4 != 4'h0 ? _GEN_4487 : _GEN_4039; // @[executor.scala 470:55]
  wire [7:0] _GEN_4808 = opcode_4 != 4'h0 ? _GEN_4492 : _GEN_4040; // @[executor.scala 470:55]
  wire [7:0] _GEN_4809 = opcode_4 != 4'h0 ? _GEN_4493 : _GEN_4041; // @[executor.scala 470:55]
  wire [7:0] _GEN_4810 = opcode_4 != 4'h0 ? _GEN_4494 : _GEN_4042; // @[executor.scala 470:55]
  wire [7:0] _GEN_4811 = opcode_4 != 4'h0 ? _GEN_4495 : _GEN_4043; // @[executor.scala 470:55]
  wire [7:0] _GEN_4812 = opcode_4 != 4'h0 ? _GEN_4500 : _GEN_4044; // @[executor.scala 470:55]
  wire [7:0] _GEN_4813 = opcode_4 != 4'h0 ? _GEN_4501 : _GEN_4045; // @[executor.scala 470:55]
  wire [7:0] _GEN_4814 = opcode_4 != 4'h0 ? _GEN_4502 : _GEN_4046; // @[executor.scala 470:55]
  wire [7:0] _GEN_4815 = opcode_4 != 4'h0 ? _GEN_4503 : _GEN_4047; // @[executor.scala 470:55]
  wire [7:0] _GEN_4816 = opcode_4 != 4'h0 ? _GEN_4508 : _GEN_4048; // @[executor.scala 470:55]
  wire [7:0] _GEN_4817 = opcode_4 != 4'h0 ? _GEN_4509 : _GEN_4049; // @[executor.scala 470:55]
  wire [7:0] _GEN_4818 = opcode_4 != 4'h0 ? _GEN_4510 : _GEN_4050; // @[executor.scala 470:55]
  wire [7:0] _GEN_4819 = opcode_4 != 4'h0 ? _GEN_4511 : _GEN_4051; // @[executor.scala 470:55]
  wire [7:0] _GEN_4820 = opcode_4 != 4'h0 ? _GEN_4516 : _GEN_4052; // @[executor.scala 470:55]
  wire [7:0] _GEN_4821 = opcode_4 != 4'h0 ? _GEN_4517 : _GEN_4053; // @[executor.scala 470:55]
  wire [7:0] _GEN_4822 = opcode_4 != 4'h0 ? _GEN_4518 : _GEN_4054; // @[executor.scala 470:55]
  wire [7:0] _GEN_4823 = opcode_4 != 4'h0 ? _GEN_4519 : _GEN_4055; // @[executor.scala 470:55]
  wire [7:0] _GEN_4824 = opcode_4 != 4'h0 ? _GEN_4524 : _GEN_4056; // @[executor.scala 470:55]
  wire [7:0] _GEN_4825 = opcode_4 != 4'h0 ? _GEN_4525 : _GEN_4057; // @[executor.scala 470:55]
  wire [7:0] _GEN_4826 = opcode_4 != 4'h0 ? _GEN_4526 : _GEN_4058; // @[executor.scala 470:55]
  wire [7:0] _GEN_4827 = opcode_4 != 4'h0 ? _GEN_4527 : _GEN_4059; // @[executor.scala 470:55]
  wire [7:0] _GEN_4828 = opcode_4 != 4'h0 ? _GEN_4532 : _GEN_4060; // @[executor.scala 470:55]
  wire [7:0] _GEN_4829 = opcode_4 != 4'h0 ? _GEN_4533 : _GEN_4061; // @[executor.scala 470:55]
  wire [7:0] _GEN_4830 = opcode_4 != 4'h0 ? _GEN_4534 : _GEN_4062; // @[executor.scala 470:55]
  wire [7:0] _GEN_4831 = opcode_4 != 4'h0 ? _GEN_4535 : _GEN_4063; // @[executor.scala 470:55]
  wire [7:0] _GEN_4832 = opcode_4 != 4'h0 ? _GEN_4540 : _GEN_4064; // @[executor.scala 470:55]
  wire [7:0] _GEN_4833 = opcode_4 != 4'h0 ? _GEN_4541 : _GEN_4065; // @[executor.scala 470:55]
  wire [7:0] _GEN_4834 = opcode_4 != 4'h0 ? _GEN_4542 : _GEN_4066; // @[executor.scala 470:55]
  wire [7:0] _GEN_4835 = opcode_4 != 4'h0 ? _GEN_4543 : _GEN_4067; // @[executor.scala 470:55]
  wire [7:0] _GEN_4836 = opcode_4 != 4'h0 ? _GEN_4548 : _GEN_4068; // @[executor.scala 470:55]
  wire [7:0] _GEN_4837 = opcode_4 != 4'h0 ? _GEN_4549 : _GEN_4069; // @[executor.scala 470:55]
  wire [7:0] _GEN_4838 = opcode_4 != 4'h0 ? _GEN_4550 : _GEN_4070; // @[executor.scala 470:55]
  wire [7:0] _GEN_4839 = opcode_4 != 4'h0 ? _GEN_4551 : _GEN_4071; // @[executor.scala 470:55]
  wire [7:0] _GEN_4840 = opcode_4 != 4'h0 ? _GEN_4556 : _GEN_4072; // @[executor.scala 470:55]
  wire [7:0] _GEN_4841 = opcode_4 != 4'h0 ? _GEN_4557 : _GEN_4073; // @[executor.scala 470:55]
  wire [7:0] _GEN_4842 = opcode_4 != 4'h0 ? _GEN_4558 : _GEN_4074; // @[executor.scala 470:55]
  wire [7:0] _GEN_4843 = opcode_4 != 4'h0 ? _GEN_4559 : _GEN_4075; // @[executor.scala 470:55]
  wire [7:0] _GEN_4844 = opcode_4 != 4'h0 ? _GEN_4564 : _GEN_4076; // @[executor.scala 470:55]
  wire [7:0] _GEN_4845 = opcode_4 != 4'h0 ? _GEN_4565 : _GEN_4077; // @[executor.scala 470:55]
  wire [7:0] _GEN_4846 = opcode_4 != 4'h0 ? _GEN_4566 : _GEN_4078; // @[executor.scala 470:55]
  wire [7:0] _GEN_4847 = opcode_4 != 4'h0 ? _GEN_4567 : _GEN_4079; // @[executor.scala 470:55]
  wire [7:0] _GEN_4848 = opcode_4 != 4'h0 ? _GEN_4572 : _GEN_4080; // @[executor.scala 470:55]
  wire [7:0] _GEN_4849 = opcode_4 != 4'h0 ? _GEN_4573 : _GEN_4081; // @[executor.scala 470:55]
  wire [7:0] _GEN_4850 = opcode_4 != 4'h0 ? _GEN_4574 : _GEN_4082; // @[executor.scala 470:55]
  wire [7:0] _GEN_4851 = opcode_4 != 4'h0 ? _GEN_4575 : _GEN_4083; // @[executor.scala 470:55]
  wire [7:0] _GEN_4852 = opcode_4 != 4'h0 ? _GEN_4580 : _GEN_4084; // @[executor.scala 470:55]
  wire [7:0] _GEN_4853 = opcode_4 != 4'h0 ? _GEN_4581 : _GEN_4085; // @[executor.scala 470:55]
  wire [7:0] _GEN_4854 = opcode_4 != 4'h0 ? _GEN_4582 : _GEN_4086; // @[executor.scala 470:55]
  wire [7:0] _GEN_4855 = opcode_4 != 4'h0 ? _GEN_4583 : _GEN_4087; // @[executor.scala 470:55]
  wire [7:0] _GEN_4856 = opcode_4 != 4'h0 ? _GEN_4588 : _GEN_4088; // @[executor.scala 470:55]
  wire [7:0] _GEN_4857 = opcode_4 != 4'h0 ? _GEN_4589 : _GEN_4089; // @[executor.scala 470:55]
  wire [7:0] _GEN_4858 = opcode_4 != 4'h0 ? _GEN_4590 : _GEN_4090; // @[executor.scala 470:55]
  wire [7:0] _GEN_4859 = opcode_4 != 4'h0 ? _GEN_4591 : _GEN_4091; // @[executor.scala 470:55]
  wire [7:0] _GEN_4860 = opcode_4 != 4'h0 ? _GEN_4596 : _GEN_4092; // @[executor.scala 470:55]
  wire [7:0] _GEN_4861 = opcode_4 != 4'h0 ? _GEN_4597 : _GEN_4093; // @[executor.scala 470:55]
  wire [7:0] _GEN_4862 = opcode_4 != 4'h0 ? _GEN_4598 : _GEN_4094; // @[executor.scala 470:55]
  wire [7:0] _GEN_4863 = opcode_4 != 4'h0 ? _GEN_4599 : _GEN_4095; // @[executor.scala 470:55]
  wire [7:0] _GEN_4864 = opcode_4 != 4'h0 ? _GEN_4604 : _GEN_4096; // @[executor.scala 470:55]
  wire [7:0] _GEN_4865 = opcode_4 != 4'h0 ? _GEN_4605 : _GEN_4097; // @[executor.scala 470:55]
  wire [7:0] _GEN_4866 = opcode_4 != 4'h0 ? _GEN_4606 : _GEN_4098; // @[executor.scala 470:55]
  wire [7:0] _GEN_4867 = opcode_4 != 4'h0 ? _GEN_4607 : _GEN_4099; // @[executor.scala 470:55]
  wire [7:0] _GEN_4868 = opcode_4 != 4'h0 ? _GEN_4612 : _GEN_4100; // @[executor.scala 470:55]
  wire [7:0] _GEN_4869 = opcode_4 != 4'h0 ? _GEN_4613 : _GEN_4101; // @[executor.scala 470:55]
  wire [7:0] _GEN_4870 = opcode_4 != 4'h0 ? _GEN_4614 : _GEN_4102; // @[executor.scala 470:55]
  wire [7:0] _GEN_4871 = opcode_4 != 4'h0 ? _GEN_4615 : _GEN_4103; // @[executor.scala 470:55]
  wire [3:0] _GEN_4872 = opcode_4 == 4'hf ? parameter_2_4[13:10] : _GEN_3846; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_4873 = opcode_4 == 4'hf ? parameter_2_4[0] : _GEN_3847; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_4874 = opcode_4 == 4'hf ? _GEN_3848 : _GEN_4616; // @[executor.scala 466:52]
  wire [7:0] _GEN_4875 = opcode_4 == 4'hf ? _GEN_3849 : _GEN_4617; // @[executor.scala 466:52]
  wire [7:0] _GEN_4876 = opcode_4 == 4'hf ? _GEN_3850 : _GEN_4618; // @[executor.scala 466:52]
  wire [7:0] _GEN_4877 = opcode_4 == 4'hf ? _GEN_3851 : _GEN_4619; // @[executor.scala 466:52]
  wire [7:0] _GEN_4878 = opcode_4 == 4'hf ? _GEN_3852 : _GEN_4620; // @[executor.scala 466:52]
  wire [7:0] _GEN_4879 = opcode_4 == 4'hf ? _GEN_3853 : _GEN_4621; // @[executor.scala 466:52]
  wire [7:0] _GEN_4880 = opcode_4 == 4'hf ? _GEN_3854 : _GEN_4622; // @[executor.scala 466:52]
  wire [7:0] _GEN_4881 = opcode_4 == 4'hf ? _GEN_3855 : _GEN_4623; // @[executor.scala 466:52]
  wire [7:0] _GEN_4882 = opcode_4 == 4'hf ? _GEN_3856 : _GEN_4624; // @[executor.scala 466:52]
  wire [7:0] _GEN_4883 = opcode_4 == 4'hf ? _GEN_3857 : _GEN_4625; // @[executor.scala 466:52]
  wire [7:0] _GEN_4884 = opcode_4 == 4'hf ? _GEN_3858 : _GEN_4626; // @[executor.scala 466:52]
  wire [7:0] _GEN_4885 = opcode_4 == 4'hf ? _GEN_3859 : _GEN_4627; // @[executor.scala 466:52]
  wire [7:0] _GEN_4886 = opcode_4 == 4'hf ? _GEN_3860 : _GEN_4628; // @[executor.scala 466:52]
  wire [7:0] _GEN_4887 = opcode_4 == 4'hf ? _GEN_3861 : _GEN_4629; // @[executor.scala 466:52]
  wire [7:0] _GEN_4888 = opcode_4 == 4'hf ? _GEN_3862 : _GEN_4630; // @[executor.scala 466:52]
  wire [7:0] _GEN_4889 = opcode_4 == 4'hf ? _GEN_3863 : _GEN_4631; // @[executor.scala 466:52]
  wire [7:0] _GEN_4890 = opcode_4 == 4'hf ? _GEN_3864 : _GEN_4632; // @[executor.scala 466:52]
  wire [7:0] _GEN_4891 = opcode_4 == 4'hf ? _GEN_3865 : _GEN_4633; // @[executor.scala 466:52]
  wire [7:0] _GEN_4892 = opcode_4 == 4'hf ? _GEN_3866 : _GEN_4634; // @[executor.scala 466:52]
  wire [7:0] _GEN_4893 = opcode_4 == 4'hf ? _GEN_3867 : _GEN_4635; // @[executor.scala 466:52]
  wire [7:0] _GEN_4894 = opcode_4 == 4'hf ? _GEN_3868 : _GEN_4636; // @[executor.scala 466:52]
  wire [7:0] _GEN_4895 = opcode_4 == 4'hf ? _GEN_3869 : _GEN_4637; // @[executor.scala 466:52]
  wire [7:0] _GEN_4896 = opcode_4 == 4'hf ? _GEN_3870 : _GEN_4638; // @[executor.scala 466:52]
  wire [7:0] _GEN_4897 = opcode_4 == 4'hf ? _GEN_3871 : _GEN_4639; // @[executor.scala 466:52]
  wire [7:0] _GEN_4898 = opcode_4 == 4'hf ? _GEN_3872 : _GEN_4640; // @[executor.scala 466:52]
  wire [7:0] _GEN_4899 = opcode_4 == 4'hf ? _GEN_3873 : _GEN_4641; // @[executor.scala 466:52]
  wire [7:0] _GEN_4900 = opcode_4 == 4'hf ? _GEN_3874 : _GEN_4642; // @[executor.scala 466:52]
  wire [7:0] _GEN_4901 = opcode_4 == 4'hf ? _GEN_3875 : _GEN_4643; // @[executor.scala 466:52]
  wire [7:0] _GEN_4902 = opcode_4 == 4'hf ? _GEN_3876 : _GEN_4644; // @[executor.scala 466:52]
  wire [7:0] _GEN_4903 = opcode_4 == 4'hf ? _GEN_3877 : _GEN_4645; // @[executor.scala 466:52]
  wire [7:0] _GEN_4904 = opcode_4 == 4'hf ? _GEN_3878 : _GEN_4646; // @[executor.scala 466:52]
  wire [7:0] _GEN_4905 = opcode_4 == 4'hf ? _GEN_3879 : _GEN_4647; // @[executor.scala 466:52]
  wire [7:0] _GEN_4906 = opcode_4 == 4'hf ? _GEN_3880 : _GEN_4648; // @[executor.scala 466:52]
  wire [7:0] _GEN_4907 = opcode_4 == 4'hf ? _GEN_3881 : _GEN_4649; // @[executor.scala 466:52]
  wire [7:0] _GEN_4908 = opcode_4 == 4'hf ? _GEN_3882 : _GEN_4650; // @[executor.scala 466:52]
  wire [7:0] _GEN_4909 = opcode_4 == 4'hf ? _GEN_3883 : _GEN_4651; // @[executor.scala 466:52]
  wire [7:0] _GEN_4910 = opcode_4 == 4'hf ? _GEN_3884 : _GEN_4652; // @[executor.scala 466:52]
  wire [7:0] _GEN_4911 = opcode_4 == 4'hf ? _GEN_3885 : _GEN_4653; // @[executor.scala 466:52]
  wire [7:0] _GEN_4912 = opcode_4 == 4'hf ? _GEN_3886 : _GEN_4654; // @[executor.scala 466:52]
  wire [7:0] _GEN_4913 = opcode_4 == 4'hf ? _GEN_3887 : _GEN_4655; // @[executor.scala 466:52]
  wire [7:0] _GEN_4914 = opcode_4 == 4'hf ? _GEN_3888 : _GEN_4656; // @[executor.scala 466:52]
  wire [7:0] _GEN_4915 = opcode_4 == 4'hf ? _GEN_3889 : _GEN_4657; // @[executor.scala 466:52]
  wire [7:0] _GEN_4916 = opcode_4 == 4'hf ? _GEN_3890 : _GEN_4658; // @[executor.scala 466:52]
  wire [7:0] _GEN_4917 = opcode_4 == 4'hf ? _GEN_3891 : _GEN_4659; // @[executor.scala 466:52]
  wire [7:0] _GEN_4918 = opcode_4 == 4'hf ? _GEN_3892 : _GEN_4660; // @[executor.scala 466:52]
  wire [7:0] _GEN_4919 = opcode_4 == 4'hf ? _GEN_3893 : _GEN_4661; // @[executor.scala 466:52]
  wire [7:0] _GEN_4920 = opcode_4 == 4'hf ? _GEN_3894 : _GEN_4662; // @[executor.scala 466:52]
  wire [7:0] _GEN_4921 = opcode_4 == 4'hf ? _GEN_3895 : _GEN_4663; // @[executor.scala 466:52]
  wire [7:0] _GEN_4922 = opcode_4 == 4'hf ? _GEN_3896 : _GEN_4664; // @[executor.scala 466:52]
  wire [7:0] _GEN_4923 = opcode_4 == 4'hf ? _GEN_3897 : _GEN_4665; // @[executor.scala 466:52]
  wire [7:0] _GEN_4924 = opcode_4 == 4'hf ? _GEN_3898 : _GEN_4666; // @[executor.scala 466:52]
  wire [7:0] _GEN_4925 = opcode_4 == 4'hf ? _GEN_3899 : _GEN_4667; // @[executor.scala 466:52]
  wire [7:0] _GEN_4926 = opcode_4 == 4'hf ? _GEN_3900 : _GEN_4668; // @[executor.scala 466:52]
  wire [7:0] _GEN_4927 = opcode_4 == 4'hf ? _GEN_3901 : _GEN_4669; // @[executor.scala 466:52]
  wire [7:0] _GEN_4928 = opcode_4 == 4'hf ? _GEN_3902 : _GEN_4670; // @[executor.scala 466:52]
  wire [7:0] _GEN_4929 = opcode_4 == 4'hf ? _GEN_3903 : _GEN_4671; // @[executor.scala 466:52]
  wire [7:0] _GEN_4930 = opcode_4 == 4'hf ? _GEN_3904 : _GEN_4672; // @[executor.scala 466:52]
  wire [7:0] _GEN_4931 = opcode_4 == 4'hf ? _GEN_3905 : _GEN_4673; // @[executor.scala 466:52]
  wire [7:0] _GEN_4932 = opcode_4 == 4'hf ? _GEN_3906 : _GEN_4674; // @[executor.scala 466:52]
  wire [7:0] _GEN_4933 = opcode_4 == 4'hf ? _GEN_3907 : _GEN_4675; // @[executor.scala 466:52]
  wire [7:0] _GEN_4934 = opcode_4 == 4'hf ? _GEN_3908 : _GEN_4676; // @[executor.scala 466:52]
  wire [7:0] _GEN_4935 = opcode_4 == 4'hf ? _GEN_3909 : _GEN_4677; // @[executor.scala 466:52]
  wire [7:0] _GEN_4936 = opcode_4 == 4'hf ? _GEN_3910 : _GEN_4678; // @[executor.scala 466:52]
  wire [7:0] _GEN_4937 = opcode_4 == 4'hf ? _GEN_3911 : _GEN_4679; // @[executor.scala 466:52]
  wire [7:0] _GEN_4938 = opcode_4 == 4'hf ? _GEN_3912 : _GEN_4680; // @[executor.scala 466:52]
  wire [7:0] _GEN_4939 = opcode_4 == 4'hf ? _GEN_3913 : _GEN_4681; // @[executor.scala 466:52]
  wire [7:0] _GEN_4940 = opcode_4 == 4'hf ? _GEN_3914 : _GEN_4682; // @[executor.scala 466:52]
  wire [7:0] _GEN_4941 = opcode_4 == 4'hf ? _GEN_3915 : _GEN_4683; // @[executor.scala 466:52]
  wire [7:0] _GEN_4942 = opcode_4 == 4'hf ? _GEN_3916 : _GEN_4684; // @[executor.scala 466:52]
  wire [7:0] _GEN_4943 = opcode_4 == 4'hf ? _GEN_3917 : _GEN_4685; // @[executor.scala 466:52]
  wire [7:0] _GEN_4944 = opcode_4 == 4'hf ? _GEN_3918 : _GEN_4686; // @[executor.scala 466:52]
  wire [7:0] _GEN_4945 = opcode_4 == 4'hf ? _GEN_3919 : _GEN_4687; // @[executor.scala 466:52]
  wire [7:0] _GEN_4946 = opcode_4 == 4'hf ? _GEN_3920 : _GEN_4688; // @[executor.scala 466:52]
  wire [7:0] _GEN_4947 = opcode_4 == 4'hf ? _GEN_3921 : _GEN_4689; // @[executor.scala 466:52]
  wire [7:0] _GEN_4948 = opcode_4 == 4'hf ? _GEN_3922 : _GEN_4690; // @[executor.scala 466:52]
  wire [7:0] _GEN_4949 = opcode_4 == 4'hf ? _GEN_3923 : _GEN_4691; // @[executor.scala 466:52]
  wire [7:0] _GEN_4950 = opcode_4 == 4'hf ? _GEN_3924 : _GEN_4692; // @[executor.scala 466:52]
  wire [7:0] _GEN_4951 = opcode_4 == 4'hf ? _GEN_3925 : _GEN_4693; // @[executor.scala 466:52]
  wire [7:0] _GEN_4952 = opcode_4 == 4'hf ? _GEN_3926 : _GEN_4694; // @[executor.scala 466:52]
  wire [7:0] _GEN_4953 = opcode_4 == 4'hf ? _GEN_3927 : _GEN_4695; // @[executor.scala 466:52]
  wire [7:0] _GEN_4954 = opcode_4 == 4'hf ? _GEN_3928 : _GEN_4696; // @[executor.scala 466:52]
  wire [7:0] _GEN_4955 = opcode_4 == 4'hf ? _GEN_3929 : _GEN_4697; // @[executor.scala 466:52]
  wire [7:0] _GEN_4956 = opcode_4 == 4'hf ? _GEN_3930 : _GEN_4698; // @[executor.scala 466:52]
  wire [7:0] _GEN_4957 = opcode_4 == 4'hf ? _GEN_3931 : _GEN_4699; // @[executor.scala 466:52]
  wire [7:0] _GEN_4958 = opcode_4 == 4'hf ? _GEN_3932 : _GEN_4700; // @[executor.scala 466:52]
  wire [7:0] _GEN_4959 = opcode_4 == 4'hf ? _GEN_3933 : _GEN_4701; // @[executor.scala 466:52]
  wire [7:0] _GEN_4960 = opcode_4 == 4'hf ? _GEN_3934 : _GEN_4702; // @[executor.scala 466:52]
  wire [7:0] _GEN_4961 = opcode_4 == 4'hf ? _GEN_3935 : _GEN_4703; // @[executor.scala 466:52]
  wire [7:0] _GEN_4962 = opcode_4 == 4'hf ? _GEN_3936 : _GEN_4704; // @[executor.scala 466:52]
  wire [7:0] _GEN_4963 = opcode_4 == 4'hf ? _GEN_3937 : _GEN_4705; // @[executor.scala 466:52]
  wire [7:0] _GEN_4964 = opcode_4 == 4'hf ? _GEN_3938 : _GEN_4706; // @[executor.scala 466:52]
  wire [7:0] _GEN_4965 = opcode_4 == 4'hf ? _GEN_3939 : _GEN_4707; // @[executor.scala 466:52]
  wire [7:0] _GEN_4966 = opcode_4 == 4'hf ? _GEN_3940 : _GEN_4708; // @[executor.scala 466:52]
  wire [7:0] _GEN_4967 = opcode_4 == 4'hf ? _GEN_3941 : _GEN_4709; // @[executor.scala 466:52]
  wire [7:0] _GEN_4968 = opcode_4 == 4'hf ? _GEN_3942 : _GEN_4710; // @[executor.scala 466:52]
  wire [7:0] _GEN_4969 = opcode_4 == 4'hf ? _GEN_3943 : _GEN_4711; // @[executor.scala 466:52]
  wire [7:0] _GEN_4970 = opcode_4 == 4'hf ? _GEN_3944 : _GEN_4712; // @[executor.scala 466:52]
  wire [7:0] _GEN_4971 = opcode_4 == 4'hf ? _GEN_3945 : _GEN_4713; // @[executor.scala 466:52]
  wire [7:0] _GEN_4972 = opcode_4 == 4'hf ? _GEN_3946 : _GEN_4714; // @[executor.scala 466:52]
  wire [7:0] _GEN_4973 = opcode_4 == 4'hf ? _GEN_3947 : _GEN_4715; // @[executor.scala 466:52]
  wire [7:0] _GEN_4974 = opcode_4 == 4'hf ? _GEN_3948 : _GEN_4716; // @[executor.scala 466:52]
  wire [7:0] _GEN_4975 = opcode_4 == 4'hf ? _GEN_3949 : _GEN_4717; // @[executor.scala 466:52]
  wire [7:0] _GEN_4976 = opcode_4 == 4'hf ? _GEN_3950 : _GEN_4718; // @[executor.scala 466:52]
  wire [7:0] _GEN_4977 = opcode_4 == 4'hf ? _GEN_3951 : _GEN_4719; // @[executor.scala 466:52]
  wire [7:0] _GEN_4978 = opcode_4 == 4'hf ? _GEN_3952 : _GEN_4720; // @[executor.scala 466:52]
  wire [7:0] _GEN_4979 = opcode_4 == 4'hf ? _GEN_3953 : _GEN_4721; // @[executor.scala 466:52]
  wire [7:0] _GEN_4980 = opcode_4 == 4'hf ? _GEN_3954 : _GEN_4722; // @[executor.scala 466:52]
  wire [7:0] _GEN_4981 = opcode_4 == 4'hf ? _GEN_3955 : _GEN_4723; // @[executor.scala 466:52]
  wire [7:0] _GEN_4982 = opcode_4 == 4'hf ? _GEN_3956 : _GEN_4724; // @[executor.scala 466:52]
  wire [7:0] _GEN_4983 = opcode_4 == 4'hf ? _GEN_3957 : _GEN_4725; // @[executor.scala 466:52]
  wire [7:0] _GEN_4984 = opcode_4 == 4'hf ? _GEN_3958 : _GEN_4726; // @[executor.scala 466:52]
  wire [7:0] _GEN_4985 = opcode_4 == 4'hf ? _GEN_3959 : _GEN_4727; // @[executor.scala 466:52]
  wire [7:0] _GEN_4986 = opcode_4 == 4'hf ? _GEN_3960 : _GEN_4728; // @[executor.scala 466:52]
  wire [7:0] _GEN_4987 = opcode_4 == 4'hf ? _GEN_3961 : _GEN_4729; // @[executor.scala 466:52]
  wire [7:0] _GEN_4988 = opcode_4 == 4'hf ? _GEN_3962 : _GEN_4730; // @[executor.scala 466:52]
  wire [7:0] _GEN_4989 = opcode_4 == 4'hf ? _GEN_3963 : _GEN_4731; // @[executor.scala 466:52]
  wire [7:0] _GEN_4990 = opcode_4 == 4'hf ? _GEN_3964 : _GEN_4732; // @[executor.scala 466:52]
  wire [7:0] _GEN_4991 = opcode_4 == 4'hf ? _GEN_3965 : _GEN_4733; // @[executor.scala 466:52]
  wire [7:0] _GEN_4992 = opcode_4 == 4'hf ? _GEN_3966 : _GEN_4734; // @[executor.scala 466:52]
  wire [7:0] _GEN_4993 = opcode_4 == 4'hf ? _GEN_3967 : _GEN_4735; // @[executor.scala 466:52]
  wire [7:0] _GEN_4994 = opcode_4 == 4'hf ? _GEN_3968 : _GEN_4736; // @[executor.scala 466:52]
  wire [7:0] _GEN_4995 = opcode_4 == 4'hf ? _GEN_3969 : _GEN_4737; // @[executor.scala 466:52]
  wire [7:0] _GEN_4996 = opcode_4 == 4'hf ? _GEN_3970 : _GEN_4738; // @[executor.scala 466:52]
  wire [7:0] _GEN_4997 = opcode_4 == 4'hf ? _GEN_3971 : _GEN_4739; // @[executor.scala 466:52]
  wire [7:0] _GEN_4998 = opcode_4 == 4'hf ? _GEN_3972 : _GEN_4740; // @[executor.scala 466:52]
  wire [7:0] _GEN_4999 = opcode_4 == 4'hf ? _GEN_3973 : _GEN_4741; // @[executor.scala 466:52]
  wire [7:0] _GEN_5000 = opcode_4 == 4'hf ? _GEN_3974 : _GEN_4742; // @[executor.scala 466:52]
  wire [7:0] _GEN_5001 = opcode_4 == 4'hf ? _GEN_3975 : _GEN_4743; // @[executor.scala 466:52]
  wire [7:0] _GEN_5002 = opcode_4 == 4'hf ? _GEN_3976 : _GEN_4744; // @[executor.scala 466:52]
  wire [7:0] _GEN_5003 = opcode_4 == 4'hf ? _GEN_3977 : _GEN_4745; // @[executor.scala 466:52]
  wire [7:0] _GEN_5004 = opcode_4 == 4'hf ? _GEN_3978 : _GEN_4746; // @[executor.scala 466:52]
  wire [7:0] _GEN_5005 = opcode_4 == 4'hf ? _GEN_3979 : _GEN_4747; // @[executor.scala 466:52]
  wire [7:0] _GEN_5006 = opcode_4 == 4'hf ? _GEN_3980 : _GEN_4748; // @[executor.scala 466:52]
  wire [7:0] _GEN_5007 = opcode_4 == 4'hf ? _GEN_3981 : _GEN_4749; // @[executor.scala 466:52]
  wire [7:0] _GEN_5008 = opcode_4 == 4'hf ? _GEN_3982 : _GEN_4750; // @[executor.scala 466:52]
  wire [7:0] _GEN_5009 = opcode_4 == 4'hf ? _GEN_3983 : _GEN_4751; // @[executor.scala 466:52]
  wire [7:0] _GEN_5010 = opcode_4 == 4'hf ? _GEN_3984 : _GEN_4752; // @[executor.scala 466:52]
  wire [7:0] _GEN_5011 = opcode_4 == 4'hf ? _GEN_3985 : _GEN_4753; // @[executor.scala 466:52]
  wire [7:0] _GEN_5012 = opcode_4 == 4'hf ? _GEN_3986 : _GEN_4754; // @[executor.scala 466:52]
  wire [7:0] _GEN_5013 = opcode_4 == 4'hf ? _GEN_3987 : _GEN_4755; // @[executor.scala 466:52]
  wire [7:0] _GEN_5014 = opcode_4 == 4'hf ? _GEN_3988 : _GEN_4756; // @[executor.scala 466:52]
  wire [7:0] _GEN_5015 = opcode_4 == 4'hf ? _GEN_3989 : _GEN_4757; // @[executor.scala 466:52]
  wire [7:0] _GEN_5016 = opcode_4 == 4'hf ? _GEN_3990 : _GEN_4758; // @[executor.scala 466:52]
  wire [7:0] _GEN_5017 = opcode_4 == 4'hf ? _GEN_3991 : _GEN_4759; // @[executor.scala 466:52]
  wire [7:0] _GEN_5018 = opcode_4 == 4'hf ? _GEN_3992 : _GEN_4760; // @[executor.scala 466:52]
  wire [7:0] _GEN_5019 = opcode_4 == 4'hf ? _GEN_3993 : _GEN_4761; // @[executor.scala 466:52]
  wire [7:0] _GEN_5020 = opcode_4 == 4'hf ? _GEN_3994 : _GEN_4762; // @[executor.scala 466:52]
  wire [7:0] _GEN_5021 = opcode_4 == 4'hf ? _GEN_3995 : _GEN_4763; // @[executor.scala 466:52]
  wire [7:0] _GEN_5022 = opcode_4 == 4'hf ? _GEN_3996 : _GEN_4764; // @[executor.scala 466:52]
  wire [7:0] _GEN_5023 = opcode_4 == 4'hf ? _GEN_3997 : _GEN_4765; // @[executor.scala 466:52]
  wire [7:0] _GEN_5024 = opcode_4 == 4'hf ? _GEN_3998 : _GEN_4766; // @[executor.scala 466:52]
  wire [7:0] _GEN_5025 = opcode_4 == 4'hf ? _GEN_3999 : _GEN_4767; // @[executor.scala 466:52]
  wire [7:0] _GEN_5026 = opcode_4 == 4'hf ? _GEN_4000 : _GEN_4768; // @[executor.scala 466:52]
  wire [7:0] _GEN_5027 = opcode_4 == 4'hf ? _GEN_4001 : _GEN_4769; // @[executor.scala 466:52]
  wire [7:0] _GEN_5028 = opcode_4 == 4'hf ? _GEN_4002 : _GEN_4770; // @[executor.scala 466:52]
  wire [7:0] _GEN_5029 = opcode_4 == 4'hf ? _GEN_4003 : _GEN_4771; // @[executor.scala 466:52]
  wire [7:0] _GEN_5030 = opcode_4 == 4'hf ? _GEN_4004 : _GEN_4772; // @[executor.scala 466:52]
  wire [7:0] _GEN_5031 = opcode_4 == 4'hf ? _GEN_4005 : _GEN_4773; // @[executor.scala 466:52]
  wire [7:0] _GEN_5032 = opcode_4 == 4'hf ? _GEN_4006 : _GEN_4774; // @[executor.scala 466:52]
  wire [7:0] _GEN_5033 = opcode_4 == 4'hf ? _GEN_4007 : _GEN_4775; // @[executor.scala 466:52]
  wire [7:0] _GEN_5034 = opcode_4 == 4'hf ? _GEN_4008 : _GEN_4776; // @[executor.scala 466:52]
  wire [7:0] _GEN_5035 = opcode_4 == 4'hf ? _GEN_4009 : _GEN_4777; // @[executor.scala 466:52]
  wire [7:0] _GEN_5036 = opcode_4 == 4'hf ? _GEN_4010 : _GEN_4778; // @[executor.scala 466:52]
  wire [7:0] _GEN_5037 = opcode_4 == 4'hf ? _GEN_4011 : _GEN_4779; // @[executor.scala 466:52]
  wire [7:0] _GEN_5038 = opcode_4 == 4'hf ? _GEN_4012 : _GEN_4780; // @[executor.scala 466:52]
  wire [7:0] _GEN_5039 = opcode_4 == 4'hf ? _GEN_4013 : _GEN_4781; // @[executor.scala 466:52]
  wire [7:0] _GEN_5040 = opcode_4 == 4'hf ? _GEN_4014 : _GEN_4782; // @[executor.scala 466:52]
  wire [7:0] _GEN_5041 = opcode_4 == 4'hf ? _GEN_4015 : _GEN_4783; // @[executor.scala 466:52]
  wire [7:0] _GEN_5042 = opcode_4 == 4'hf ? _GEN_4016 : _GEN_4784; // @[executor.scala 466:52]
  wire [7:0] _GEN_5043 = opcode_4 == 4'hf ? _GEN_4017 : _GEN_4785; // @[executor.scala 466:52]
  wire [7:0] _GEN_5044 = opcode_4 == 4'hf ? _GEN_4018 : _GEN_4786; // @[executor.scala 466:52]
  wire [7:0] _GEN_5045 = opcode_4 == 4'hf ? _GEN_4019 : _GEN_4787; // @[executor.scala 466:52]
  wire [7:0] _GEN_5046 = opcode_4 == 4'hf ? _GEN_4020 : _GEN_4788; // @[executor.scala 466:52]
  wire [7:0] _GEN_5047 = opcode_4 == 4'hf ? _GEN_4021 : _GEN_4789; // @[executor.scala 466:52]
  wire [7:0] _GEN_5048 = opcode_4 == 4'hf ? _GEN_4022 : _GEN_4790; // @[executor.scala 466:52]
  wire [7:0] _GEN_5049 = opcode_4 == 4'hf ? _GEN_4023 : _GEN_4791; // @[executor.scala 466:52]
  wire [7:0] _GEN_5050 = opcode_4 == 4'hf ? _GEN_4024 : _GEN_4792; // @[executor.scala 466:52]
  wire [7:0] _GEN_5051 = opcode_4 == 4'hf ? _GEN_4025 : _GEN_4793; // @[executor.scala 466:52]
  wire [7:0] _GEN_5052 = opcode_4 == 4'hf ? _GEN_4026 : _GEN_4794; // @[executor.scala 466:52]
  wire [7:0] _GEN_5053 = opcode_4 == 4'hf ? _GEN_4027 : _GEN_4795; // @[executor.scala 466:52]
  wire [7:0] _GEN_5054 = opcode_4 == 4'hf ? _GEN_4028 : _GEN_4796; // @[executor.scala 466:52]
  wire [7:0] _GEN_5055 = opcode_4 == 4'hf ? _GEN_4029 : _GEN_4797; // @[executor.scala 466:52]
  wire [7:0] _GEN_5056 = opcode_4 == 4'hf ? _GEN_4030 : _GEN_4798; // @[executor.scala 466:52]
  wire [7:0] _GEN_5057 = opcode_4 == 4'hf ? _GEN_4031 : _GEN_4799; // @[executor.scala 466:52]
  wire [7:0] _GEN_5058 = opcode_4 == 4'hf ? _GEN_4032 : _GEN_4800; // @[executor.scala 466:52]
  wire [7:0] _GEN_5059 = opcode_4 == 4'hf ? _GEN_4033 : _GEN_4801; // @[executor.scala 466:52]
  wire [7:0] _GEN_5060 = opcode_4 == 4'hf ? _GEN_4034 : _GEN_4802; // @[executor.scala 466:52]
  wire [7:0] _GEN_5061 = opcode_4 == 4'hf ? _GEN_4035 : _GEN_4803; // @[executor.scala 466:52]
  wire [7:0] _GEN_5062 = opcode_4 == 4'hf ? _GEN_4036 : _GEN_4804; // @[executor.scala 466:52]
  wire [7:0] _GEN_5063 = opcode_4 == 4'hf ? _GEN_4037 : _GEN_4805; // @[executor.scala 466:52]
  wire [7:0] _GEN_5064 = opcode_4 == 4'hf ? _GEN_4038 : _GEN_4806; // @[executor.scala 466:52]
  wire [7:0] _GEN_5065 = opcode_4 == 4'hf ? _GEN_4039 : _GEN_4807; // @[executor.scala 466:52]
  wire [7:0] _GEN_5066 = opcode_4 == 4'hf ? _GEN_4040 : _GEN_4808; // @[executor.scala 466:52]
  wire [7:0] _GEN_5067 = opcode_4 == 4'hf ? _GEN_4041 : _GEN_4809; // @[executor.scala 466:52]
  wire [7:0] _GEN_5068 = opcode_4 == 4'hf ? _GEN_4042 : _GEN_4810; // @[executor.scala 466:52]
  wire [7:0] _GEN_5069 = opcode_4 == 4'hf ? _GEN_4043 : _GEN_4811; // @[executor.scala 466:52]
  wire [7:0] _GEN_5070 = opcode_4 == 4'hf ? _GEN_4044 : _GEN_4812; // @[executor.scala 466:52]
  wire [7:0] _GEN_5071 = opcode_4 == 4'hf ? _GEN_4045 : _GEN_4813; // @[executor.scala 466:52]
  wire [7:0] _GEN_5072 = opcode_4 == 4'hf ? _GEN_4046 : _GEN_4814; // @[executor.scala 466:52]
  wire [7:0] _GEN_5073 = opcode_4 == 4'hf ? _GEN_4047 : _GEN_4815; // @[executor.scala 466:52]
  wire [7:0] _GEN_5074 = opcode_4 == 4'hf ? _GEN_4048 : _GEN_4816; // @[executor.scala 466:52]
  wire [7:0] _GEN_5075 = opcode_4 == 4'hf ? _GEN_4049 : _GEN_4817; // @[executor.scala 466:52]
  wire [7:0] _GEN_5076 = opcode_4 == 4'hf ? _GEN_4050 : _GEN_4818; // @[executor.scala 466:52]
  wire [7:0] _GEN_5077 = opcode_4 == 4'hf ? _GEN_4051 : _GEN_4819; // @[executor.scala 466:52]
  wire [7:0] _GEN_5078 = opcode_4 == 4'hf ? _GEN_4052 : _GEN_4820; // @[executor.scala 466:52]
  wire [7:0] _GEN_5079 = opcode_4 == 4'hf ? _GEN_4053 : _GEN_4821; // @[executor.scala 466:52]
  wire [7:0] _GEN_5080 = opcode_4 == 4'hf ? _GEN_4054 : _GEN_4822; // @[executor.scala 466:52]
  wire [7:0] _GEN_5081 = opcode_4 == 4'hf ? _GEN_4055 : _GEN_4823; // @[executor.scala 466:52]
  wire [7:0] _GEN_5082 = opcode_4 == 4'hf ? _GEN_4056 : _GEN_4824; // @[executor.scala 466:52]
  wire [7:0] _GEN_5083 = opcode_4 == 4'hf ? _GEN_4057 : _GEN_4825; // @[executor.scala 466:52]
  wire [7:0] _GEN_5084 = opcode_4 == 4'hf ? _GEN_4058 : _GEN_4826; // @[executor.scala 466:52]
  wire [7:0] _GEN_5085 = opcode_4 == 4'hf ? _GEN_4059 : _GEN_4827; // @[executor.scala 466:52]
  wire [7:0] _GEN_5086 = opcode_4 == 4'hf ? _GEN_4060 : _GEN_4828; // @[executor.scala 466:52]
  wire [7:0] _GEN_5087 = opcode_4 == 4'hf ? _GEN_4061 : _GEN_4829; // @[executor.scala 466:52]
  wire [7:0] _GEN_5088 = opcode_4 == 4'hf ? _GEN_4062 : _GEN_4830; // @[executor.scala 466:52]
  wire [7:0] _GEN_5089 = opcode_4 == 4'hf ? _GEN_4063 : _GEN_4831; // @[executor.scala 466:52]
  wire [7:0] _GEN_5090 = opcode_4 == 4'hf ? _GEN_4064 : _GEN_4832; // @[executor.scala 466:52]
  wire [7:0] _GEN_5091 = opcode_4 == 4'hf ? _GEN_4065 : _GEN_4833; // @[executor.scala 466:52]
  wire [7:0] _GEN_5092 = opcode_4 == 4'hf ? _GEN_4066 : _GEN_4834; // @[executor.scala 466:52]
  wire [7:0] _GEN_5093 = opcode_4 == 4'hf ? _GEN_4067 : _GEN_4835; // @[executor.scala 466:52]
  wire [7:0] _GEN_5094 = opcode_4 == 4'hf ? _GEN_4068 : _GEN_4836; // @[executor.scala 466:52]
  wire [7:0] _GEN_5095 = opcode_4 == 4'hf ? _GEN_4069 : _GEN_4837; // @[executor.scala 466:52]
  wire [7:0] _GEN_5096 = opcode_4 == 4'hf ? _GEN_4070 : _GEN_4838; // @[executor.scala 466:52]
  wire [7:0] _GEN_5097 = opcode_4 == 4'hf ? _GEN_4071 : _GEN_4839; // @[executor.scala 466:52]
  wire [7:0] _GEN_5098 = opcode_4 == 4'hf ? _GEN_4072 : _GEN_4840; // @[executor.scala 466:52]
  wire [7:0] _GEN_5099 = opcode_4 == 4'hf ? _GEN_4073 : _GEN_4841; // @[executor.scala 466:52]
  wire [7:0] _GEN_5100 = opcode_4 == 4'hf ? _GEN_4074 : _GEN_4842; // @[executor.scala 466:52]
  wire [7:0] _GEN_5101 = opcode_4 == 4'hf ? _GEN_4075 : _GEN_4843; // @[executor.scala 466:52]
  wire [7:0] _GEN_5102 = opcode_4 == 4'hf ? _GEN_4076 : _GEN_4844; // @[executor.scala 466:52]
  wire [7:0] _GEN_5103 = opcode_4 == 4'hf ? _GEN_4077 : _GEN_4845; // @[executor.scala 466:52]
  wire [7:0] _GEN_5104 = opcode_4 == 4'hf ? _GEN_4078 : _GEN_4846; // @[executor.scala 466:52]
  wire [7:0] _GEN_5105 = opcode_4 == 4'hf ? _GEN_4079 : _GEN_4847; // @[executor.scala 466:52]
  wire [7:0] _GEN_5106 = opcode_4 == 4'hf ? _GEN_4080 : _GEN_4848; // @[executor.scala 466:52]
  wire [7:0] _GEN_5107 = opcode_4 == 4'hf ? _GEN_4081 : _GEN_4849; // @[executor.scala 466:52]
  wire [7:0] _GEN_5108 = opcode_4 == 4'hf ? _GEN_4082 : _GEN_4850; // @[executor.scala 466:52]
  wire [7:0] _GEN_5109 = opcode_4 == 4'hf ? _GEN_4083 : _GEN_4851; // @[executor.scala 466:52]
  wire [7:0] _GEN_5110 = opcode_4 == 4'hf ? _GEN_4084 : _GEN_4852; // @[executor.scala 466:52]
  wire [7:0] _GEN_5111 = opcode_4 == 4'hf ? _GEN_4085 : _GEN_4853; // @[executor.scala 466:52]
  wire [7:0] _GEN_5112 = opcode_4 == 4'hf ? _GEN_4086 : _GEN_4854; // @[executor.scala 466:52]
  wire [7:0] _GEN_5113 = opcode_4 == 4'hf ? _GEN_4087 : _GEN_4855; // @[executor.scala 466:52]
  wire [7:0] _GEN_5114 = opcode_4 == 4'hf ? _GEN_4088 : _GEN_4856; // @[executor.scala 466:52]
  wire [7:0] _GEN_5115 = opcode_4 == 4'hf ? _GEN_4089 : _GEN_4857; // @[executor.scala 466:52]
  wire [7:0] _GEN_5116 = opcode_4 == 4'hf ? _GEN_4090 : _GEN_4858; // @[executor.scala 466:52]
  wire [7:0] _GEN_5117 = opcode_4 == 4'hf ? _GEN_4091 : _GEN_4859; // @[executor.scala 466:52]
  wire [7:0] _GEN_5118 = opcode_4 == 4'hf ? _GEN_4092 : _GEN_4860; // @[executor.scala 466:52]
  wire [7:0] _GEN_5119 = opcode_4 == 4'hf ? _GEN_4093 : _GEN_4861; // @[executor.scala 466:52]
  wire [7:0] _GEN_5120 = opcode_4 == 4'hf ? _GEN_4094 : _GEN_4862; // @[executor.scala 466:52]
  wire [7:0] _GEN_5121 = opcode_4 == 4'hf ? _GEN_4095 : _GEN_4863; // @[executor.scala 466:52]
  wire [7:0] _GEN_5122 = opcode_4 == 4'hf ? _GEN_4096 : _GEN_4864; // @[executor.scala 466:52]
  wire [7:0] _GEN_5123 = opcode_4 == 4'hf ? _GEN_4097 : _GEN_4865; // @[executor.scala 466:52]
  wire [7:0] _GEN_5124 = opcode_4 == 4'hf ? _GEN_4098 : _GEN_4866; // @[executor.scala 466:52]
  wire [7:0] _GEN_5125 = opcode_4 == 4'hf ? _GEN_4099 : _GEN_4867; // @[executor.scala 466:52]
  wire [7:0] _GEN_5126 = opcode_4 == 4'hf ? _GEN_4100 : _GEN_4868; // @[executor.scala 466:52]
  wire [7:0] _GEN_5127 = opcode_4 == 4'hf ? _GEN_4101 : _GEN_4869; // @[executor.scala 466:52]
  wire [7:0] _GEN_5128 = opcode_4 == 4'hf ? _GEN_4102 : _GEN_4870; // @[executor.scala 466:52]
  wire [7:0] _GEN_5129 = opcode_4 == 4'hf ? _GEN_4103 : _GEN_4871; // @[executor.scala 466:52]
  wire [3:0] opcode_5 = vliw_5[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_5 = vliw_5[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8786 = {{2'd0}, dst_offset_5}; // @[executor.scala 473:49]
  wire [7:0] byte_1280 = field_5[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_5130 = mask_5[0] ? byte_1280 : _GEN_4874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1281 = field_5[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_5131 = mask_5[1] ? byte_1281 : _GEN_4875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1282 = field_5[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_5132 = mask_5[2] ? byte_1282 : _GEN_4876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1283 = field_5[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_5133 = mask_5[3] ? byte_1283 : _GEN_4877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5134 = _GEN_8786 == 8'h0 ? _GEN_5130 : _GEN_4874; // @[executor.scala 473:84]
  wire [7:0] _GEN_5135 = _GEN_8786 == 8'h0 ? _GEN_5131 : _GEN_4875; // @[executor.scala 473:84]
  wire [7:0] _GEN_5136 = _GEN_8786 == 8'h0 ? _GEN_5132 : _GEN_4876; // @[executor.scala 473:84]
  wire [7:0] _GEN_5137 = _GEN_8786 == 8'h0 ? _GEN_5133 : _GEN_4877; // @[executor.scala 473:84]
  wire [7:0] _GEN_5138 = mask_5[0] ? byte_1280 : _GEN_4878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5139 = mask_5[1] ? byte_1281 : _GEN_4879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5140 = mask_5[2] ? byte_1282 : _GEN_4880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5141 = mask_5[3] ? byte_1283 : _GEN_4881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5142 = _GEN_8786 == 8'h1 ? _GEN_5138 : _GEN_4878; // @[executor.scala 473:84]
  wire [7:0] _GEN_5143 = _GEN_8786 == 8'h1 ? _GEN_5139 : _GEN_4879; // @[executor.scala 473:84]
  wire [7:0] _GEN_5144 = _GEN_8786 == 8'h1 ? _GEN_5140 : _GEN_4880; // @[executor.scala 473:84]
  wire [7:0] _GEN_5145 = _GEN_8786 == 8'h1 ? _GEN_5141 : _GEN_4881; // @[executor.scala 473:84]
  wire [7:0] _GEN_5146 = mask_5[0] ? byte_1280 : _GEN_4882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5147 = mask_5[1] ? byte_1281 : _GEN_4883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5148 = mask_5[2] ? byte_1282 : _GEN_4884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5149 = mask_5[3] ? byte_1283 : _GEN_4885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5150 = _GEN_8786 == 8'h2 ? _GEN_5146 : _GEN_4882; // @[executor.scala 473:84]
  wire [7:0] _GEN_5151 = _GEN_8786 == 8'h2 ? _GEN_5147 : _GEN_4883; // @[executor.scala 473:84]
  wire [7:0] _GEN_5152 = _GEN_8786 == 8'h2 ? _GEN_5148 : _GEN_4884; // @[executor.scala 473:84]
  wire [7:0] _GEN_5153 = _GEN_8786 == 8'h2 ? _GEN_5149 : _GEN_4885; // @[executor.scala 473:84]
  wire [7:0] _GEN_5154 = mask_5[0] ? byte_1280 : _GEN_4886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5155 = mask_5[1] ? byte_1281 : _GEN_4887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5156 = mask_5[2] ? byte_1282 : _GEN_4888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5157 = mask_5[3] ? byte_1283 : _GEN_4889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5158 = _GEN_8786 == 8'h3 ? _GEN_5154 : _GEN_4886; // @[executor.scala 473:84]
  wire [7:0] _GEN_5159 = _GEN_8786 == 8'h3 ? _GEN_5155 : _GEN_4887; // @[executor.scala 473:84]
  wire [7:0] _GEN_5160 = _GEN_8786 == 8'h3 ? _GEN_5156 : _GEN_4888; // @[executor.scala 473:84]
  wire [7:0] _GEN_5161 = _GEN_8786 == 8'h3 ? _GEN_5157 : _GEN_4889; // @[executor.scala 473:84]
  wire [7:0] _GEN_5162 = mask_5[0] ? byte_1280 : _GEN_4890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5163 = mask_5[1] ? byte_1281 : _GEN_4891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5164 = mask_5[2] ? byte_1282 : _GEN_4892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5165 = mask_5[3] ? byte_1283 : _GEN_4893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5166 = _GEN_8786 == 8'h4 ? _GEN_5162 : _GEN_4890; // @[executor.scala 473:84]
  wire [7:0] _GEN_5167 = _GEN_8786 == 8'h4 ? _GEN_5163 : _GEN_4891; // @[executor.scala 473:84]
  wire [7:0] _GEN_5168 = _GEN_8786 == 8'h4 ? _GEN_5164 : _GEN_4892; // @[executor.scala 473:84]
  wire [7:0] _GEN_5169 = _GEN_8786 == 8'h4 ? _GEN_5165 : _GEN_4893; // @[executor.scala 473:84]
  wire [7:0] _GEN_5170 = mask_5[0] ? byte_1280 : _GEN_4894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5171 = mask_5[1] ? byte_1281 : _GEN_4895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5172 = mask_5[2] ? byte_1282 : _GEN_4896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5173 = mask_5[3] ? byte_1283 : _GEN_4897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5174 = _GEN_8786 == 8'h5 ? _GEN_5170 : _GEN_4894; // @[executor.scala 473:84]
  wire [7:0] _GEN_5175 = _GEN_8786 == 8'h5 ? _GEN_5171 : _GEN_4895; // @[executor.scala 473:84]
  wire [7:0] _GEN_5176 = _GEN_8786 == 8'h5 ? _GEN_5172 : _GEN_4896; // @[executor.scala 473:84]
  wire [7:0] _GEN_5177 = _GEN_8786 == 8'h5 ? _GEN_5173 : _GEN_4897; // @[executor.scala 473:84]
  wire [7:0] _GEN_5178 = mask_5[0] ? byte_1280 : _GEN_4898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5179 = mask_5[1] ? byte_1281 : _GEN_4899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5180 = mask_5[2] ? byte_1282 : _GEN_4900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5181 = mask_5[3] ? byte_1283 : _GEN_4901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5182 = _GEN_8786 == 8'h6 ? _GEN_5178 : _GEN_4898; // @[executor.scala 473:84]
  wire [7:0] _GEN_5183 = _GEN_8786 == 8'h6 ? _GEN_5179 : _GEN_4899; // @[executor.scala 473:84]
  wire [7:0] _GEN_5184 = _GEN_8786 == 8'h6 ? _GEN_5180 : _GEN_4900; // @[executor.scala 473:84]
  wire [7:0] _GEN_5185 = _GEN_8786 == 8'h6 ? _GEN_5181 : _GEN_4901; // @[executor.scala 473:84]
  wire [7:0] _GEN_5186 = mask_5[0] ? byte_1280 : _GEN_4902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5187 = mask_5[1] ? byte_1281 : _GEN_4903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5188 = mask_5[2] ? byte_1282 : _GEN_4904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5189 = mask_5[3] ? byte_1283 : _GEN_4905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5190 = _GEN_8786 == 8'h7 ? _GEN_5186 : _GEN_4902; // @[executor.scala 473:84]
  wire [7:0] _GEN_5191 = _GEN_8786 == 8'h7 ? _GEN_5187 : _GEN_4903; // @[executor.scala 473:84]
  wire [7:0] _GEN_5192 = _GEN_8786 == 8'h7 ? _GEN_5188 : _GEN_4904; // @[executor.scala 473:84]
  wire [7:0] _GEN_5193 = _GEN_8786 == 8'h7 ? _GEN_5189 : _GEN_4905; // @[executor.scala 473:84]
  wire [7:0] _GEN_5194 = mask_5[0] ? byte_1280 : _GEN_4906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5195 = mask_5[1] ? byte_1281 : _GEN_4907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5196 = mask_5[2] ? byte_1282 : _GEN_4908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5197 = mask_5[3] ? byte_1283 : _GEN_4909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5198 = _GEN_8786 == 8'h8 ? _GEN_5194 : _GEN_4906; // @[executor.scala 473:84]
  wire [7:0] _GEN_5199 = _GEN_8786 == 8'h8 ? _GEN_5195 : _GEN_4907; // @[executor.scala 473:84]
  wire [7:0] _GEN_5200 = _GEN_8786 == 8'h8 ? _GEN_5196 : _GEN_4908; // @[executor.scala 473:84]
  wire [7:0] _GEN_5201 = _GEN_8786 == 8'h8 ? _GEN_5197 : _GEN_4909; // @[executor.scala 473:84]
  wire [7:0] _GEN_5202 = mask_5[0] ? byte_1280 : _GEN_4910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5203 = mask_5[1] ? byte_1281 : _GEN_4911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5204 = mask_5[2] ? byte_1282 : _GEN_4912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5205 = mask_5[3] ? byte_1283 : _GEN_4913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5206 = _GEN_8786 == 8'h9 ? _GEN_5202 : _GEN_4910; // @[executor.scala 473:84]
  wire [7:0] _GEN_5207 = _GEN_8786 == 8'h9 ? _GEN_5203 : _GEN_4911; // @[executor.scala 473:84]
  wire [7:0] _GEN_5208 = _GEN_8786 == 8'h9 ? _GEN_5204 : _GEN_4912; // @[executor.scala 473:84]
  wire [7:0] _GEN_5209 = _GEN_8786 == 8'h9 ? _GEN_5205 : _GEN_4913; // @[executor.scala 473:84]
  wire [7:0] _GEN_5210 = mask_5[0] ? byte_1280 : _GEN_4914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5211 = mask_5[1] ? byte_1281 : _GEN_4915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5212 = mask_5[2] ? byte_1282 : _GEN_4916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5213 = mask_5[3] ? byte_1283 : _GEN_4917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5214 = _GEN_8786 == 8'ha ? _GEN_5210 : _GEN_4914; // @[executor.scala 473:84]
  wire [7:0] _GEN_5215 = _GEN_8786 == 8'ha ? _GEN_5211 : _GEN_4915; // @[executor.scala 473:84]
  wire [7:0] _GEN_5216 = _GEN_8786 == 8'ha ? _GEN_5212 : _GEN_4916; // @[executor.scala 473:84]
  wire [7:0] _GEN_5217 = _GEN_8786 == 8'ha ? _GEN_5213 : _GEN_4917; // @[executor.scala 473:84]
  wire [7:0] _GEN_5218 = mask_5[0] ? byte_1280 : _GEN_4918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5219 = mask_5[1] ? byte_1281 : _GEN_4919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5220 = mask_5[2] ? byte_1282 : _GEN_4920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5221 = mask_5[3] ? byte_1283 : _GEN_4921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5222 = _GEN_8786 == 8'hb ? _GEN_5218 : _GEN_4918; // @[executor.scala 473:84]
  wire [7:0] _GEN_5223 = _GEN_8786 == 8'hb ? _GEN_5219 : _GEN_4919; // @[executor.scala 473:84]
  wire [7:0] _GEN_5224 = _GEN_8786 == 8'hb ? _GEN_5220 : _GEN_4920; // @[executor.scala 473:84]
  wire [7:0] _GEN_5225 = _GEN_8786 == 8'hb ? _GEN_5221 : _GEN_4921; // @[executor.scala 473:84]
  wire [7:0] _GEN_5226 = mask_5[0] ? byte_1280 : _GEN_4922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5227 = mask_5[1] ? byte_1281 : _GEN_4923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5228 = mask_5[2] ? byte_1282 : _GEN_4924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5229 = mask_5[3] ? byte_1283 : _GEN_4925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5230 = _GEN_8786 == 8'hc ? _GEN_5226 : _GEN_4922; // @[executor.scala 473:84]
  wire [7:0] _GEN_5231 = _GEN_8786 == 8'hc ? _GEN_5227 : _GEN_4923; // @[executor.scala 473:84]
  wire [7:0] _GEN_5232 = _GEN_8786 == 8'hc ? _GEN_5228 : _GEN_4924; // @[executor.scala 473:84]
  wire [7:0] _GEN_5233 = _GEN_8786 == 8'hc ? _GEN_5229 : _GEN_4925; // @[executor.scala 473:84]
  wire [7:0] _GEN_5234 = mask_5[0] ? byte_1280 : _GEN_4926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5235 = mask_5[1] ? byte_1281 : _GEN_4927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5236 = mask_5[2] ? byte_1282 : _GEN_4928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5237 = mask_5[3] ? byte_1283 : _GEN_4929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5238 = _GEN_8786 == 8'hd ? _GEN_5234 : _GEN_4926; // @[executor.scala 473:84]
  wire [7:0] _GEN_5239 = _GEN_8786 == 8'hd ? _GEN_5235 : _GEN_4927; // @[executor.scala 473:84]
  wire [7:0] _GEN_5240 = _GEN_8786 == 8'hd ? _GEN_5236 : _GEN_4928; // @[executor.scala 473:84]
  wire [7:0] _GEN_5241 = _GEN_8786 == 8'hd ? _GEN_5237 : _GEN_4929; // @[executor.scala 473:84]
  wire [7:0] _GEN_5242 = mask_5[0] ? byte_1280 : _GEN_4930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5243 = mask_5[1] ? byte_1281 : _GEN_4931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5244 = mask_5[2] ? byte_1282 : _GEN_4932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5245 = mask_5[3] ? byte_1283 : _GEN_4933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5246 = _GEN_8786 == 8'he ? _GEN_5242 : _GEN_4930; // @[executor.scala 473:84]
  wire [7:0] _GEN_5247 = _GEN_8786 == 8'he ? _GEN_5243 : _GEN_4931; // @[executor.scala 473:84]
  wire [7:0] _GEN_5248 = _GEN_8786 == 8'he ? _GEN_5244 : _GEN_4932; // @[executor.scala 473:84]
  wire [7:0] _GEN_5249 = _GEN_8786 == 8'he ? _GEN_5245 : _GEN_4933; // @[executor.scala 473:84]
  wire [7:0] _GEN_5250 = mask_5[0] ? byte_1280 : _GEN_4934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5251 = mask_5[1] ? byte_1281 : _GEN_4935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5252 = mask_5[2] ? byte_1282 : _GEN_4936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5253 = mask_5[3] ? byte_1283 : _GEN_4937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5254 = _GEN_8786 == 8'hf ? _GEN_5250 : _GEN_4934; // @[executor.scala 473:84]
  wire [7:0] _GEN_5255 = _GEN_8786 == 8'hf ? _GEN_5251 : _GEN_4935; // @[executor.scala 473:84]
  wire [7:0] _GEN_5256 = _GEN_8786 == 8'hf ? _GEN_5252 : _GEN_4936; // @[executor.scala 473:84]
  wire [7:0] _GEN_5257 = _GEN_8786 == 8'hf ? _GEN_5253 : _GEN_4937; // @[executor.scala 473:84]
  wire [7:0] _GEN_5258 = mask_5[0] ? byte_1280 : _GEN_4938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5259 = mask_5[1] ? byte_1281 : _GEN_4939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5260 = mask_5[2] ? byte_1282 : _GEN_4940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5261 = mask_5[3] ? byte_1283 : _GEN_4941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5262 = _GEN_8786 == 8'h10 ? _GEN_5258 : _GEN_4938; // @[executor.scala 473:84]
  wire [7:0] _GEN_5263 = _GEN_8786 == 8'h10 ? _GEN_5259 : _GEN_4939; // @[executor.scala 473:84]
  wire [7:0] _GEN_5264 = _GEN_8786 == 8'h10 ? _GEN_5260 : _GEN_4940; // @[executor.scala 473:84]
  wire [7:0] _GEN_5265 = _GEN_8786 == 8'h10 ? _GEN_5261 : _GEN_4941; // @[executor.scala 473:84]
  wire [7:0] _GEN_5266 = mask_5[0] ? byte_1280 : _GEN_4942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5267 = mask_5[1] ? byte_1281 : _GEN_4943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5268 = mask_5[2] ? byte_1282 : _GEN_4944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5269 = mask_5[3] ? byte_1283 : _GEN_4945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5270 = _GEN_8786 == 8'h11 ? _GEN_5266 : _GEN_4942; // @[executor.scala 473:84]
  wire [7:0] _GEN_5271 = _GEN_8786 == 8'h11 ? _GEN_5267 : _GEN_4943; // @[executor.scala 473:84]
  wire [7:0] _GEN_5272 = _GEN_8786 == 8'h11 ? _GEN_5268 : _GEN_4944; // @[executor.scala 473:84]
  wire [7:0] _GEN_5273 = _GEN_8786 == 8'h11 ? _GEN_5269 : _GEN_4945; // @[executor.scala 473:84]
  wire [7:0] _GEN_5274 = mask_5[0] ? byte_1280 : _GEN_4946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5275 = mask_5[1] ? byte_1281 : _GEN_4947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5276 = mask_5[2] ? byte_1282 : _GEN_4948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5277 = mask_5[3] ? byte_1283 : _GEN_4949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5278 = _GEN_8786 == 8'h12 ? _GEN_5274 : _GEN_4946; // @[executor.scala 473:84]
  wire [7:0] _GEN_5279 = _GEN_8786 == 8'h12 ? _GEN_5275 : _GEN_4947; // @[executor.scala 473:84]
  wire [7:0] _GEN_5280 = _GEN_8786 == 8'h12 ? _GEN_5276 : _GEN_4948; // @[executor.scala 473:84]
  wire [7:0] _GEN_5281 = _GEN_8786 == 8'h12 ? _GEN_5277 : _GEN_4949; // @[executor.scala 473:84]
  wire [7:0] _GEN_5282 = mask_5[0] ? byte_1280 : _GEN_4950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5283 = mask_5[1] ? byte_1281 : _GEN_4951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5284 = mask_5[2] ? byte_1282 : _GEN_4952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5285 = mask_5[3] ? byte_1283 : _GEN_4953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5286 = _GEN_8786 == 8'h13 ? _GEN_5282 : _GEN_4950; // @[executor.scala 473:84]
  wire [7:0] _GEN_5287 = _GEN_8786 == 8'h13 ? _GEN_5283 : _GEN_4951; // @[executor.scala 473:84]
  wire [7:0] _GEN_5288 = _GEN_8786 == 8'h13 ? _GEN_5284 : _GEN_4952; // @[executor.scala 473:84]
  wire [7:0] _GEN_5289 = _GEN_8786 == 8'h13 ? _GEN_5285 : _GEN_4953; // @[executor.scala 473:84]
  wire [7:0] _GEN_5290 = mask_5[0] ? byte_1280 : _GEN_4954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5291 = mask_5[1] ? byte_1281 : _GEN_4955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5292 = mask_5[2] ? byte_1282 : _GEN_4956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5293 = mask_5[3] ? byte_1283 : _GEN_4957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5294 = _GEN_8786 == 8'h14 ? _GEN_5290 : _GEN_4954; // @[executor.scala 473:84]
  wire [7:0] _GEN_5295 = _GEN_8786 == 8'h14 ? _GEN_5291 : _GEN_4955; // @[executor.scala 473:84]
  wire [7:0] _GEN_5296 = _GEN_8786 == 8'h14 ? _GEN_5292 : _GEN_4956; // @[executor.scala 473:84]
  wire [7:0] _GEN_5297 = _GEN_8786 == 8'h14 ? _GEN_5293 : _GEN_4957; // @[executor.scala 473:84]
  wire [7:0] _GEN_5298 = mask_5[0] ? byte_1280 : _GEN_4958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5299 = mask_5[1] ? byte_1281 : _GEN_4959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5300 = mask_5[2] ? byte_1282 : _GEN_4960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5301 = mask_5[3] ? byte_1283 : _GEN_4961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5302 = _GEN_8786 == 8'h15 ? _GEN_5298 : _GEN_4958; // @[executor.scala 473:84]
  wire [7:0] _GEN_5303 = _GEN_8786 == 8'h15 ? _GEN_5299 : _GEN_4959; // @[executor.scala 473:84]
  wire [7:0] _GEN_5304 = _GEN_8786 == 8'h15 ? _GEN_5300 : _GEN_4960; // @[executor.scala 473:84]
  wire [7:0] _GEN_5305 = _GEN_8786 == 8'h15 ? _GEN_5301 : _GEN_4961; // @[executor.scala 473:84]
  wire [7:0] _GEN_5306 = mask_5[0] ? byte_1280 : _GEN_4962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5307 = mask_5[1] ? byte_1281 : _GEN_4963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5308 = mask_5[2] ? byte_1282 : _GEN_4964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5309 = mask_5[3] ? byte_1283 : _GEN_4965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5310 = _GEN_8786 == 8'h16 ? _GEN_5306 : _GEN_4962; // @[executor.scala 473:84]
  wire [7:0] _GEN_5311 = _GEN_8786 == 8'h16 ? _GEN_5307 : _GEN_4963; // @[executor.scala 473:84]
  wire [7:0] _GEN_5312 = _GEN_8786 == 8'h16 ? _GEN_5308 : _GEN_4964; // @[executor.scala 473:84]
  wire [7:0] _GEN_5313 = _GEN_8786 == 8'h16 ? _GEN_5309 : _GEN_4965; // @[executor.scala 473:84]
  wire [7:0] _GEN_5314 = mask_5[0] ? byte_1280 : _GEN_4966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5315 = mask_5[1] ? byte_1281 : _GEN_4967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5316 = mask_5[2] ? byte_1282 : _GEN_4968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5317 = mask_5[3] ? byte_1283 : _GEN_4969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5318 = _GEN_8786 == 8'h17 ? _GEN_5314 : _GEN_4966; // @[executor.scala 473:84]
  wire [7:0] _GEN_5319 = _GEN_8786 == 8'h17 ? _GEN_5315 : _GEN_4967; // @[executor.scala 473:84]
  wire [7:0] _GEN_5320 = _GEN_8786 == 8'h17 ? _GEN_5316 : _GEN_4968; // @[executor.scala 473:84]
  wire [7:0] _GEN_5321 = _GEN_8786 == 8'h17 ? _GEN_5317 : _GEN_4969; // @[executor.scala 473:84]
  wire [7:0] _GEN_5322 = mask_5[0] ? byte_1280 : _GEN_4970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5323 = mask_5[1] ? byte_1281 : _GEN_4971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5324 = mask_5[2] ? byte_1282 : _GEN_4972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5325 = mask_5[3] ? byte_1283 : _GEN_4973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5326 = _GEN_8786 == 8'h18 ? _GEN_5322 : _GEN_4970; // @[executor.scala 473:84]
  wire [7:0] _GEN_5327 = _GEN_8786 == 8'h18 ? _GEN_5323 : _GEN_4971; // @[executor.scala 473:84]
  wire [7:0] _GEN_5328 = _GEN_8786 == 8'h18 ? _GEN_5324 : _GEN_4972; // @[executor.scala 473:84]
  wire [7:0] _GEN_5329 = _GEN_8786 == 8'h18 ? _GEN_5325 : _GEN_4973; // @[executor.scala 473:84]
  wire [7:0] _GEN_5330 = mask_5[0] ? byte_1280 : _GEN_4974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5331 = mask_5[1] ? byte_1281 : _GEN_4975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5332 = mask_5[2] ? byte_1282 : _GEN_4976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5333 = mask_5[3] ? byte_1283 : _GEN_4977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5334 = _GEN_8786 == 8'h19 ? _GEN_5330 : _GEN_4974; // @[executor.scala 473:84]
  wire [7:0] _GEN_5335 = _GEN_8786 == 8'h19 ? _GEN_5331 : _GEN_4975; // @[executor.scala 473:84]
  wire [7:0] _GEN_5336 = _GEN_8786 == 8'h19 ? _GEN_5332 : _GEN_4976; // @[executor.scala 473:84]
  wire [7:0] _GEN_5337 = _GEN_8786 == 8'h19 ? _GEN_5333 : _GEN_4977; // @[executor.scala 473:84]
  wire [7:0] _GEN_5338 = mask_5[0] ? byte_1280 : _GEN_4978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5339 = mask_5[1] ? byte_1281 : _GEN_4979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5340 = mask_5[2] ? byte_1282 : _GEN_4980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5341 = mask_5[3] ? byte_1283 : _GEN_4981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5342 = _GEN_8786 == 8'h1a ? _GEN_5338 : _GEN_4978; // @[executor.scala 473:84]
  wire [7:0] _GEN_5343 = _GEN_8786 == 8'h1a ? _GEN_5339 : _GEN_4979; // @[executor.scala 473:84]
  wire [7:0] _GEN_5344 = _GEN_8786 == 8'h1a ? _GEN_5340 : _GEN_4980; // @[executor.scala 473:84]
  wire [7:0] _GEN_5345 = _GEN_8786 == 8'h1a ? _GEN_5341 : _GEN_4981; // @[executor.scala 473:84]
  wire [7:0] _GEN_5346 = mask_5[0] ? byte_1280 : _GEN_4982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5347 = mask_5[1] ? byte_1281 : _GEN_4983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5348 = mask_5[2] ? byte_1282 : _GEN_4984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5349 = mask_5[3] ? byte_1283 : _GEN_4985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5350 = _GEN_8786 == 8'h1b ? _GEN_5346 : _GEN_4982; // @[executor.scala 473:84]
  wire [7:0] _GEN_5351 = _GEN_8786 == 8'h1b ? _GEN_5347 : _GEN_4983; // @[executor.scala 473:84]
  wire [7:0] _GEN_5352 = _GEN_8786 == 8'h1b ? _GEN_5348 : _GEN_4984; // @[executor.scala 473:84]
  wire [7:0] _GEN_5353 = _GEN_8786 == 8'h1b ? _GEN_5349 : _GEN_4985; // @[executor.scala 473:84]
  wire [7:0] _GEN_5354 = mask_5[0] ? byte_1280 : _GEN_4986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5355 = mask_5[1] ? byte_1281 : _GEN_4987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5356 = mask_5[2] ? byte_1282 : _GEN_4988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5357 = mask_5[3] ? byte_1283 : _GEN_4989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5358 = _GEN_8786 == 8'h1c ? _GEN_5354 : _GEN_4986; // @[executor.scala 473:84]
  wire [7:0] _GEN_5359 = _GEN_8786 == 8'h1c ? _GEN_5355 : _GEN_4987; // @[executor.scala 473:84]
  wire [7:0] _GEN_5360 = _GEN_8786 == 8'h1c ? _GEN_5356 : _GEN_4988; // @[executor.scala 473:84]
  wire [7:0] _GEN_5361 = _GEN_8786 == 8'h1c ? _GEN_5357 : _GEN_4989; // @[executor.scala 473:84]
  wire [7:0] _GEN_5362 = mask_5[0] ? byte_1280 : _GEN_4990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5363 = mask_5[1] ? byte_1281 : _GEN_4991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5364 = mask_5[2] ? byte_1282 : _GEN_4992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5365 = mask_5[3] ? byte_1283 : _GEN_4993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5366 = _GEN_8786 == 8'h1d ? _GEN_5362 : _GEN_4990; // @[executor.scala 473:84]
  wire [7:0] _GEN_5367 = _GEN_8786 == 8'h1d ? _GEN_5363 : _GEN_4991; // @[executor.scala 473:84]
  wire [7:0] _GEN_5368 = _GEN_8786 == 8'h1d ? _GEN_5364 : _GEN_4992; // @[executor.scala 473:84]
  wire [7:0] _GEN_5369 = _GEN_8786 == 8'h1d ? _GEN_5365 : _GEN_4993; // @[executor.scala 473:84]
  wire [7:0] _GEN_5370 = mask_5[0] ? byte_1280 : _GEN_4994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5371 = mask_5[1] ? byte_1281 : _GEN_4995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5372 = mask_5[2] ? byte_1282 : _GEN_4996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5373 = mask_5[3] ? byte_1283 : _GEN_4997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5374 = _GEN_8786 == 8'h1e ? _GEN_5370 : _GEN_4994; // @[executor.scala 473:84]
  wire [7:0] _GEN_5375 = _GEN_8786 == 8'h1e ? _GEN_5371 : _GEN_4995; // @[executor.scala 473:84]
  wire [7:0] _GEN_5376 = _GEN_8786 == 8'h1e ? _GEN_5372 : _GEN_4996; // @[executor.scala 473:84]
  wire [7:0] _GEN_5377 = _GEN_8786 == 8'h1e ? _GEN_5373 : _GEN_4997; // @[executor.scala 473:84]
  wire [7:0] _GEN_5378 = mask_5[0] ? byte_1280 : _GEN_4998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5379 = mask_5[1] ? byte_1281 : _GEN_4999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5380 = mask_5[2] ? byte_1282 : _GEN_5000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5381 = mask_5[3] ? byte_1283 : _GEN_5001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5382 = _GEN_8786 == 8'h1f ? _GEN_5378 : _GEN_4998; // @[executor.scala 473:84]
  wire [7:0] _GEN_5383 = _GEN_8786 == 8'h1f ? _GEN_5379 : _GEN_4999; // @[executor.scala 473:84]
  wire [7:0] _GEN_5384 = _GEN_8786 == 8'h1f ? _GEN_5380 : _GEN_5000; // @[executor.scala 473:84]
  wire [7:0] _GEN_5385 = _GEN_8786 == 8'h1f ? _GEN_5381 : _GEN_5001; // @[executor.scala 473:84]
  wire [7:0] _GEN_5386 = mask_5[0] ? byte_1280 : _GEN_5002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5387 = mask_5[1] ? byte_1281 : _GEN_5003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5388 = mask_5[2] ? byte_1282 : _GEN_5004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5389 = mask_5[3] ? byte_1283 : _GEN_5005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5390 = _GEN_8786 == 8'h20 ? _GEN_5386 : _GEN_5002; // @[executor.scala 473:84]
  wire [7:0] _GEN_5391 = _GEN_8786 == 8'h20 ? _GEN_5387 : _GEN_5003; // @[executor.scala 473:84]
  wire [7:0] _GEN_5392 = _GEN_8786 == 8'h20 ? _GEN_5388 : _GEN_5004; // @[executor.scala 473:84]
  wire [7:0] _GEN_5393 = _GEN_8786 == 8'h20 ? _GEN_5389 : _GEN_5005; // @[executor.scala 473:84]
  wire [7:0] _GEN_5394 = mask_5[0] ? byte_1280 : _GEN_5006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5395 = mask_5[1] ? byte_1281 : _GEN_5007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5396 = mask_5[2] ? byte_1282 : _GEN_5008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5397 = mask_5[3] ? byte_1283 : _GEN_5009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5398 = _GEN_8786 == 8'h21 ? _GEN_5394 : _GEN_5006; // @[executor.scala 473:84]
  wire [7:0] _GEN_5399 = _GEN_8786 == 8'h21 ? _GEN_5395 : _GEN_5007; // @[executor.scala 473:84]
  wire [7:0] _GEN_5400 = _GEN_8786 == 8'h21 ? _GEN_5396 : _GEN_5008; // @[executor.scala 473:84]
  wire [7:0] _GEN_5401 = _GEN_8786 == 8'h21 ? _GEN_5397 : _GEN_5009; // @[executor.scala 473:84]
  wire [7:0] _GEN_5402 = mask_5[0] ? byte_1280 : _GEN_5010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5403 = mask_5[1] ? byte_1281 : _GEN_5011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5404 = mask_5[2] ? byte_1282 : _GEN_5012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5405 = mask_5[3] ? byte_1283 : _GEN_5013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5406 = _GEN_8786 == 8'h22 ? _GEN_5402 : _GEN_5010; // @[executor.scala 473:84]
  wire [7:0] _GEN_5407 = _GEN_8786 == 8'h22 ? _GEN_5403 : _GEN_5011; // @[executor.scala 473:84]
  wire [7:0] _GEN_5408 = _GEN_8786 == 8'h22 ? _GEN_5404 : _GEN_5012; // @[executor.scala 473:84]
  wire [7:0] _GEN_5409 = _GEN_8786 == 8'h22 ? _GEN_5405 : _GEN_5013; // @[executor.scala 473:84]
  wire [7:0] _GEN_5410 = mask_5[0] ? byte_1280 : _GEN_5014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5411 = mask_5[1] ? byte_1281 : _GEN_5015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5412 = mask_5[2] ? byte_1282 : _GEN_5016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5413 = mask_5[3] ? byte_1283 : _GEN_5017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5414 = _GEN_8786 == 8'h23 ? _GEN_5410 : _GEN_5014; // @[executor.scala 473:84]
  wire [7:0] _GEN_5415 = _GEN_8786 == 8'h23 ? _GEN_5411 : _GEN_5015; // @[executor.scala 473:84]
  wire [7:0] _GEN_5416 = _GEN_8786 == 8'h23 ? _GEN_5412 : _GEN_5016; // @[executor.scala 473:84]
  wire [7:0] _GEN_5417 = _GEN_8786 == 8'h23 ? _GEN_5413 : _GEN_5017; // @[executor.scala 473:84]
  wire [7:0] _GEN_5418 = mask_5[0] ? byte_1280 : _GEN_5018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5419 = mask_5[1] ? byte_1281 : _GEN_5019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5420 = mask_5[2] ? byte_1282 : _GEN_5020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5421 = mask_5[3] ? byte_1283 : _GEN_5021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5422 = _GEN_8786 == 8'h24 ? _GEN_5418 : _GEN_5018; // @[executor.scala 473:84]
  wire [7:0] _GEN_5423 = _GEN_8786 == 8'h24 ? _GEN_5419 : _GEN_5019; // @[executor.scala 473:84]
  wire [7:0] _GEN_5424 = _GEN_8786 == 8'h24 ? _GEN_5420 : _GEN_5020; // @[executor.scala 473:84]
  wire [7:0] _GEN_5425 = _GEN_8786 == 8'h24 ? _GEN_5421 : _GEN_5021; // @[executor.scala 473:84]
  wire [7:0] _GEN_5426 = mask_5[0] ? byte_1280 : _GEN_5022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5427 = mask_5[1] ? byte_1281 : _GEN_5023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5428 = mask_5[2] ? byte_1282 : _GEN_5024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5429 = mask_5[3] ? byte_1283 : _GEN_5025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5430 = _GEN_8786 == 8'h25 ? _GEN_5426 : _GEN_5022; // @[executor.scala 473:84]
  wire [7:0] _GEN_5431 = _GEN_8786 == 8'h25 ? _GEN_5427 : _GEN_5023; // @[executor.scala 473:84]
  wire [7:0] _GEN_5432 = _GEN_8786 == 8'h25 ? _GEN_5428 : _GEN_5024; // @[executor.scala 473:84]
  wire [7:0] _GEN_5433 = _GEN_8786 == 8'h25 ? _GEN_5429 : _GEN_5025; // @[executor.scala 473:84]
  wire [7:0] _GEN_5434 = mask_5[0] ? byte_1280 : _GEN_5026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5435 = mask_5[1] ? byte_1281 : _GEN_5027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5436 = mask_5[2] ? byte_1282 : _GEN_5028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5437 = mask_5[3] ? byte_1283 : _GEN_5029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5438 = _GEN_8786 == 8'h26 ? _GEN_5434 : _GEN_5026; // @[executor.scala 473:84]
  wire [7:0] _GEN_5439 = _GEN_8786 == 8'h26 ? _GEN_5435 : _GEN_5027; // @[executor.scala 473:84]
  wire [7:0] _GEN_5440 = _GEN_8786 == 8'h26 ? _GEN_5436 : _GEN_5028; // @[executor.scala 473:84]
  wire [7:0] _GEN_5441 = _GEN_8786 == 8'h26 ? _GEN_5437 : _GEN_5029; // @[executor.scala 473:84]
  wire [7:0] _GEN_5442 = mask_5[0] ? byte_1280 : _GEN_5030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5443 = mask_5[1] ? byte_1281 : _GEN_5031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5444 = mask_5[2] ? byte_1282 : _GEN_5032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5445 = mask_5[3] ? byte_1283 : _GEN_5033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5446 = _GEN_8786 == 8'h27 ? _GEN_5442 : _GEN_5030; // @[executor.scala 473:84]
  wire [7:0] _GEN_5447 = _GEN_8786 == 8'h27 ? _GEN_5443 : _GEN_5031; // @[executor.scala 473:84]
  wire [7:0] _GEN_5448 = _GEN_8786 == 8'h27 ? _GEN_5444 : _GEN_5032; // @[executor.scala 473:84]
  wire [7:0] _GEN_5449 = _GEN_8786 == 8'h27 ? _GEN_5445 : _GEN_5033; // @[executor.scala 473:84]
  wire [7:0] _GEN_5450 = mask_5[0] ? byte_1280 : _GEN_5034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5451 = mask_5[1] ? byte_1281 : _GEN_5035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5452 = mask_5[2] ? byte_1282 : _GEN_5036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5453 = mask_5[3] ? byte_1283 : _GEN_5037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5454 = _GEN_8786 == 8'h28 ? _GEN_5450 : _GEN_5034; // @[executor.scala 473:84]
  wire [7:0] _GEN_5455 = _GEN_8786 == 8'h28 ? _GEN_5451 : _GEN_5035; // @[executor.scala 473:84]
  wire [7:0] _GEN_5456 = _GEN_8786 == 8'h28 ? _GEN_5452 : _GEN_5036; // @[executor.scala 473:84]
  wire [7:0] _GEN_5457 = _GEN_8786 == 8'h28 ? _GEN_5453 : _GEN_5037; // @[executor.scala 473:84]
  wire [7:0] _GEN_5458 = mask_5[0] ? byte_1280 : _GEN_5038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5459 = mask_5[1] ? byte_1281 : _GEN_5039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5460 = mask_5[2] ? byte_1282 : _GEN_5040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5461 = mask_5[3] ? byte_1283 : _GEN_5041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5462 = _GEN_8786 == 8'h29 ? _GEN_5458 : _GEN_5038; // @[executor.scala 473:84]
  wire [7:0] _GEN_5463 = _GEN_8786 == 8'h29 ? _GEN_5459 : _GEN_5039; // @[executor.scala 473:84]
  wire [7:0] _GEN_5464 = _GEN_8786 == 8'h29 ? _GEN_5460 : _GEN_5040; // @[executor.scala 473:84]
  wire [7:0] _GEN_5465 = _GEN_8786 == 8'h29 ? _GEN_5461 : _GEN_5041; // @[executor.scala 473:84]
  wire [7:0] _GEN_5466 = mask_5[0] ? byte_1280 : _GEN_5042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5467 = mask_5[1] ? byte_1281 : _GEN_5043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5468 = mask_5[2] ? byte_1282 : _GEN_5044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5469 = mask_5[3] ? byte_1283 : _GEN_5045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5470 = _GEN_8786 == 8'h2a ? _GEN_5466 : _GEN_5042; // @[executor.scala 473:84]
  wire [7:0] _GEN_5471 = _GEN_8786 == 8'h2a ? _GEN_5467 : _GEN_5043; // @[executor.scala 473:84]
  wire [7:0] _GEN_5472 = _GEN_8786 == 8'h2a ? _GEN_5468 : _GEN_5044; // @[executor.scala 473:84]
  wire [7:0] _GEN_5473 = _GEN_8786 == 8'h2a ? _GEN_5469 : _GEN_5045; // @[executor.scala 473:84]
  wire [7:0] _GEN_5474 = mask_5[0] ? byte_1280 : _GEN_5046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5475 = mask_5[1] ? byte_1281 : _GEN_5047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5476 = mask_5[2] ? byte_1282 : _GEN_5048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5477 = mask_5[3] ? byte_1283 : _GEN_5049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5478 = _GEN_8786 == 8'h2b ? _GEN_5474 : _GEN_5046; // @[executor.scala 473:84]
  wire [7:0] _GEN_5479 = _GEN_8786 == 8'h2b ? _GEN_5475 : _GEN_5047; // @[executor.scala 473:84]
  wire [7:0] _GEN_5480 = _GEN_8786 == 8'h2b ? _GEN_5476 : _GEN_5048; // @[executor.scala 473:84]
  wire [7:0] _GEN_5481 = _GEN_8786 == 8'h2b ? _GEN_5477 : _GEN_5049; // @[executor.scala 473:84]
  wire [7:0] _GEN_5482 = mask_5[0] ? byte_1280 : _GEN_5050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5483 = mask_5[1] ? byte_1281 : _GEN_5051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5484 = mask_5[2] ? byte_1282 : _GEN_5052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5485 = mask_5[3] ? byte_1283 : _GEN_5053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5486 = _GEN_8786 == 8'h2c ? _GEN_5482 : _GEN_5050; // @[executor.scala 473:84]
  wire [7:0] _GEN_5487 = _GEN_8786 == 8'h2c ? _GEN_5483 : _GEN_5051; // @[executor.scala 473:84]
  wire [7:0] _GEN_5488 = _GEN_8786 == 8'h2c ? _GEN_5484 : _GEN_5052; // @[executor.scala 473:84]
  wire [7:0] _GEN_5489 = _GEN_8786 == 8'h2c ? _GEN_5485 : _GEN_5053; // @[executor.scala 473:84]
  wire [7:0] _GEN_5490 = mask_5[0] ? byte_1280 : _GEN_5054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5491 = mask_5[1] ? byte_1281 : _GEN_5055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5492 = mask_5[2] ? byte_1282 : _GEN_5056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5493 = mask_5[3] ? byte_1283 : _GEN_5057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5494 = _GEN_8786 == 8'h2d ? _GEN_5490 : _GEN_5054; // @[executor.scala 473:84]
  wire [7:0] _GEN_5495 = _GEN_8786 == 8'h2d ? _GEN_5491 : _GEN_5055; // @[executor.scala 473:84]
  wire [7:0] _GEN_5496 = _GEN_8786 == 8'h2d ? _GEN_5492 : _GEN_5056; // @[executor.scala 473:84]
  wire [7:0] _GEN_5497 = _GEN_8786 == 8'h2d ? _GEN_5493 : _GEN_5057; // @[executor.scala 473:84]
  wire [7:0] _GEN_5498 = mask_5[0] ? byte_1280 : _GEN_5058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5499 = mask_5[1] ? byte_1281 : _GEN_5059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5500 = mask_5[2] ? byte_1282 : _GEN_5060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5501 = mask_5[3] ? byte_1283 : _GEN_5061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5502 = _GEN_8786 == 8'h2e ? _GEN_5498 : _GEN_5058; // @[executor.scala 473:84]
  wire [7:0] _GEN_5503 = _GEN_8786 == 8'h2e ? _GEN_5499 : _GEN_5059; // @[executor.scala 473:84]
  wire [7:0] _GEN_5504 = _GEN_8786 == 8'h2e ? _GEN_5500 : _GEN_5060; // @[executor.scala 473:84]
  wire [7:0] _GEN_5505 = _GEN_8786 == 8'h2e ? _GEN_5501 : _GEN_5061; // @[executor.scala 473:84]
  wire [7:0] _GEN_5506 = mask_5[0] ? byte_1280 : _GEN_5062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5507 = mask_5[1] ? byte_1281 : _GEN_5063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5508 = mask_5[2] ? byte_1282 : _GEN_5064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5509 = mask_5[3] ? byte_1283 : _GEN_5065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5510 = _GEN_8786 == 8'h2f ? _GEN_5506 : _GEN_5062; // @[executor.scala 473:84]
  wire [7:0] _GEN_5511 = _GEN_8786 == 8'h2f ? _GEN_5507 : _GEN_5063; // @[executor.scala 473:84]
  wire [7:0] _GEN_5512 = _GEN_8786 == 8'h2f ? _GEN_5508 : _GEN_5064; // @[executor.scala 473:84]
  wire [7:0] _GEN_5513 = _GEN_8786 == 8'h2f ? _GEN_5509 : _GEN_5065; // @[executor.scala 473:84]
  wire [7:0] _GEN_5514 = mask_5[0] ? byte_1280 : _GEN_5066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5515 = mask_5[1] ? byte_1281 : _GEN_5067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5516 = mask_5[2] ? byte_1282 : _GEN_5068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5517 = mask_5[3] ? byte_1283 : _GEN_5069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5518 = _GEN_8786 == 8'h30 ? _GEN_5514 : _GEN_5066; // @[executor.scala 473:84]
  wire [7:0] _GEN_5519 = _GEN_8786 == 8'h30 ? _GEN_5515 : _GEN_5067; // @[executor.scala 473:84]
  wire [7:0] _GEN_5520 = _GEN_8786 == 8'h30 ? _GEN_5516 : _GEN_5068; // @[executor.scala 473:84]
  wire [7:0] _GEN_5521 = _GEN_8786 == 8'h30 ? _GEN_5517 : _GEN_5069; // @[executor.scala 473:84]
  wire [7:0] _GEN_5522 = mask_5[0] ? byte_1280 : _GEN_5070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5523 = mask_5[1] ? byte_1281 : _GEN_5071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5524 = mask_5[2] ? byte_1282 : _GEN_5072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5525 = mask_5[3] ? byte_1283 : _GEN_5073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5526 = _GEN_8786 == 8'h31 ? _GEN_5522 : _GEN_5070; // @[executor.scala 473:84]
  wire [7:0] _GEN_5527 = _GEN_8786 == 8'h31 ? _GEN_5523 : _GEN_5071; // @[executor.scala 473:84]
  wire [7:0] _GEN_5528 = _GEN_8786 == 8'h31 ? _GEN_5524 : _GEN_5072; // @[executor.scala 473:84]
  wire [7:0] _GEN_5529 = _GEN_8786 == 8'h31 ? _GEN_5525 : _GEN_5073; // @[executor.scala 473:84]
  wire [7:0] _GEN_5530 = mask_5[0] ? byte_1280 : _GEN_5074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5531 = mask_5[1] ? byte_1281 : _GEN_5075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5532 = mask_5[2] ? byte_1282 : _GEN_5076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5533 = mask_5[3] ? byte_1283 : _GEN_5077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5534 = _GEN_8786 == 8'h32 ? _GEN_5530 : _GEN_5074; // @[executor.scala 473:84]
  wire [7:0] _GEN_5535 = _GEN_8786 == 8'h32 ? _GEN_5531 : _GEN_5075; // @[executor.scala 473:84]
  wire [7:0] _GEN_5536 = _GEN_8786 == 8'h32 ? _GEN_5532 : _GEN_5076; // @[executor.scala 473:84]
  wire [7:0] _GEN_5537 = _GEN_8786 == 8'h32 ? _GEN_5533 : _GEN_5077; // @[executor.scala 473:84]
  wire [7:0] _GEN_5538 = mask_5[0] ? byte_1280 : _GEN_5078; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5539 = mask_5[1] ? byte_1281 : _GEN_5079; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5540 = mask_5[2] ? byte_1282 : _GEN_5080; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5541 = mask_5[3] ? byte_1283 : _GEN_5081; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5542 = _GEN_8786 == 8'h33 ? _GEN_5538 : _GEN_5078; // @[executor.scala 473:84]
  wire [7:0] _GEN_5543 = _GEN_8786 == 8'h33 ? _GEN_5539 : _GEN_5079; // @[executor.scala 473:84]
  wire [7:0] _GEN_5544 = _GEN_8786 == 8'h33 ? _GEN_5540 : _GEN_5080; // @[executor.scala 473:84]
  wire [7:0] _GEN_5545 = _GEN_8786 == 8'h33 ? _GEN_5541 : _GEN_5081; // @[executor.scala 473:84]
  wire [7:0] _GEN_5546 = mask_5[0] ? byte_1280 : _GEN_5082; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5547 = mask_5[1] ? byte_1281 : _GEN_5083; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5548 = mask_5[2] ? byte_1282 : _GEN_5084; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5549 = mask_5[3] ? byte_1283 : _GEN_5085; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5550 = _GEN_8786 == 8'h34 ? _GEN_5546 : _GEN_5082; // @[executor.scala 473:84]
  wire [7:0] _GEN_5551 = _GEN_8786 == 8'h34 ? _GEN_5547 : _GEN_5083; // @[executor.scala 473:84]
  wire [7:0] _GEN_5552 = _GEN_8786 == 8'h34 ? _GEN_5548 : _GEN_5084; // @[executor.scala 473:84]
  wire [7:0] _GEN_5553 = _GEN_8786 == 8'h34 ? _GEN_5549 : _GEN_5085; // @[executor.scala 473:84]
  wire [7:0] _GEN_5554 = mask_5[0] ? byte_1280 : _GEN_5086; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5555 = mask_5[1] ? byte_1281 : _GEN_5087; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5556 = mask_5[2] ? byte_1282 : _GEN_5088; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5557 = mask_5[3] ? byte_1283 : _GEN_5089; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5558 = _GEN_8786 == 8'h35 ? _GEN_5554 : _GEN_5086; // @[executor.scala 473:84]
  wire [7:0] _GEN_5559 = _GEN_8786 == 8'h35 ? _GEN_5555 : _GEN_5087; // @[executor.scala 473:84]
  wire [7:0] _GEN_5560 = _GEN_8786 == 8'h35 ? _GEN_5556 : _GEN_5088; // @[executor.scala 473:84]
  wire [7:0] _GEN_5561 = _GEN_8786 == 8'h35 ? _GEN_5557 : _GEN_5089; // @[executor.scala 473:84]
  wire [7:0] _GEN_5562 = mask_5[0] ? byte_1280 : _GEN_5090; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5563 = mask_5[1] ? byte_1281 : _GEN_5091; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5564 = mask_5[2] ? byte_1282 : _GEN_5092; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5565 = mask_5[3] ? byte_1283 : _GEN_5093; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5566 = _GEN_8786 == 8'h36 ? _GEN_5562 : _GEN_5090; // @[executor.scala 473:84]
  wire [7:0] _GEN_5567 = _GEN_8786 == 8'h36 ? _GEN_5563 : _GEN_5091; // @[executor.scala 473:84]
  wire [7:0] _GEN_5568 = _GEN_8786 == 8'h36 ? _GEN_5564 : _GEN_5092; // @[executor.scala 473:84]
  wire [7:0] _GEN_5569 = _GEN_8786 == 8'h36 ? _GEN_5565 : _GEN_5093; // @[executor.scala 473:84]
  wire [7:0] _GEN_5570 = mask_5[0] ? byte_1280 : _GEN_5094; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5571 = mask_5[1] ? byte_1281 : _GEN_5095; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5572 = mask_5[2] ? byte_1282 : _GEN_5096; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5573 = mask_5[3] ? byte_1283 : _GEN_5097; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5574 = _GEN_8786 == 8'h37 ? _GEN_5570 : _GEN_5094; // @[executor.scala 473:84]
  wire [7:0] _GEN_5575 = _GEN_8786 == 8'h37 ? _GEN_5571 : _GEN_5095; // @[executor.scala 473:84]
  wire [7:0] _GEN_5576 = _GEN_8786 == 8'h37 ? _GEN_5572 : _GEN_5096; // @[executor.scala 473:84]
  wire [7:0] _GEN_5577 = _GEN_8786 == 8'h37 ? _GEN_5573 : _GEN_5097; // @[executor.scala 473:84]
  wire [7:0] _GEN_5578 = mask_5[0] ? byte_1280 : _GEN_5098; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5579 = mask_5[1] ? byte_1281 : _GEN_5099; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5580 = mask_5[2] ? byte_1282 : _GEN_5100; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5581 = mask_5[3] ? byte_1283 : _GEN_5101; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5582 = _GEN_8786 == 8'h38 ? _GEN_5578 : _GEN_5098; // @[executor.scala 473:84]
  wire [7:0] _GEN_5583 = _GEN_8786 == 8'h38 ? _GEN_5579 : _GEN_5099; // @[executor.scala 473:84]
  wire [7:0] _GEN_5584 = _GEN_8786 == 8'h38 ? _GEN_5580 : _GEN_5100; // @[executor.scala 473:84]
  wire [7:0] _GEN_5585 = _GEN_8786 == 8'h38 ? _GEN_5581 : _GEN_5101; // @[executor.scala 473:84]
  wire [7:0] _GEN_5586 = mask_5[0] ? byte_1280 : _GEN_5102; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5587 = mask_5[1] ? byte_1281 : _GEN_5103; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5588 = mask_5[2] ? byte_1282 : _GEN_5104; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5589 = mask_5[3] ? byte_1283 : _GEN_5105; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5590 = _GEN_8786 == 8'h39 ? _GEN_5586 : _GEN_5102; // @[executor.scala 473:84]
  wire [7:0] _GEN_5591 = _GEN_8786 == 8'h39 ? _GEN_5587 : _GEN_5103; // @[executor.scala 473:84]
  wire [7:0] _GEN_5592 = _GEN_8786 == 8'h39 ? _GEN_5588 : _GEN_5104; // @[executor.scala 473:84]
  wire [7:0] _GEN_5593 = _GEN_8786 == 8'h39 ? _GEN_5589 : _GEN_5105; // @[executor.scala 473:84]
  wire [7:0] _GEN_5594 = mask_5[0] ? byte_1280 : _GEN_5106; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5595 = mask_5[1] ? byte_1281 : _GEN_5107; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5596 = mask_5[2] ? byte_1282 : _GEN_5108; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5597 = mask_5[3] ? byte_1283 : _GEN_5109; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5598 = _GEN_8786 == 8'h3a ? _GEN_5594 : _GEN_5106; // @[executor.scala 473:84]
  wire [7:0] _GEN_5599 = _GEN_8786 == 8'h3a ? _GEN_5595 : _GEN_5107; // @[executor.scala 473:84]
  wire [7:0] _GEN_5600 = _GEN_8786 == 8'h3a ? _GEN_5596 : _GEN_5108; // @[executor.scala 473:84]
  wire [7:0] _GEN_5601 = _GEN_8786 == 8'h3a ? _GEN_5597 : _GEN_5109; // @[executor.scala 473:84]
  wire [7:0] _GEN_5602 = mask_5[0] ? byte_1280 : _GEN_5110; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5603 = mask_5[1] ? byte_1281 : _GEN_5111; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5604 = mask_5[2] ? byte_1282 : _GEN_5112; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5605 = mask_5[3] ? byte_1283 : _GEN_5113; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5606 = _GEN_8786 == 8'h3b ? _GEN_5602 : _GEN_5110; // @[executor.scala 473:84]
  wire [7:0] _GEN_5607 = _GEN_8786 == 8'h3b ? _GEN_5603 : _GEN_5111; // @[executor.scala 473:84]
  wire [7:0] _GEN_5608 = _GEN_8786 == 8'h3b ? _GEN_5604 : _GEN_5112; // @[executor.scala 473:84]
  wire [7:0] _GEN_5609 = _GEN_8786 == 8'h3b ? _GEN_5605 : _GEN_5113; // @[executor.scala 473:84]
  wire [7:0] _GEN_5610 = mask_5[0] ? byte_1280 : _GEN_5114; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5611 = mask_5[1] ? byte_1281 : _GEN_5115; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5612 = mask_5[2] ? byte_1282 : _GEN_5116; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5613 = mask_5[3] ? byte_1283 : _GEN_5117; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5614 = _GEN_8786 == 8'h3c ? _GEN_5610 : _GEN_5114; // @[executor.scala 473:84]
  wire [7:0] _GEN_5615 = _GEN_8786 == 8'h3c ? _GEN_5611 : _GEN_5115; // @[executor.scala 473:84]
  wire [7:0] _GEN_5616 = _GEN_8786 == 8'h3c ? _GEN_5612 : _GEN_5116; // @[executor.scala 473:84]
  wire [7:0] _GEN_5617 = _GEN_8786 == 8'h3c ? _GEN_5613 : _GEN_5117; // @[executor.scala 473:84]
  wire [7:0] _GEN_5618 = mask_5[0] ? byte_1280 : _GEN_5118; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5619 = mask_5[1] ? byte_1281 : _GEN_5119; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5620 = mask_5[2] ? byte_1282 : _GEN_5120; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5621 = mask_5[3] ? byte_1283 : _GEN_5121; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5622 = _GEN_8786 == 8'h3d ? _GEN_5618 : _GEN_5118; // @[executor.scala 473:84]
  wire [7:0] _GEN_5623 = _GEN_8786 == 8'h3d ? _GEN_5619 : _GEN_5119; // @[executor.scala 473:84]
  wire [7:0] _GEN_5624 = _GEN_8786 == 8'h3d ? _GEN_5620 : _GEN_5120; // @[executor.scala 473:84]
  wire [7:0] _GEN_5625 = _GEN_8786 == 8'h3d ? _GEN_5621 : _GEN_5121; // @[executor.scala 473:84]
  wire [7:0] _GEN_5626 = mask_5[0] ? byte_1280 : _GEN_5122; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5627 = mask_5[1] ? byte_1281 : _GEN_5123; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5628 = mask_5[2] ? byte_1282 : _GEN_5124; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5629 = mask_5[3] ? byte_1283 : _GEN_5125; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5630 = _GEN_8786 == 8'h3e ? _GEN_5626 : _GEN_5122; // @[executor.scala 473:84]
  wire [7:0] _GEN_5631 = _GEN_8786 == 8'h3e ? _GEN_5627 : _GEN_5123; // @[executor.scala 473:84]
  wire [7:0] _GEN_5632 = _GEN_8786 == 8'h3e ? _GEN_5628 : _GEN_5124; // @[executor.scala 473:84]
  wire [7:0] _GEN_5633 = _GEN_8786 == 8'h3e ? _GEN_5629 : _GEN_5125; // @[executor.scala 473:84]
  wire [7:0] _GEN_5634 = mask_5[0] ? byte_1280 : _GEN_5126; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5635 = mask_5[1] ? byte_1281 : _GEN_5127; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5636 = mask_5[2] ? byte_1282 : _GEN_5128; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5637 = mask_5[3] ? byte_1283 : _GEN_5129; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5638 = _GEN_8786 == 8'h3f ? _GEN_5634 : _GEN_5126; // @[executor.scala 473:84]
  wire [7:0] _GEN_5639 = _GEN_8786 == 8'h3f ? _GEN_5635 : _GEN_5127; // @[executor.scala 473:84]
  wire [7:0] _GEN_5640 = _GEN_8786 == 8'h3f ? _GEN_5636 : _GEN_5128; // @[executor.scala 473:84]
  wire [7:0] _GEN_5641 = _GEN_8786 == 8'h3f ? _GEN_5637 : _GEN_5129; // @[executor.scala 473:84]
  wire [7:0] _GEN_5642 = opcode_5 != 4'h0 ? _GEN_5134 : _GEN_4874; // @[executor.scala 470:55]
  wire [7:0] _GEN_5643 = opcode_5 != 4'h0 ? _GEN_5135 : _GEN_4875; // @[executor.scala 470:55]
  wire [7:0] _GEN_5644 = opcode_5 != 4'h0 ? _GEN_5136 : _GEN_4876; // @[executor.scala 470:55]
  wire [7:0] _GEN_5645 = opcode_5 != 4'h0 ? _GEN_5137 : _GEN_4877; // @[executor.scala 470:55]
  wire [7:0] _GEN_5646 = opcode_5 != 4'h0 ? _GEN_5142 : _GEN_4878; // @[executor.scala 470:55]
  wire [7:0] _GEN_5647 = opcode_5 != 4'h0 ? _GEN_5143 : _GEN_4879; // @[executor.scala 470:55]
  wire [7:0] _GEN_5648 = opcode_5 != 4'h0 ? _GEN_5144 : _GEN_4880; // @[executor.scala 470:55]
  wire [7:0] _GEN_5649 = opcode_5 != 4'h0 ? _GEN_5145 : _GEN_4881; // @[executor.scala 470:55]
  wire [7:0] _GEN_5650 = opcode_5 != 4'h0 ? _GEN_5150 : _GEN_4882; // @[executor.scala 470:55]
  wire [7:0] _GEN_5651 = opcode_5 != 4'h0 ? _GEN_5151 : _GEN_4883; // @[executor.scala 470:55]
  wire [7:0] _GEN_5652 = opcode_5 != 4'h0 ? _GEN_5152 : _GEN_4884; // @[executor.scala 470:55]
  wire [7:0] _GEN_5653 = opcode_5 != 4'h0 ? _GEN_5153 : _GEN_4885; // @[executor.scala 470:55]
  wire [7:0] _GEN_5654 = opcode_5 != 4'h0 ? _GEN_5158 : _GEN_4886; // @[executor.scala 470:55]
  wire [7:0] _GEN_5655 = opcode_5 != 4'h0 ? _GEN_5159 : _GEN_4887; // @[executor.scala 470:55]
  wire [7:0] _GEN_5656 = opcode_5 != 4'h0 ? _GEN_5160 : _GEN_4888; // @[executor.scala 470:55]
  wire [7:0] _GEN_5657 = opcode_5 != 4'h0 ? _GEN_5161 : _GEN_4889; // @[executor.scala 470:55]
  wire [7:0] _GEN_5658 = opcode_5 != 4'h0 ? _GEN_5166 : _GEN_4890; // @[executor.scala 470:55]
  wire [7:0] _GEN_5659 = opcode_5 != 4'h0 ? _GEN_5167 : _GEN_4891; // @[executor.scala 470:55]
  wire [7:0] _GEN_5660 = opcode_5 != 4'h0 ? _GEN_5168 : _GEN_4892; // @[executor.scala 470:55]
  wire [7:0] _GEN_5661 = opcode_5 != 4'h0 ? _GEN_5169 : _GEN_4893; // @[executor.scala 470:55]
  wire [7:0] _GEN_5662 = opcode_5 != 4'h0 ? _GEN_5174 : _GEN_4894; // @[executor.scala 470:55]
  wire [7:0] _GEN_5663 = opcode_5 != 4'h0 ? _GEN_5175 : _GEN_4895; // @[executor.scala 470:55]
  wire [7:0] _GEN_5664 = opcode_5 != 4'h0 ? _GEN_5176 : _GEN_4896; // @[executor.scala 470:55]
  wire [7:0] _GEN_5665 = opcode_5 != 4'h0 ? _GEN_5177 : _GEN_4897; // @[executor.scala 470:55]
  wire [7:0] _GEN_5666 = opcode_5 != 4'h0 ? _GEN_5182 : _GEN_4898; // @[executor.scala 470:55]
  wire [7:0] _GEN_5667 = opcode_5 != 4'h0 ? _GEN_5183 : _GEN_4899; // @[executor.scala 470:55]
  wire [7:0] _GEN_5668 = opcode_5 != 4'h0 ? _GEN_5184 : _GEN_4900; // @[executor.scala 470:55]
  wire [7:0] _GEN_5669 = opcode_5 != 4'h0 ? _GEN_5185 : _GEN_4901; // @[executor.scala 470:55]
  wire [7:0] _GEN_5670 = opcode_5 != 4'h0 ? _GEN_5190 : _GEN_4902; // @[executor.scala 470:55]
  wire [7:0] _GEN_5671 = opcode_5 != 4'h0 ? _GEN_5191 : _GEN_4903; // @[executor.scala 470:55]
  wire [7:0] _GEN_5672 = opcode_5 != 4'h0 ? _GEN_5192 : _GEN_4904; // @[executor.scala 470:55]
  wire [7:0] _GEN_5673 = opcode_5 != 4'h0 ? _GEN_5193 : _GEN_4905; // @[executor.scala 470:55]
  wire [7:0] _GEN_5674 = opcode_5 != 4'h0 ? _GEN_5198 : _GEN_4906; // @[executor.scala 470:55]
  wire [7:0] _GEN_5675 = opcode_5 != 4'h0 ? _GEN_5199 : _GEN_4907; // @[executor.scala 470:55]
  wire [7:0] _GEN_5676 = opcode_5 != 4'h0 ? _GEN_5200 : _GEN_4908; // @[executor.scala 470:55]
  wire [7:0] _GEN_5677 = opcode_5 != 4'h0 ? _GEN_5201 : _GEN_4909; // @[executor.scala 470:55]
  wire [7:0] _GEN_5678 = opcode_5 != 4'h0 ? _GEN_5206 : _GEN_4910; // @[executor.scala 470:55]
  wire [7:0] _GEN_5679 = opcode_5 != 4'h0 ? _GEN_5207 : _GEN_4911; // @[executor.scala 470:55]
  wire [7:0] _GEN_5680 = opcode_5 != 4'h0 ? _GEN_5208 : _GEN_4912; // @[executor.scala 470:55]
  wire [7:0] _GEN_5681 = opcode_5 != 4'h0 ? _GEN_5209 : _GEN_4913; // @[executor.scala 470:55]
  wire [7:0] _GEN_5682 = opcode_5 != 4'h0 ? _GEN_5214 : _GEN_4914; // @[executor.scala 470:55]
  wire [7:0] _GEN_5683 = opcode_5 != 4'h0 ? _GEN_5215 : _GEN_4915; // @[executor.scala 470:55]
  wire [7:0] _GEN_5684 = opcode_5 != 4'h0 ? _GEN_5216 : _GEN_4916; // @[executor.scala 470:55]
  wire [7:0] _GEN_5685 = opcode_5 != 4'h0 ? _GEN_5217 : _GEN_4917; // @[executor.scala 470:55]
  wire [7:0] _GEN_5686 = opcode_5 != 4'h0 ? _GEN_5222 : _GEN_4918; // @[executor.scala 470:55]
  wire [7:0] _GEN_5687 = opcode_5 != 4'h0 ? _GEN_5223 : _GEN_4919; // @[executor.scala 470:55]
  wire [7:0] _GEN_5688 = opcode_5 != 4'h0 ? _GEN_5224 : _GEN_4920; // @[executor.scala 470:55]
  wire [7:0] _GEN_5689 = opcode_5 != 4'h0 ? _GEN_5225 : _GEN_4921; // @[executor.scala 470:55]
  wire [7:0] _GEN_5690 = opcode_5 != 4'h0 ? _GEN_5230 : _GEN_4922; // @[executor.scala 470:55]
  wire [7:0] _GEN_5691 = opcode_5 != 4'h0 ? _GEN_5231 : _GEN_4923; // @[executor.scala 470:55]
  wire [7:0] _GEN_5692 = opcode_5 != 4'h0 ? _GEN_5232 : _GEN_4924; // @[executor.scala 470:55]
  wire [7:0] _GEN_5693 = opcode_5 != 4'h0 ? _GEN_5233 : _GEN_4925; // @[executor.scala 470:55]
  wire [7:0] _GEN_5694 = opcode_5 != 4'h0 ? _GEN_5238 : _GEN_4926; // @[executor.scala 470:55]
  wire [7:0] _GEN_5695 = opcode_5 != 4'h0 ? _GEN_5239 : _GEN_4927; // @[executor.scala 470:55]
  wire [7:0] _GEN_5696 = opcode_5 != 4'h0 ? _GEN_5240 : _GEN_4928; // @[executor.scala 470:55]
  wire [7:0] _GEN_5697 = opcode_5 != 4'h0 ? _GEN_5241 : _GEN_4929; // @[executor.scala 470:55]
  wire [7:0] _GEN_5698 = opcode_5 != 4'h0 ? _GEN_5246 : _GEN_4930; // @[executor.scala 470:55]
  wire [7:0] _GEN_5699 = opcode_5 != 4'h0 ? _GEN_5247 : _GEN_4931; // @[executor.scala 470:55]
  wire [7:0] _GEN_5700 = opcode_5 != 4'h0 ? _GEN_5248 : _GEN_4932; // @[executor.scala 470:55]
  wire [7:0] _GEN_5701 = opcode_5 != 4'h0 ? _GEN_5249 : _GEN_4933; // @[executor.scala 470:55]
  wire [7:0] _GEN_5702 = opcode_5 != 4'h0 ? _GEN_5254 : _GEN_4934; // @[executor.scala 470:55]
  wire [7:0] _GEN_5703 = opcode_5 != 4'h0 ? _GEN_5255 : _GEN_4935; // @[executor.scala 470:55]
  wire [7:0] _GEN_5704 = opcode_5 != 4'h0 ? _GEN_5256 : _GEN_4936; // @[executor.scala 470:55]
  wire [7:0] _GEN_5705 = opcode_5 != 4'h0 ? _GEN_5257 : _GEN_4937; // @[executor.scala 470:55]
  wire [7:0] _GEN_5706 = opcode_5 != 4'h0 ? _GEN_5262 : _GEN_4938; // @[executor.scala 470:55]
  wire [7:0] _GEN_5707 = opcode_5 != 4'h0 ? _GEN_5263 : _GEN_4939; // @[executor.scala 470:55]
  wire [7:0] _GEN_5708 = opcode_5 != 4'h0 ? _GEN_5264 : _GEN_4940; // @[executor.scala 470:55]
  wire [7:0] _GEN_5709 = opcode_5 != 4'h0 ? _GEN_5265 : _GEN_4941; // @[executor.scala 470:55]
  wire [7:0] _GEN_5710 = opcode_5 != 4'h0 ? _GEN_5270 : _GEN_4942; // @[executor.scala 470:55]
  wire [7:0] _GEN_5711 = opcode_5 != 4'h0 ? _GEN_5271 : _GEN_4943; // @[executor.scala 470:55]
  wire [7:0] _GEN_5712 = opcode_5 != 4'h0 ? _GEN_5272 : _GEN_4944; // @[executor.scala 470:55]
  wire [7:0] _GEN_5713 = opcode_5 != 4'h0 ? _GEN_5273 : _GEN_4945; // @[executor.scala 470:55]
  wire [7:0] _GEN_5714 = opcode_5 != 4'h0 ? _GEN_5278 : _GEN_4946; // @[executor.scala 470:55]
  wire [7:0] _GEN_5715 = opcode_5 != 4'h0 ? _GEN_5279 : _GEN_4947; // @[executor.scala 470:55]
  wire [7:0] _GEN_5716 = opcode_5 != 4'h0 ? _GEN_5280 : _GEN_4948; // @[executor.scala 470:55]
  wire [7:0] _GEN_5717 = opcode_5 != 4'h0 ? _GEN_5281 : _GEN_4949; // @[executor.scala 470:55]
  wire [7:0] _GEN_5718 = opcode_5 != 4'h0 ? _GEN_5286 : _GEN_4950; // @[executor.scala 470:55]
  wire [7:0] _GEN_5719 = opcode_5 != 4'h0 ? _GEN_5287 : _GEN_4951; // @[executor.scala 470:55]
  wire [7:0] _GEN_5720 = opcode_5 != 4'h0 ? _GEN_5288 : _GEN_4952; // @[executor.scala 470:55]
  wire [7:0] _GEN_5721 = opcode_5 != 4'h0 ? _GEN_5289 : _GEN_4953; // @[executor.scala 470:55]
  wire [7:0] _GEN_5722 = opcode_5 != 4'h0 ? _GEN_5294 : _GEN_4954; // @[executor.scala 470:55]
  wire [7:0] _GEN_5723 = opcode_5 != 4'h0 ? _GEN_5295 : _GEN_4955; // @[executor.scala 470:55]
  wire [7:0] _GEN_5724 = opcode_5 != 4'h0 ? _GEN_5296 : _GEN_4956; // @[executor.scala 470:55]
  wire [7:0] _GEN_5725 = opcode_5 != 4'h0 ? _GEN_5297 : _GEN_4957; // @[executor.scala 470:55]
  wire [7:0] _GEN_5726 = opcode_5 != 4'h0 ? _GEN_5302 : _GEN_4958; // @[executor.scala 470:55]
  wire [7:0] _GEN_5727 = opcode_5 != 4'h0 ? _GEN_5303 : _GEN_4959; // @[executor.scala 470:55]
  wire [7:0] _GEN_5728 = opcode_5 != 4'h0 ? _GEN_5304 : _GEN_4960; // @[executor.scala 470:55]
  wire [7:0] _GEN_5729 = opcode_5 != 4'h0 ? _GEN_5305 : _GEN_4961; // @[executor.scala 470:55]
  wire [7:0] _GEN_5730 = opcode_5 != 4'h0 ? _GEN_5310 : _GEN_4962; // @[executor.scala 470:55]
  wire [7:0] _GEN_5731 = opcode_5 != 4'h0 ? _GEN_5311 : _GEN_4963; // @[executor.scala 470:55]
  wire [7:0] _GEN_5732 = opcode_5 != 4'h0 ? _GEN_5312 : _GEN_4964; // @[executor.scala 470:55]
  wire [7:0] _GEN_5733 = opcode_5 != 4'h0 ? _GEN_5313 : _GEN_4965; // @[executor.scala 470:55]
  wire [7:0] _GEN_5734 = opcode_5 != 4'h0 ? _GEN_5318 : _GEN_4966; // @[executor.scala 470:55]
  wire [7:0] _GEN_5735 = opcode_5 != 4'h0 ? _GEN_5319 : _GEN_4967; // @[executor.scala 470:55]
  wire [7:0] _GEN_5736 = opcode_5 != 4'h0 ? _GEN_5320 : _GEN_4968; // @[executor.scala 470:55]
  wire [7:0] _GEN_5737 = opcode_5 != 4'h0 ? _GEN_5321 : _GEN_4969; // @[executor.scala 470:55]
  wire [7:0] _GEN_5738 = opcode_5 != 4'h0 ? _GEN_5326 : _GEN_4970; // @[executor.scala 470:55]
  wire [7:0] _GEN_5739 = opcode_5 != 4'h0 ? _GEN_5327 : _GEN_4971; // @[executor.scala 470:55]
  wire [7:0] _GEN_5740 = opcode_5 != 4'h0 ? _GEN_5328 : _GEN_4972; // @[executor.scala 470:55]
  wire [7:0] _GEN_5741 = opcode_5 != 4'h0 ? _GEN_5329 : _GEN_4973; // @[executor.scala 470:55]
  wire [7:0] _GEN_5742 = opcode_5 != 4'h0 ? _GEN_5334 : _GEN_4974; // @[executor.scala 470:55]
  wire [7:0] _GEN_5743 = opcode_5 != 4'h0 ? _GEN_5335 : _GEN_4975; // @[executor.scala 470:55]
  wire [7:0] _GEN_5744 = opcode_5 != 4'h0 ? _GEN_5336 : _GEN_4976; // @[executor.scala 470:55]
  wire [7:0] _GEN_5745 = opcode_5 != 4'h0 ? _GEN_5337 : _GEN_4977; // @[executor.scala 470:55]
  wire [7:0] _GEN_5746 = opcode_5 != 4'h0 ? _GEN_5342 : _GEN_4978; // @[executor.scala 470:55]
  wire [7:0] _GEN_5747 = opcode_5 != 4'h0 ? _GEN_5343 : _GEN_4979; // @[executor.scala 470:55]
  wire [7:0] _GEN_5748 = opcode_5 != 4'h0 ? _GEN_5344 : _GEN_4980; // @[executor.scala 470:55]
  wire [7:0] _GEN_5749 = opcode_5 != 4'h0 ? _GEN_5345 : _GEN_4981; // @[executor.scala 470:55]
  wire [7:0] _GEN_5750 = opcode_5 != 4'h0 ? _GEN_5350 : _GEN_4982; // @[executor.scala 470:55]
  wire [7:0] _GEN_5751 = opcode_5 != 4'h0 ? _GEN_5351 : _GEN_4983; // @[executor.scala 470:55]
  wire [7:0] _GEN_5752 = opcode_5 != 4'h0 ? _GEN_5352 : _GEN_4984; // @[executor.scala 470:55]
  wire [7:0] _GEN_5753 = opcode_5 != 4'h0 ? _GEN_5353 : _GEN_4985; // @[executor.scala 470:55]
  wire [7:0] _GEN_5754 = opcode_5 != 4'h0 ? _GEN_5358 : _GEN_4986; // @[executor.scala 470:55]
  wire [7:0] _GEN_5755 = opcode_5 != 4'h0 ? _GEN_5359 : _GEN_4987; // @[executor.scala 470:55]
  wire [7:0] _GEN_5756 = opcode_5 != 4'h0 ? _GEN_5360 : _GEN_4988; // @[executor.scala 470:55]
  wire [7:0] _GEN_5757 = opcode_5 != 4'h0 ? _GEN_5361 : _GEN_4989; // @[executor.scala 470:55]
  wire [7:0] _GEN_5758 = opcode_5 != 4'h0 ? _GEN_5366 : _GEN_4990; // @[executor.scala 470:55]
  wire [7:0] _GEN_5759 = opcode_5 != 4'h0 ? _GEN_5367 : _GEN_4991; // @[executor.scala 470:55]
  wire [7:0] _GEN_5760 = opcode_5 != 4'h0 ? _GEN_5368 : _GEN_4992; // @[executor.scala 470:55]
  wire [7:0] _GEN_5761 = opcode_5 != 4'h0 ? _GEN_5369 : _GEN_4993; // @[executor.scala 470:55]
  wire [7:0] _GEN_5762 = opcode_5 != 4'h0 ? _GEN_5374 : _GEN_4994; // @[executor.scala 470:55]
  wire [7:0] _GEN_5763 = opcode_5 != 4'h0 ? _GEN_5375 : _GEN_4995; // @[executor.scala 470:55]
  wire [7:0] _GEN_5764 = opcode_5 != 4'h0 ? _GEN_5376 : _GEN_4996; // @[executor.scala 470:55]
  wire [7:0] _GEN_5765 = opcode_5 != 4'h0 ? _GEN_5377 : _GEN_4997; // @[executor.scala 470:55]
  wire [7:0] _GEN_5766 = opcode_5 != 4'h0 ? _GEN_5382 : _GEN_4998; // @[executor.scala 470:55]
  wire [7:0] _GEN_5767 = opcode_5 != 4'h0 ? _GEN_5383 : _GEN_4999; // @[executor.scala 470:55]
  wire [7:0] _GEN_5768 = opcode_5 != 4'h0 ? _GEN_5384 : _GEN_5000; // @[executor.scala 470:55]
  wire [7:0] _GEN_5769 = opcode_5 != 4'h0 ? _GEN_5385 : _GEN_5001; // @[executor.scala 470:55]
  wire [7:0] _GEN_5770 = opcode_5 != 4'h0 ? _GEN_5390 : _GEN_5002; // @[executor.scala 470:55]
  wire [7:0] _GEN_5771 = opcode_5 != 4'h0 ? _GEN_5391 : _GEN_5003; // @[executor.scala 470:55]
  wire [7:0] _GEN_5772 = opcode_5 != 4'h0 ? _GEN_5392 : _GEN_5004; // @[executor.scala 470:55]
  wire [7:0] _GEN_5773 = opcode_5 != 4'h0 ? _GEN_5393 : _GEN_5005; // @[executor.scala 470:55]
  wire [7:0] _GEN_5774 = opcode_5 != 4'h0 ? _GEN_5398 : _GEN_5006; // @[executor.scala 470:55]
  wire [7:0] _GEN_5775 = opcode_5 != 4'h0 ? _GEN_5399 : _GEN_5007; // @[executor.scala 470:55]
  wire [7:0] _GEN_5776 = opcode_5 != 4'h0 ? _GEN_5400 : _GEN_5008; // @[executor.scala 470:55]
  wire [7:0] _GEN_5777 = opcode_5 != 4'h0 ? _GEN_5401 : _GEN_5009; // @[executor.scala 470:55]
  wire [7:0] _GEN_5778 = opcode_5 != 4'h0 ? _GEN_5406 : _GEN_5010; // @[executor.scala 470:55]
  wire [7:0] _GEN_5779 = opcode_5 != 4'h0 ? _GEN_5407 : _GEN_5011; // @[executor.scala 470:55]
  wire [7:0] _GEN_5780 = opcode_5 != 4'h0 ? _GEN_5408 : _GEN_5012; // @[executor.scala 470:55]
  wire [7:0] _GEN_5781 = opcode_5 != 4'h0 ? _GEN_5409 : _GEN_5013; // @[executor.scala 470:55]
  wire [7:0] _GEN_5782 = opcode_5 != 4'h0 ? _GEN_5414 : _GEN_5014; // @[executor.scala 470:55]
  wire [7:0] _GEN_5783 = opcode_5 != 4'h0 ? _GEN_5415 : _GEN_5015; // @[executor.scala 470:55]
  wire [7:0] _GEN_5784 = opcode_5 != 4'h0 ? _GEN_5416 : _GEN_5016; // @[executor.scala 470:55]
  wire [7:0] _GEN_5785 = opcode_5 != 4'h0 ? _GEN_5417 : _GEN_5017; // @[executor.scala 470:55]
  wire [7:0] _GEN_5786 = opcode_5 != 4'h0 ? _GEN_5422 : _GEN_5018; // @[executor.scala 470:55]
  wire [7:0] _GEN_5787 = opcode_5 != 4'h0 ? _GEN_5423 : _GEN_5019; // @[executor.scala 470:55]
  wire [7:0] _GEN_5788 = opcode_5 != 4'h0 ? _GEN_5424 : _GEN_5020; // @[executor.scala 470:55]
  wire [7:0] _GEN_5789 = opcode_5 != 4'h0 ? _GEN_5425 : _GEN_5021; // @[executor.scala 470:55]
  wire [7:0] _GEN_5790 = opcode_5 != 4'h0 ? _GEN_5430 : _GEN_5022; // @[executor.scala 470:55]
  wire [7:0] _GEN_5791 = opcode_5 != 4'h0 ? _GEN_5431 : _GEN_5023; // @[executor.scala 470:55]
  wire [7:0] _GEN_5792 = opcode_5 != 4'h0 ? _GEN_5432 : _GEN_5024; // @[executor.scala 470:55]
  wire [7:0] _GEN_5793 = opcode_5 != 4'h0 ? _GEN_5433 : _GEN_5025; // @[executor.scala 470:55]
  wire [7:0] _GEN_5794 = opcode_5 != 4'h0 ? _GEN_5438 : _GEN_5026; // @[executor.scala 470:55]
  wire [7:0] _GEN_5795 = opcode_5 != 4'h0 ? _GEN_5439 : _GEN_5027; // @[executor.scala 470:55]
  wire [7:0] _GEN_5796 = opcode_5 != 4'h0 ? _GEN_5440 : _GEN_5028; // @[executor.scala 470:55]
  wire [7:0] _GEN_5797 = opcode_5 != 4'h0 ? _GEN_5441 : _GEN_5029; // @[executor.scala 470:55]
  wire [7:0] _GEN_5798 = opcode_5 != 4'h0 ? _GEN_5446 : _GEN_5030; // @[executor.scala 470:55]
  wire [7:0] _GEN_5799 = opcode_5 != 4'h0 ? _GEN_5447 : _GEN_5031; // @[executor.scala 470:55]
  wire [7:0] _GEN_5800 = opcode_5 != 4'h0 ? _GEN_5448 : _GEN_5032; // @[executor.scala 470:55]
  wire [7:0] _GEN_5801 = opcode_5 != 4'h0 ? _GEN_5449 : _GEN_5033; // @[executor.scala 470:55]
  wire [7:0] _GEN_5802 = opcode_5 != 4'h0 ? _GEN_5454 : _GEN_5034; // @[executor.scala 470:55]
  wire [7:0] _GEN_5803 = opcode_5 != 4'h0 ? _GEN_5455 : _GEN_5035; // @[executor.scala 470:55]
  wire [7:0] _GEN_5804 = opcode_5 != 4'h0 ? _GEN_5456 : _GEN_5036; // @[executor.scala 470:55]
  wire [7:0] _GEN_5805 = opcode_5 != 4'h0 ? _GEN_5457 : _GEN_5037; // @[executor.scala 470:55]
  wire [7:0] _GEN_5806 = opcode_5 != 4'h0 ? _GEN_5462 : _GEN_5038; // @[executor.scala 470:55]
  wire [7:0] _GEN_5807 = opcode_5 != 4'h0 ? _GEN_5463 : _GEN_5039; // @[executor.scala 470:55]
  wire [7:0] _GEN_5808 = opcode_5 != 4'h0 ? _GEN_5464 : _GEN_5040; // @[executor.scala 470:55]
  wire [7:0] _GEN_5809 = opcode_5 != 4'h0 ? _GEN_5465 : _GEN_5041; // @[executor.scala 470:55]
  wire [7:0] _GEN_5810 = opcode_5 != 4'h0 ? _GEN_5470 : _GEN_5042; // @[executor.scala 470:55]
  wire [7:0] _GEN_5811 = opcode_5 != 4'h0 ? _GEN_5471 : _GEN_5043; // @[executor.scala 470:55]
  wire [7:0] _GEN_5812 = opcode_5 != 4'h0 ? _GEN_5472 : _GEN_5044; // @[executor.scala 470:55]
  wire [7:0] _GEN_5813 = opcode_5 != 4'h0 ? _GEN_5473 : _GEN_5045; // @[executor.scala 470:55]
  wire [7:0] _GEN_5814 = opcode_5 != 4'h0 ? _GEN_5478 : _GEN_5046; // @[executor.scala 470:55]
  wire [7:0] _GEN_5815 = opcode_5 != 4'h0 ? _GEN_5479 : _GEN_5047; // @[executor.scala 470:55]
  wire [7:0] _GEN_5816 = opcode_5 != 4'h0 ? _GEN_5480 : _GEN_5048; // @[executor.scala 470:55]
  wire [7:0] _GEN_5817 = opcode_5 != 4'h0 ? _GEN_5481 : _GEN_5049; // @[executor.scala 470:55]
  wire [7:0] _GEN_5818 = opcode_5 != 4'h0 ? _GEN_5486 : _GEN_5050; // @[executor.scala 470:55]
  wire [7:0] _GEN_5819 = opcode_5 != 4'h0 ? _GEN_5487 : _GEN_5051; // @[executor.scala 470:55]
  wire [7:0] _GEN_5820 = opcode_5 != 4'h0 ? _GEN_5488 : _GEN_5052; // @[executor.scala 470:55]
  wire [7:0] _GEN_5821 = opcode_5 != 4'h0 ? _GEN_5489 : _GEN_5053; // @[executor.scala 470:55]
  wire [7:0] _GEN_5822 = opcode_5 != 4'h0 ? _GEN_5494 : _GEN_5054; // @[executor.scala 470:55]
  wire [7:0] _GEN_5823 = opcode_5 != 4'h0 ? _GEN_5495 : _GEN_5055; // @[executor.scala 470:55]
  wire [7:0] _GEN_5824 = opcode_5 != 4'h0 ? _GEN_5496 : _GEN_5056; // @[executor.scala 470:55]
  wire [7:0] _GEN_5825 = opcode_5 != 4'h0 ? _GEN_5497 : _GEN_5057; // @[executor.scala 470:55]
  wire [7:0] _GEN_5826 = opcode_5 != 4'h0 ? _GEN_5502 : _GEN_5058; // @[executor.scala 470:55]
  wire [7:0] _GEN_5827 = opcode_5 != 4'h0 ? _GEN_5503 : _GEN_5059; // @[executor.scala 470:55]
  wire [7:0] _GEN_5828 = opcode_5 != 4'h0 ? _GEN_5504 : _GEN_5060; // @[executor.scala 470:55]
  wire [7:0] _GEN_5829 = opcode_5 != 4'h0 ? _GEN_5505 : _GEN_5061; // @[executor.scala 470:55]
  wire [7:0] _GEN_5830 = opcode_5 != 4'h0 ? _GEN_5510 : _GEN_5062; // @[executor.scala 470:55]
  wire [7:0] _GEN_5831 = opcode_5 != 4'h0 ? _GEN_5511 : _GEN_5063; // @[executor.scala 470:55]
  wire [7:0] _GEN_5832 = opcode_5 != 4'h0 ? _GEN_5512 : _GEN_5064; // @[executor.scala 470:55]
  wire [7:0] _GEN_5833 = opcode_5 != 4'h0 ? _GEN_5513 : _GEN_5065; // @[executor.scala 470:55]
  wire [7:0] _GEN_5834 = opcode_5 != 4'h0 ? _GEN_5518 : _GEN_5066; // @[executor.scala 470:55]
  wire [7:0] _GEN_5835 = opcode_5 != 4'h0 ? _GEN_5519 : _GEN_5067; // @[executor.scala 470:55]
  wire [7:0] _GEN_5836 = opcode_5 != 4'h0 ? _GEN_5520 : _GEN_5068; // @[executor.scala 470:55]
  wire [7:0] _GEN_5837 = opcode_5 != 4'h0 ? _GEN_5521 : _GEN_5069; // @[executor.scala 470:55]
  wire [7:0] _GEN_5838 = opcode_5 != 4'h0 ? _GEN_5526 : _GEN_5070; // @[executor.scala 470:55]
  wire [7:0] _GEN_5839 = opcode_5 != 4'h0 ? _GEN_5527 : _GEN_5071; // @[executor.scala 470:55]
  wire [7:0] _GEN_5840 = opcode_5 != 4'h0 ? _GEN_5528 : _GEN_5072; // @[executor.scala 470:55]
  wire [7:0] _GEN_5841 = opcode_5 != 4'h0 ? _GEN_5529 : _GEN_5073; // @[executor.scala 470:55]
  wire [7:0] _GEN_5842 = opcode_5 != 4'h0 ? _GEN_5534 : _GEN_5074; // @[executor.scala 470:55]
  wire [7:0] _GEN_5843 = opcode_5 != 4'h0 ? _GEN_5535 : _GEN_5075; // @[executor.scala 470:55]
  wire [7:0] _GEN_5844 = opcode_5 != 4'h0 ? _GEN_5536 : _GEN_5076; // @[executor.scala 470:55]
  wire [7:0] _GEN_5845 = opcode_5 != 4'h0 ? _GEN_5537 : _GEN_5077; // @[executor.scala 470:55]
  wire [7:0] _GEN_5846 = opcode_5 != 4'h0 ? _GEN_5542 : _GEN_5078; // @[executor.scala 470:55]
  wire [7:0] _GEN_5847 = opcode_5 != 4'h0 ? _GEN_5543 : _GEN_5079; // @[executor.scala 470:55]
  wire [7:0] _GEN_5848 = opcode_5 != 4'h0 ? _GEN_5544 : _GEN_5080; // @[executor.scala 470:55]
  wire [7:0] _GEN_5849 = opcode_5 != 4'h0 ? _GEN_5545 : _GEN_5081; // @[executor.scala 470:55]
  wire [7:0] _GEN_5850 = opcode_5 != 4'h0 ? _GEN_5550 : _GEN_5082; // @[executor.scala 470:55]
  wire [7:0] _GEN_5851 = opcode_5 != 4'h0 ? _GEN_5551 : _GEN_5083; // @[executor.scala 470:55]
  wire [7:0] _GEN_5852 = opcode_5 != 4'h0 ? _GEN_5552 : _GEN_5084; // @[executor.scala 470:55]
  wire [7:0] _GEN_5853 = opcode_5 != 4'h0 ? _GEN_5553 : _GEN_5085; // @[executor.scala 470:55]
  wire [7:0] _GEN_5854 = opcode_5 != 4'h0 ? _GEN_5558 : _GEN_5086; // @[executor.scala 470:55]
  wire [7:0] _GEN_5855 = opcode_5 != 4'h0 ? _GEN_5559 : _GEN_5087; // @[executor.scala 470:55]
  wire [7:0] _GEN_5856 = opcode_5 != 4'h0 ? _GEN_5560 : _GEN_5088; // @[executor.scala 470:55]
  wire [7:0] _GEN_5857 = opcode_5 != 4'h0 ? _GEN_5561 : _GEN_5089; // @[executor.scala 470:55]
  wire [7:0] _GEN_5858 = opcode_5 != 4'h0 ? _GEN_5566 : _GEN_5090; // @[executor.scala 470:55]
  wire [7:0] _GEN_5859 = opcode_5 != 4'h0 ? _GEN_5567 : _GEN_5091; // @[executor.scala 470:55]
  wire [7:0] _GEN_5860 = opcode_5 != 4'h0 ? _GEN_5568 : _GEN_5092; // @[executor.scala 470:55]
  wire [7:0] _GEN_5861 = opcode_5 != 4'h0 ? _GEN_5569 : _GEN_5093; // @[executor.scala 470:55]
  wire [7:0] _GEN_5862 = opcode_5 != 4'h0 ? _GEN_5574 : _GEN_5094; // @[executor.scala 470:55]
  wire [7:0] _GEN_5863 = opcode_5 != 4'h0 ? _GEN_5575 : _GEN_5095; // @[executor.scala 470:55]
  wire [7:0] _GEN_5864 = opcode_5 != 4'h0 ? _GEN_5576 : _GEN_5096; // @[executor.scala 470:55]
  wire [7:0] _GEN_5865 = opcode_5 != 4'h0 ? _GEN_5577 : _GEN_5097; // @[executor.scala 470:55]
  wire [7:0] _GEN_5866 = opcode_5 != 4'h0 ? _GEN_5582 : _GEN_5098; // @[executor.scala 470:55]
  wire [7:0] _GEN_5867 = opcode_5 != 4'h0 ? _GEN_5583 : _GEN_5099; // @[executor.scala 470:55]
  wire [7:0] _GEN_5868 = opcode_5 != 4'h0 ? _GEN_5584 : _GEN_5100; // @[executor.scala 470:55]
  wire [7:0] _GEN_5869 = opcode_5 != 4'h0 ? _GEN_5585 : _GEN_5101; // @[executor.scala 470:55]
  wire [7:0] _GEN_5870 = opcode_5 != 4'h0 ? _GEN_5590 : _GEN_5102; // @[executor.scala 470:55]
  wire [7:0] _GEN_5871 = opcode_5 != 4'h0 ? _GEN_5591 : _GEN_5103; // @[executor.scala 470:55]
  wire [7:0] _GEN_5872 = opcode_5 != 4'h0 ? _GEN_5592 : _GEN_5104; // @[executor.scala 470:55]
  wire [7:0] _GEN_5873 = opcode_5 != 4'h0 ? _GEN_5593 : _GEN_5105; // @[executor.scala 470:55]
  wire [7:0] _GEN_5874 = opcode_5 != 4'h0 ? _GEN_5598 : _GEN_5106; // @[executor.scala 470:55]
  wire [7:0] _GEN_5875 = opcode_5 != 4'h0 ? _GEN_5599 : _GEN_5107; // @[executor.scala 470:55]
  wire [7:0] _GEN_5876 = opcode_5 != 4'h0 ? _GEN_5600 : _GEN_5108; // @[executor.scala 470:55]
  wire [7:0] _GEN_5877 = opcode_5 != 4'h0 ? _GEN_5601 : _GEN_5109; // @[executor.scala 470:55]
  wire [7:0] _GEN_5878 = opcode_5 != 4'h0 ? _GEN_5606 : _GEN_5110; // @[executor.scala 470:55]
  wire [7:0] _GEN_5879 = opcode_5 != 4'h0 ? _GEN_5607 : _GEN_5111; // @[executor.scala 470:55]
  wire [7:0] _GEN_5880 = opcode_5 != 4'h0 ? _GEN_5608 : _GEN_5112; // @[executor.scala 470:55]
  wire [7:0] _GEN_5881 = opcode_5 != 4'h0 ? _GEN_5609 : _GEN_5113; // @[executor.scala 470:55]
  wire [7:0] _GEN_5882 = opcode_5 != 4'h0 ? _GEN_5614 : _GEN_5114; // @[executor.scala 470:55]
  wire [7:0] _GEN_5883 = opcode_5 != 4'h0 ? _GEN_5615 : _GEN_5115; // @[executor.scala 470:55]
  wire [7:0] _GEN_5884 = opcode_5 != 4'h0 ? _GEN_5616 : _GEN_5116; // @[executor.scala 470:55]
  wire [7:0] _GEN_5885 = opcode_5 != 4'h0 ? _GEN_5617 : _GEN_5117; // @[executor.scala 470:55]
  wire [7:0] _GEN_5886 = opcode_5 != 4'h0 ? _GEN_5622 : _GEN_5118; // @[executor.scala 470:55]
  wire [7:0] _GEN_5887 = opcode_5 != 4'h0 ? _GEN_5623 : _GEN_5119; // @[executor.scala 470:55]
  wire [7:0] _GEN_5888 = opcode_5 != 4'h0 ? _GEN_5624 : _GEN_5120; // @[executor.scala 470:55]
  wire [7:0] _GEN_5889 = opcode_5 != 4'h0 ? _GEN_5625 : _GEN_5121; // @[executor.scala 470:55]
  wire [7:0] _GEN_5890 = opcode_5 != 4'h0 ? _GEN_5630 : _GEN_5122; // @[executor.scala 470:55]
  wire [7:0] _GEN_5891 = opcode_5 != 4'h0 ? _GEN_5631 : _GEN_5123; // @[executor.scala 470:55]
  wire [7:0] _GEN_5892 = opcode_5 != 4'h0 ? _GEN_5632 : _GEN_5124; // @[executor.scala 470:55]
  wire [7:0] _GEN_5893 = opcode_5 != 4'h0 ? _GEN_5633 : _GEN_5125; // @[executor.scala 470:55]
  wire [7:0] _GEN_5894 = opcode_5 != 4'h0 ? _GEN_5638 : _GEN_5126; // @[executor.scala 470:55]
  wire [7:0] _GEN_5895 = opcode_5 != 4'h0 ? _GEN_5639 : _GEN_5127; // @[executor.scala 470:55]
  wire [7:0] _GEN_5896 = opcode_5 != 4'h0 ? _GEN_5640 : _GEN_5128; // @[executor.scala 470:55]
  wire [7:0] _GEN_5897 = opcode_5 != 4'h0 ? _GEN_5641 : _GEN_5129; // @[executor.scala 470:55]
  wire [3:0] _GEN_5898 = opcode_5 == 4'hf ? parameter_2_5[13:10] : _GEN_4872; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_5899 = opcode_5 == 4'hf ? parameter_2_5[0] : _GEN_4873; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_5900 = opcode_5 == 4'hf ? _GEN_4874 : _GEN_5642; // @[executor.scala 466:52]
  wire [7:0] _GEN_5901 = opcode_5 == 4'hf ? _GEN_4875 : _GEN_5643; // @[executor.scala 466:52]
  wire [7:0] _GEN_5902 = opcode_5 == 4'hf ? _GEN_4876 : _GEN_5644; // @[executor.scala 466:52]
  wire [7:0] _GEN_5903 = opcode_5 == 4'hf ? _GEN_4877 : _GEN_5645; // @[executor.scala 466:52]
  wire [7:0] _GEN_5904 = opcode_5 == 4'hf ? _GEN_4878 : _GEN_5646; // @[executor.scala 466:52]
  wire [7:0] _GEN_5905 = opcode_5 == 4'hf ? _GEN_4879 : _GEN_5647; // @[executor.scala 466:52]
  wire [7:0] _GEN_5906 = opcode_5 == 4'hf ? _GEN_4880 : _GEN_5648; // @[executor.scala 466:52]
  wire [7:0] _GEN_5907 = opcode_5 == 4'hf ? _GEN_4881 : _GEN_5649; // @[executor.scala 466:52]
  wire [7:0] _GEN_5908 = opcode_5 == 4'hf ? _GEN_4882 : _GEN_5650; // @[executor.scala 466:52]
  wire [7:0] _GEN_5909 = opcode_5 == 4'hf ? _GEN_4883 : _GEN_5651; // @[executor.scala 466:52]
  wire [7:0] _GEN_5910 = opcode_5 == 4'hf ? _GEN_4884 : _GEN_5652; // @[executor.scala 466:52]
  wire [7:0] _GEN_5911 = opcode_5 == 4'hf ? _GEN_4885 : _GEN_5653; // @[executor.scala 466:52]
  wire [7:0] _GEN_5912 = opcode_5 == 4'hf ? _GEN_4886 : _GEN_5654; // @[executor.scala 466:52]
  wire [7:0] _GEN_5913 = opcode_5 == 4'hf ? _GEN_4887 : _GEN_5655; // @[executor.scala 466:52]
  wire [7:0] _GEN_5914 = opcode_5 == 4'hf ? _GEN_4888 : _GEN_5656; // @[executor.scala 466:52]
  wire [7:0] _GEN_5915 = opcode_5 == 4'hf ? _GEN_4889 : _GEN_5657; // @[executor.scala 466:52]
  wire [7:0] _GEN_5916 = opcode_5 == 4'hf ? _GEN_4890 : _GEN_5658; // @[executor.scala 466:52]
  wire [7:0] _GEN_5917 = opcode_5 == 4'hf ? _GEN_4891 : _GEN_5659; // @[executor.scala 466:52]
  wire [7:0] _GEN_5918 = opcode_5 == 4'hf ? _GEN_4892 : _GEN_5660; // @[executor.scala 466:52]
  wire [7:0] _GEN_5919 = opcode_5 == 4'hf ? _GEN_4893 : _GEN_5661; // @[executor.scala 466:52]
  wire [7:0] _GEN_5920 = opcode_5 == 4'hf ? _GEN_4894 : _GEN_5662; // @[executor.scala 466:52]
  wire [7:0] _GEN_5921 = opcode_5 == 4'hf ? _GEN_4895 : _GEN_5663; // @[executor.scala 466:52]
  wire [7:0] _GEN_5922 = opcode_5 == 4'hf ? _GEN_4896 : _GEN_5664; // @[executor.scala 466:52]
  wire [7:0] _GEN_5923 = opcode_5 == 4'hf ? _GEN_4897 : _GEN_5665; // @[executor.scala 466:52]
  wire [7:0] _GEN_5924 = opcode_5 == 4'hf ? _GEN_4898 : _GEN_5666; // @[executor.scala 466:52]
  wire [7:0] _GEN_5925 = opcode_5 == 4'hf ? _GEN_4899 : _GEN_5667; // @[executor.scala 466:52]
  wire [7:0] _GEN_5926 = opcode_5 == 4'hf ? _GEN_4900 : _GEN_5668; // @[executor.scala 466:52]
  wire [7:0] _GEN_5927 = opcode_5 == 4'hf ? _GEN_4901 : _GEN_5669; // @[executor.scala 466:52]
  wire [7:0] _GEN_5928 = opcode_5 == 4'hf ? _GEN_4902 : _GEN_5670; // @[executor.scala 466:52]
  wire [7:0] _GEN_5929 = opcode_5 == 4'hf ? _GEN_4903 : _GEN_5671; // @[executor.scala 466:52]
  wire [7:0] _GEN_5930 = opcode_5 == 4'hf ? _GEN_4904 : _GEN_5672; // @[executor.scala 466:52]
  wire [7:0] _GEN_5931 = opcode_5 == 4'hf ? _GEN_4905 : _GEN_5673; // @[executor.scala 466:52]
  wire [7:0] _GEN_5932 = opcode_5 == 4'hf ? _GEN_4906 : _GEN_5674; // @[executor.scala 466:52]
  wire [7:0] _GEN_5933 = opcode_5 == 4'hf ? _GEN_4907 : _GEN_5675; // @[executor.scala 466:52]
  wire [7:0] _GEN_5934 = opcode_5 == 4'hf ? _GEN_4908 : _GEN_5676; // @[executor.scala 466:52]
  wire [7:0] _GEN_5935 = opcode_5 == 4'hf ? _GEN_4909 : _GEN_5677; // @[executor.scala 466:52]
  wire [7:0] _GEN_5936 = opcode_5 == 4'hf ? _GEN_4910 : _GEN_5678; // @[executor.scala 466:52]
  wire [7:0] _GEN_5937 = opcode_5 == 4'hf ? _GEN_4911 : _GEN_5679; // @[executor.scala 466:52]
  wire [7:0] _GEN_5938 = opcode_5 == 4'hf ? _GEN_4912 : _GEN_5680; // @[executor.scala 466:52]
  wire [7:0] _GEN_5939 = opcode_5 == 4'hf ? _GEN_4913 : _GEN_5681; // @[executor.scala 466:52]
  wire [7:0] _GEN_5940 = opcode_5 == 4'hf ? _GEN_4914 : _GEN_5682; // @[executor.scala 466:52]
  wire [7:0] _GEN_5941 = opcode_5 == 4'hf ? _GEN_4915 : _GEN_5683; // @[executor.scala 466:52]
  wire [7:0] _GEN_5942 = opcode_5 == 4'hf ? _GEN_4916 : _GEN_5684; // @[executor.scala 466:52]
  wire [7:0] _GEN_5943 = opcode_5 == 4'hf ? _GEN_4917 : _GEN_5685; // @[executor.scala 466:52]
  wire [7:0] _GEN_5944 = opcode_5 == 4'hf ? _GEN_4918 : _GEN_5686; // @[executor.scala 466:52]
  wire [7:0] _GEN_5945 = opcode_5 == 4'hf ? _GEN_4919 : _GEN_5687; // @[executor.scala 466:52]
  wire [7:0] _GEN_5946 = opcode_5 == 4'hf ? _GEN_4920 : _GEN_5688; // @[executor.scala 466:52]
  wire [7:0] _GEN_5947 = opcode_5 == 4'hf ? _GEN_4921 : _GEN_5689; // @[executor.scala 466:52]
  wire [7:0] _GEN_5948 = opcode_5 == 4'hf ? _GEN_4922 : _GEN_5690; // @[executor.scala 466:52]
  wire [7:0] _GEN_5949 = opcode_5 == 4'hf ? _GEN_4923 : _GEN_5691; // @[executor.scala 466:52]
  wire [7:0] _GEN_5950 = opcode_5 == 4'hf ? _GEN_4924 : _GEN_5692; // @[executor.scala 466:52]
  wire [7:0] _GEN_5951 = opcode_5 == 4'hf ? _GEN_4925 : _GEN_5693; // @[executor.scala 466:52]
  wire [7:0] _GEN_5952 = opcode_5 == 4'hf ? _GEN_4926 : _GEN_5694; // @[executor.scala 466:52]
  wire [7:0] _GEN_5953 = opcode_5 == 4'hf ? _GEN_4927 : _GEN_5695; // @[executor.scala 466:52]
  wire [7:0] _GEN_5954 = opcode_5 == 4'hf ? _GEN_4928 : _GEN_5696; // @[executor.scala 466:52]
  wire [7:0] _GEN_5955 = opcode_5 == 4'hf ? _GEN_4929 : _GEN_5697; // @[executor.scala 466:52]
  wire [7:0] _GEN_5956 = opcode_5 == 4'hf ? _GEN_4930 : _GEN_5698; // @[executor.scala 466:52]
  wire [7:0] _GEN_5957 = opcode_5 == 4'hf ? _GEN_4931 : _GEN_5699; // @[executor.scala 466:52]
  wire [7:0] _GEN_5958 = opcode_5 == 4'hf ? _GEN_4932 : _GEN_5700; // @[executor.scala 466:52]
  wire [7:0] _GEN_5959 = opcode_5 == 4'hf ? _GEN_4933 : _GEN_5701; // @[executor.scala 466:52]
  wire [7:0] _GEN_5960 = opcode_5 == 4'hf ? _GEN_4934 : _GEN_5702; // @[executor.scala 466:52]
  wire [7:0] _GEN_5961 = opcode_5 == 4'hf ? _GEN_4935 : _GEN_5703; // @[executor.scala 466:52]
  wire [7:0] _GEN_5962 = opcode_5 == 4'hf ? _GEN_4936 : _GEN_5704; // @[executor.scala 466:52]
  wire [7:0] _GEN_5963 = opcode_5 == 4'hf ? _GEN_4937 : _GEN_5705; // @[executor.scala 466:52]
  wire [7:0] _GEN_5964 = opcode_5 == 4'hf ? _GEN_4938 : _GEN_5706; // @[executor.scala 466:52]
  wire [7:0] _GEN_5965 = opcode_5 == 4'hf ? _GEN_4939 : _GEN_5707; // @[executor.scala 466:52]
  wire [7:0] _GEN_5966 = opcode_5 == 4'hf ? _GEN_4940 : _GEN_5708; // @[executor.scala 466:52]
  wire [7:0] _GEN_5967 = opcode_5 == 4'hf ? _GEN_4941 : _GEN_5709; // @[executor.scala 466:52]
  wire [7:0] _GEN_5968 = opcode_5 == 4'hf ? _GEN_4942 : _GEN_5710; // @[executor.scala 466:52]
  wire [7:0] _GEN_5969 = opcode_5 == 4'hf ? _GEN_4943 : _GEN_5711; // @[executor.scala 466:52]
  wire [7:0] _GEN_5970 = opcode_5 == 4'hf ? _GEN_4944 : _GEN_5712; // @[executor.scala 466:52]
  wire [7:0] _GEN_5971 = opcode_5 == 4'hf ? _GEN_4945 : _GEN_5713; // @[executor.scala 466:52]
  wire [7:0] _GEN_5972 = opcode_5 == 4'hf ? _GEN_4946 : _GEN_5714; // @[executor.scala 466:52]
  wire [7:0] _GEN_5973 = opcode_5 == 4'hf ? _GEN_4947 : _GEN_5715; // @[executor.scala 466:52]
  wire [7:0] _GEN_5974 = opcode_5 == 4'hf ? _GEN_4948 : _GEN_5716; // @[executor.scala 466:52]
  wire [7:0] _GEN_5975 = opcode_5 == 4'hf ? _GEN_4949 : _GEN_5717; // @[executor.scala 466:52]
  wire [7:0] _GEN_5976 = opcode_5 == 4'hf ? _GEN_4950 : _GEN_5718; // @[executor.scala 466:52]
  wire [7:0] _GEN_5977 = opcode_5 == 4'hf ? _GEN_4951 : _GEN_5719; // @[executor.scala 466:52]
  wire [7:0] _GEN_5978 = opcode_5 == 4'hf ? _GEN_4952 : _GEN_5720; // @[executor.scala 466:52]
  wire [7:0] _GEN_5979 = opcode_5 == 4'hf ? _GEN_4953 : _GEN_5721; // @[executor.scala 466:52]
  wire [7:0] _GEN_5980 = opcode_5 == 4'hf ? _GEN_4954 : _GEN_5722; // @[executor.scala 466:52]
  wire [7:0] _GEN_5981 = opcode_5 == 4'hf ? _GEN_4955 : _GEN_5723; // @[executor.scala 466:52]
  wire [7:0] _GEN_5982 = opcode_5 == 4'hf ? _GEN_4956 : _GEN_5724; // @[executor.scala 466:52]
  wire [7:0] _GEN_5983 = opcode_5 == 4'hf ? _GEN_4957 : _GEN_5725; // @[executor.scala 466:52]
  wire [7:0] _GEN_5984 = opcode_5 == 4'hf ? _GEN_4958 : _GEN_5726; // @[executor.scala 466:52]
  wire [7:0] _GEN_5985 = opcode_5 == 4'hf ? _GEN_4959 : _GEN_5727; // @[executor.scala 466:52]
  wire [7:0] _GEN_5986 = opcode_5 == 4'hf ? _GEN_4960 : _GEN_5728; // @[executor.scala 466:52]
  wire [7:0] _GEN_5987 = opcode_5 == 4'hf ? _GEN_4961 : _GEN_5729; // @[executor.scala 466:52]
  wire [7:0] _GEN_5988 = opcode_5 == 4'hf ? _GEN_4962 : _GEN_5730; // @[executor.scala 466:52]
  wire [7:0] _GEN_5989 = opcode_5 == 4'hf ? _GEN_4963 : _GEN_5731; // @[executor.scala 466:52]
  wire [7:0] _GEN_5990 = opcode_5 == 4'hf ? _GEN_4964 : _GEN_5732; // @[executor.scala 466:52]
  wire [7:0] _GEN_5991 = opcode_5 == 4'hf ? _GEN_4965 : _GEN_5733; // @[executor.scala 466:52]
  wire [7:0] _GEN_5992 = opcode_5 == 4'hf ? _GEN_4966 : _GEN_5734; // @[executor.scala 466:52]
  wire [7:0] _GEN_5993 = opcode_5 == 4'hf ? _GEN_4967 : _GEN_5735; // @[executor.scala 466:52]
  wire [7:0] _GEN_5994 = opcode_5 == 4'hf ? _GEN_4968 : _GEN_5736; // @[executor.scala 466:52]
  wire [7:0] _GEN_5995 = opcode_5 == 4'hf ? _GEN_4969 : _GEN_5737; // @[executor.scala 466:52]
  wire [7:0] _GEN_5996 = opcode_5 == 4'hf ? _GEN_4970 : _GEN_5738; // @[executor.scala 466:52]
  wire [7:0] _GEN_5997 = opcode_5 == 4'hf ? _GEN_4971 : _GEN_5739; // @[executor.scala 466:52]
  wire [7:0] _GEN_5998 = opcode_5 == 4'hf ? _GEN_4972 : _GEN_5740; // @[executor.scala 466:52]
  wire [7:0] _GEN_5999 = opcode_5 == 4'hf ? _GEN_4973 : _GEN_5741; // @[executor.scala 466:52]
  wire [7:0] _GEN_6000 = opcode_5 == 4'hf ? _GEN_4974 : _GEN_5742; // @[executor.scala 466:52]
  wire [7:0] _GEN_6001 = opcode_5 == 4'hf ? _GEN_4975 : _GEN_5743; // @[executor.scala 466:52]
  wire [7:0] _GEN_6002 = opcode_5 == 4'hf ? _GEN_4976 : _GEN_5744; // @[executor.scala 466:52]
  wire [7:0] _GEN_6003 = opcode_5 == 4'hf ? _GEN_4977 : _GEN_5745; // @[executor.scala 466:52]
  wire [7:0] _GEN_6004 = opcode_5 == 4'hf ? _GEN_4978 : _GEN_5746; // @[executor.scala 466:52]
  wire [7:0] _GEN_6005 = opcode_5 == 4'hf ? _GEN_4979 : _GEN_5747; // @[executor.scala 466:52]
  wire [7:0] _GEN_6006 = opcode_5 == 4'hf ? _GEN_4980 : _GEN_5748; // @[executor.scala 466:52]
  wire [7:0] _GEN_6007 = opcode_5 == 4'hf ? _GEN_4981 : _GEN_5749; // @[executor.scala 466:52]
  wire [7:0] _GEN_6008 = opcode_5 == 4'hf ? _GEN_4982 : _GEN_5750; // @[executor.scala 466:52]
  wire [7:0] _GEN_6009 = opcode_5 == 4'hf ? _GEN_4983 : _GEN_5751; // @[executor.scala 466:52]
  wire [7:0] _GEN_6010 = opcode_5 == 4'hf ? _GEN_4984 : _GEN_5752; // @[executor.scala 466:52]
  wire [7:0] _GEN_6011 = opcode_5 == 4'hf ? _GEN_4985 : _GEN_5753; // @[executor.scala 466:52]
  wire [7:0] _GEN_6012 = opcode_5 == 4'hf ? _GEN_4986 : _GEN_5754; // @[executor.scala 466:52]
  wire [7:0] _GEN_6013 = opcode_5 == 4'hf ? _GEN_4987 : _GEN_5755; // @[executor.scala 466:52]
  wire [7:0] _GEN_6014 = opcode_5 == 4'hf ? _GEN_4988 : _GEN_5756; // @[executor.scala 466:52]
  wire [7:0] _GEN_6015 = opcode_5 == 4'hf ? _GEN_4989 : _GEN_5757; // @[executor.scala 466:52]
  wire [7:0] _GEN_6016 = opcode_5 == 4'hf ? _GEN_4990 : _GEN_5758; // @[executor.scala 466:52]
  wire [7:0] _GEN_6017 = opcode_5 == 4'hf ? _GEN_4991 : _GEN_5759; // @[executor.scala 466:52]
  wire [7:0] _GEN_6018 = opcode_5 == 4'hf ? _GEN_4992 : _GEN_5760; // @[executor.scala 466:52]
  wire [7:0] _GEN_6019 = opcode_5 == 4'hf ? _GEN_4993 : _GEN_5761; // @[executor.scala 466:52]
  wire [7:0] _GEN_6020 = opcode_5 == 4'hf ? _GEN_4994 : _GEN_5762; // @[executor.scala 466:52]
  wire [7:0] _GEN_6021 = opcode_5 == 4'hf ? _GEN_4995 : _GEN_5763; // @[executor.scala 466:52]
  wire [7:0] _GEN_6022 = opcode_5 == 4'hf ? _GEN_4996 : _GEN_5764; // @[executor.scala 466:52]
  wire [7:0] _GEN_6023 = opcode_5 == 4'hf ? _GEN_4997 : _GEN_5765; // @[executor.scala 466:52]
  wire [7:0] _GEN_6024 = opcode_5 == 4'hf ? _GEN_4998 : _GEN_5766; // @[executor.scala 466:52]
  wire [7:0] _GEN_6025 = opcode_5 == 4'hf ? _GEN_4999 : _GEN_5767; // @[executor.scala 466:52]
  wire [7:0] _GEN_6026 = opcode_5 == 4'hf ? _GEN_5000 : _GEN_5768; // @[executor.scala 466:52]
  wire [7:0] _GEN_6027 = opcode_5 == 4'hf ? _GEN_5001 : _GEN_5769; // @[executor.scala 466:52]
  wire [7:0] _GEN_6028 = opcode_5 == 4'hf ? _GEN_5002 : _GEN_5770; // @[executor.scala 466:52]
  wire [7:0] _GEN_6029 = opcode_5 == 4'hf ? _GEN_5003 : _GEN_5771; // @[executor.scala 466:52]
  wire [7:0] _GEN_6030 = opcode_5 == 4'hf ? _GEN_5004 : _GEN_5772; // @[executor.scala 466:52]
  wire [7:0] _GEN_6031 = opcode_5 == 4'hf ? _GEN_5005 : _GEN_5773; // @[executor.scala 466:52]
  wire [7:0] _GEN_6032 = opcode_5 == 4'hf ? _GEN_5006 : _GEN_5774; // @[executor.scala 466:52]
  wire [7:0] _GEN_6033 = opcode_5 == 4'hf ? _GEN_5007 : _GEN_5775; // @[executor.scala 466:52]
  wire [7:0] _GEN_6034 = opcode_5 == 4'hf ? _GEN_5008 : _GEN_5776; // @[executor.scala 466:52]
  wire [7:0] _GEN_6035 = opcode_5 == 4'hf ? _GEN_5009 : _GEN_5777; // @[executor.scala 466:52]
  wire [7:0] _GEN_6036 = opcode_5 == 4'hf ? _GEN_5010 : _GEN_5778; // @[executor.scala 466:52]
  wire [7:0] _GEN_6037 = opcode_5 == 4'hf ? _GEN_5011 : _GEN_5779; // @[executor.scala 466:52]
  wire [7:0] _GEN_6038 = opcode_5 == 4'hf ? _GEN_5012 : _GEN_5780; // @[executor.scala 466:52]
  wire [7:0] _GEN_6039 = opcode_5 == 4'hf ? _GEN_5013 : _GEN_5781; // @[executor.scala 466:52]
  wire [7:0] _GEN_6040 = opcode_5 == 4'hf ? _GEN_5014 : _GEN_5782; // @[executor.scala 466:52]
  wire [7:0] _GEN_6041 = opcode_5 == 4'hf ? _GEN_5015 : _GEN_5783; // @[executor.scala 466:52]
  wire [7:0] _GEN_6042 = opcode_5 == 4'hf ? _GEN_5016 : _GEN_5784; // @[executor.scala 466:52]
  wire [7:0] _GEN_6043 = opcode_5 == 4'hf ? _GEN_5017 : _GEN_5785; // @[executor.scala 466:52]
  wire [7:0] _GEN_6044 = opcode_5 == 4'hf ? _GEN_5018 : _GEN_5786; // @[executor.scala 466:52]
  wire [7:0] _GEN_6045 = opcode_5 == 4'hf ? _GEN_5019 : _GEN_5787; // @[executor.scala 466:52]
  wire [7:0] _GEN_6046 = opcode_5 == 4'hf ? _GEN_5020 : _GEN_5788; // @[executor.scala 466:52]
  wire [7:0] _GEN_6047 = opcode_5 == 4'hf ? _GEN_5021 : _GEN_5789; // @[executor.scala 466:52]
  wire [7:0] _GEN_6048 = opcode_5 == 4'hf ? _GEN_5022 : _GEN_5790; // @[executor.scala 466:52]
  wire [7:0] _GEN_6049 = opcode_5 == 4'hf ? _GEN_5023 : _GEN_5791; // @[executor.scala 466:52]
  wire [7:0] _GEN_6050 = opcode_5 == 4'hf ? _GEN_5024 : _GEN_5792; // @[executor.scala 466:52]
  wire [7:0] _GEN_6051 = opcode_5 == 4'hf ? _GEN_5025 : _GEN_5793; // @[executor.scala 466:52]
  wire [7:0] _GEN_6052 = opcode_5 == 4'hf ? _GEN_5026 : _GEN_5794; // @[executor.scala 466:52]
  wire [7:0] _GEN_6053 = opcode_5 == 4'hf ? _GEN_5027 : _GEN_5795; // @[executor.scala 466:52]
  wire [7:0] _GEN_6054 = opcode_5 == 4'hf ? _GEN_5028 : _GEN_5796; // @[executor.scala 466:52]
  wire [7:0] _GEN_6055 = opcode_5 == 4'hf ? _GEN_5029 : _GEN_5797; // @[executor.scala 466:52]
  wire [7:0] _GEN_6056 = opcode_5 == 4'hf ? _GEN_5030 : _GEN_5798; // @[executor.scala 466:52]
  wire [7:0] _GEN_6057 = opcode_5 == 4'hf ? _GEN_5031 : _GEN_5799; // @[executor.scala 466:52]
  wire [7:0] _GEN_6058 = opcode_5 == 4'hf ? _GEN_5032 : _GEN_5800; // @[executor.scala 466:52]
  wire [7:0] _GEN_6059 = opcode_5 == 4'hf ? _GEN_5033 : _GEN_5801; // @[executor.scala 466:52]
  wire [7:0] _GEN_6060 = opcode_5 == 4'hf ? _GEN_5034 : _GEN_5802; // @[executor.scala 466:52]
  wire [7:0] _GEN_6061 = opcode_5 == 4'hf ? _GEN_5035 : _GEN_5803; // @[executor.scala 466:52]
  wire [7:0] _GEN_6062 = opcode_5 == 4'hf ? _GEN_5036 : _GEN_5804; // @[executor.scala 466:52]
  wire [7:0] _GEN_6063 = opcode_5 == 4'hf ? _GEN_5037 : _GEN_5805; // @[executor.scala 466:52]
  wire [7:0] _GEN_6064 = opcode_5 == 4'hf ? _GEN_5038 : _GEN_5806; // @[executor.scala 466:52]
  wire [7:0] _GEN_6065 = opcode_5 == 4'hf ? _GEN_5039 : _GEN_5807; // @[executor.scala 466:52]
  wire [7:0] _GEN_6066 = opcode_5 == 4'hf ? _GEN_5040 : _GEN_5808; // @[executor.scala 466:52]
  wire [7:0] _GEN_6067 = opcode_5 == 4'hf ? _GEN_5041 : _GEN_5809; // @[executor.scala 466:52]
  wire [7:0] _GEN_6068 = opcode_5 == 4'hf ? _GEN_5042 : _GEN_5810; // @[executor.scala 466:52]
  wire [7:0] _GEN_6069 = opcode_5 == 4'hf ? _GEN_5043 : _GEN_5811; // @[executor.scala 466:52]
  wire [7:0] _GEN_6070 = opcode_5 == 4'hf ? _GEN_5044 : _GEN_5812; // @[executor.scala 466:52]
  wire [7:0] _GEN_6071 = opcode_5 == 4'hf ? _GEN_5045 : _GEN_5813; // @[executor.scala 466:52]
  wire [7:0] _GEN_6072 = opcode_5 == 4'hf ? _GEN_5046 : _GEN_5814; // @[executor.scala 466:52]
  wire [7:0] _GEN_6073 = opcode_5 == 4'hf ? _GEN_5047 : _GEN_5815; // @[executor.scala 466:52]
  wire [7:0] _GEN_6074 = opcode_5 == 4'hf ? _GEN_5048 : _GEN_5816; // @[executor.scala 466:52]
  wire [7:0] _GEN_6075 = opcode_5 == 4'hf ? _GEN_5049 : _GEN_5817; // @[executor.scala 466:52]
  wire [7:0] _GEN_6076 = opcode_5 == 4'hf ? _GEN_5050 : _GEN_5818; // @[executor.scala 466:52]
  wire [7:0] _GEN_6077 = opcode_5 == 4'hf ? _GEN_5051 : _GEN_5819; // @[executor.scala 466:52]
  wire [7:0] _GEN_6078 = opcode_5 == 4'hf ? _GEN_5052 : _GEN_5820; // @[executor.scala 466:52]
  wire [7:0] _GEN_6079 = opcode_5 == 4'hf ? _GEN_5053 : _GEN_5821; // @[executor.scala 466:52]
  wire [7:0] _GEN_6080 = opcode_5 == 4'hf ? _GEN_5054 : _GEN_5822; // @[executor.scala 466:52]
  wire [7:0] _GEN_6081 = opcode_5 == 4'hf ? _GEN_5055 : _GEN_5823; // @[executor.scala 466:52]
  wire [7:0] _GEN_6082 = opcode_5 == 4'hf ? _GEN_5056 : _GEN_5824; // @[executor.scala 466:52]
  wire [7:0] _GEN_6083 = opcode_5 == 4'hf ? _GEN_5057 : _GEN_5825; // @[executor.scala 466:52]
  wire [7:0] _GEN_6084 = opcode_5 == 4'hf ? _GEN_5058 : _GEN_5826; // @[executor.scala 466:52]
  wire [7:0] _GEN_6085 = opcode_5 == 4'hf ? _GEN_5059 : _GEN_5827; // @[executor.scala 466:52]
  wire [7:0] _GEN_6086 = opcode_5 == 4'hf ? _GEN_5060 : _GEN_5828; // @[executor.scala 466:52]
  wire [7:0] _GEN_6087 = opcode_5 == 4'hf ? _GEN_5061 : _GEN_5829; // @[executor.scala 466:52]
  wire [7:0] _GEN_6088 = opcode_5 == 4'hf ? _GEN_5062 : _GEN_5830; // @[executor.scala 466:52]
  wire [7:0] _GEN_6089 = opcode_5 == 4'hf ? _GEN_5063 : _GEN_5831; // @[executor.scala 466:52]
  wire [7:0] _GEN_6090 = opcode_5 == 4'hf ? _GEN_5064 : _GEN_5832; // @[executor.scala 466:52]
  wire [7:0] _GEN_6091 = opcode_5 == 4'hf ? _GEN_5065 : _GEN_5833; // @[executor.scala 466:52]
  wire [7:0] _GEN_6092 = opcode_5 == 4'hf ? _GEN_5066 : _GEN_5834; // @[executor.scala 466:52]
  wire [7:0] _GEN_6093 = opcode_5 == 4'hf ? _GEN_5067 : _GEN_5835; // @[executor.scala 466:52]
  wire [7:0] _GEN_6094 = opcode_5 == 4'hf ? _GEN_5068 : _GEN_5836; // @[executor.scala 466:52]
  wire [7:0] _GEN_6095 = opcode_5 == 4'hf ? _GEN_5069 : _GEN_5837; // @[executor.scala 466:52]
  wire [7:0] _GEN_6096 = opcode_5 == 4'hf ? _GEN_5070 : _GEN_5838; // @[executor.scala 466:52]
  wire [7:0] _GEN_6097 = opcode_5 == 4'hf ? _GEN_5071 : _GEN_5839; // @[executor.scala 466:52]
  wire [7:0] _GEN_6098 = opcode_5 == 4'hf ? _GEN_5072 : _GEN_5840; // @[executor.scala 466:52]
  wire [7:0] _GEN_6099 = opcode_5 == 4'hf ? _GEN_5073 : _GEN_5841; // @[executor.scala 466:52]
  wire [7:0] _GEN_6100 = opcode_5 == 4'hf ? _GEN_5074 : _GEN_5842; // @[executor.scala 466:52]
  wire [7:0] _GEN_6101 = opcode_5 == 4'hf ? _GEN_5075 : _GEN_5843; // @[executor.scala 466:52]
  wire [7:0] _GEN_6102 = opcode_5 == 4'hf ? _GEN_5076 : _GEN_5844; // @[executor.scala 466:52]
  wire [7:0] _GEN_6103 = opcode_5 == 4'hf ? _GEN_5077 : _GEN_5845; // @[executor.scala 466:52]
  wire [7:0] _GEN_6104 = opcode_5 == 4'hf ? _GEN_5078 : _GEN_5846; // @[executor.scala 466:52]
  wire [7:0] _GEN_6105 = opcode_5 == 4'hf ? _GEN_5079 : _GEN_5847; // @[executor.scala 466:52]
  wire [7:0] _GEN_6106 = opcode_5 == 4'hf ? _GEN_5080 : _GEN_5848; // @[executor.scala 466:52]
  wire [7:0] _GEN_6107 = opcode_5 == 4'hf ? _GEN_5081 : _GEN_5849; // @[executor.scala 466:52]
  wire [7:0] _GEN_6108 = opcode_5 == 4'hf ? _GEN_5082 : _GEN_5850; // @[executor.scala 466:52]
  wire [7:0] _GEN_6109 = opcode_5 == 4'hf ? _GEN_5083 : _GEN_5851; // @[executor.scala 466:52]
  wire [7:0] _GEN_6110 = opcode_5 == 4'hf ? _GEN_5084 : _GEN_5852; // @[executor.scala 466:52]
  wire [7:0] _GEN_6111 = opcode_5 == 4'hf ? _GEN_5085 : _GEN_5853; // @[executor.scala 466:52]
  wire [7:0] _GEN_6112 = opcode_5 == 4'hf ? _GEN_5086 : _GEN_5854; // @[executor.scala 466:52]
  wire [7:0] _GEN_6113 = opcode_5 == 4'hf ? _GEN_5087 : _GEN_5855; // @[executor.scala 466:52]
  wire [7:0] _GEN_6114 = opcode_5 == 4'hf ? _GEN_5088 : _GEN_5856; // @[executor.scala 466:52]
  wire [7:0] _GEN_6115 = opcode_5 == 4'hf ? _GEN_5089 : _GEN_5857; // @[executor.scala 466:52]
  wire [7:0] _GEN_6116 = opcode_5 == 4'hf ? _GEN_5090 : _GEN_5858; // @[executor.scala 466:52]
  wire [7:0] _GEN_6117 = opcode_5 == 4'hf ? _GEN_5091 : _GEN_5859; // @[executor.scala 466:52]
  wire [7:0] _GEN_6118 = opcode_5 == 4'hf ? _GEN_5092 : _GEN_5860; // @[executor.scala 466:52]
  wire [7:0] _GEN_6119 = opcode_5 == 4'hf ? _GEN_5093 : _GEN_5861; // @[executor.scala 466:52]
  wire [7:0] _GEN_6120 = opcode_5 == 4'hf ? _GEN_5094 : _GEN_5862; // @[executor.scala 466:52]
  wire [7:0] _GEN_6121 = opcode_5 == 4'hf ? _GEN_5095 : _GEN_5863; // @[executor.scala 466:52]
  wire [7:0] _GEN_6122 = opcode_5 == 4'hf ? _GEN_5096 : _GEN_5864; // @[executor.scala 466:52]
  wire [7:0] _GEN_6123 = opcode_5 == 4'hf ? _GEN_5097 : _GEN_5865; // @[executor.scala 466:52]
  wire [7:0] _GEN_6124 = opcode_5 == 4'hf ? _GEN_5098 : _GEN_5866; // @[executor.scala 466:52]
  wire [7:0] _GEN_6125 = opcode_5 == 4'hf ? _GEN_5099 : _GEN_5867; // @[executor.scala 466:52]
  wire [7:0] _GEN_6126 = opcode_5 == 4'hf ? _GEN_5100 : _GEN_5868; // @[executor.scala 466:52]
  wire [7:0] _GEN_6127 = opcode_5 == 4'hf ? _GEN_5101 : _GEN_5869; // @[executor.scala 466:52]
  wire [7:0] _GEN_6128 = opcode_5 == 4'hf ? _GEN_5102 : _GEN_5870; // @[executor.scala 466:52]
  wire [7:0] _GEN_6129 = opcode_5 == 4'hf ? _GEN_5103 : _GEN_5871; // @[executor.scala 466:52]
  wire [7:0] _GEN_6130 = opcode_5 == 4'hf ? _GEN_5104 : _GEN_5872; // @[executor.scala 466:52]
  wire [7:0] _GEN_6131 = opcode_5 == 4'hf ? _GEN_5105 : _GEN_5873; // @[executor.scala 466:52]
  wire [7:0] _GEN_6132 = opcode_5 == 4'hf ? _GEN_5106 : _GEN_5874; // @[executor.scala 466:52]
  wire [7:0] _GEN_6133 = opcode_5 == 4'hf ? _GEN_5107 : _GEN_5875; // @[executor.scala 466:52]
  wire [7:0] _GEN_6134 = opcode_5 == 4'hf ? _GEN_5108 : _GEN_5876; // @[executor.scala 466:52]
  wire [7:0] _GEN_6135 = opcode_5 == 4'hf ? _GEN_5109 : _GEN_5877; // @[executor.scala 466:52]
  wire [7:0] _GEN_6136 = opcode_5 == 4'hf ? _GEN_5110 : _GEN_5878; // @[executor.scala 466:52]
  wire [7:0] _GEN_6137 = opcode_5 == 4'hf ? _GEN_5111 : _GEN_5879; // @[executor.scala 466:52]
  wire [7:0] _GEN_6138 = opcode_5 == 4'hf ? _GEN_5112 : _GEN_5880; // @[executor.scala 466:52]
  wire [7:0] _GEN_6139 = opcode_5 == 4'hf ? _GEN_5113 : _GEN_5881; // @[executor.scala 466:52]
  wire [7:0] _GEN_6140 = opcode_5 == 4'hf ? _GEN_5114 : _GEN_5882; // @[executor.scala 466:52]
  wire [7:0] _GEN_6141 = opcode_5 == 4'hf ? _GEN_5115 : _GEN_5883; // @[executor.scala 466:52]
  wire [7:0] _GEN_6142 = opcode_5 == 4'hf ? _GEN_5116 : _GEN_5884; // @[executor.scala 466:52]
  wire [7:0] _GEN_6143 = opcode_5 == 4'hf ? _GEN_5117 : _GEN_5885; // @[executor.scala 466:52]
  wire [7:0] _GEN_6144 = opcode_5 == 4'hf ? _GEN_5118 : _GEN_5886; // @[executor.scala 466:52]
  wire [7:0] _GEN_6145 = opcode_5 == 4'hf ? _GEN_5119 : _GEN_5887; // @[executor.scala 466:52]
  wire [7:0] _GEN_6146 = opcode_5 == 4'hf ? _GEN_5120 : _GEN_5888; // @[executor.scala 466:52]
  wire [7:0] _GEN_6147 = opcode_5 == 4'hf ? _GEN_5121 : _GEN_5889; // @[executor.scala 466:52]
  wire [7:0] _GEN_6148 = opcode_5 == 4'hf ? _GEN_5122 : _GEN_5890; // @[executor.scala 466:52]
  wire [7:0] _GEN_6149 = opcode_5 == 4'hf ? _GEN_5123 : _GEN_5891; // @[executor.scala 466:52]
  wire [7:0] _GEN_6150 = opcode_5 == 4'hf ? _GEN_5124 : _GEN_5892; // @[executor.scala 466:52]
  wire [7:0] _GEN_6151 = opcode_5 == 4'hf ? _GEN_5125 : _GEN_5893; // @[executor.scala 466:52]
  wire [7:0] _GEN_6152 = opcode_5 == 4'hf ? _GEN_5126 : _GEN_5894; // @[executor.scala 466:52]
  wire [7:0] _GEN_6153 = opcode_5 == 4'hf ? _GEN_5127 : _GEN_5895; // @[executor.scala 466:52]
  wire [7:0] _GEN_6154 = opcode_5 == 4'hf ? _GEN_5128 : _GEN_5896; // @[executor.scala 466:52]
  wire [7:0] _GEN_6155 = opcode_5 == 4'hf ? _GEN_5129 : _GEN_5897; // @[executor.scala 466:52]
  wire [3:0] opcode_6 = vliw_6[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_6 = vliw_6[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8850 = {{2'd0}, dst_offset_6}; // @[executor.scala 473:49]
  wire [7:0] byte_1536 = field_6[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6156 = mask_6[0] ? byte_1536 : _GEN_5900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1537 = field_6[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6157 = mask_6[1] ? byte_1537 : _GEN_5901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1538 = field_6[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6158 = mask_6[2] ? byte_1538 : _GEN_5902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1539 = field_6[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6159 = mask_6[3] ? byte_1539 : _GEN_5903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6160 = _GEN_8850 == 8'h0 ? _GEN_6156 : _GEN_5900; // @[executor.scala 473:84]
  wire [7:0] _GEN_6161 = _GEN_8850 == 8'h0 ? _GEN_6157 : _GEN_5901; // @[executor.scala 473:84]
  wire [7:0] _GEN_6162 = _GEN_8850 == 8'h0 ? _GEN_6158 : _GEN_5902; // @[executor.scala 473:84]
  wire [7:0] _GEN_6163 = _GEN_8850 == 8'h0 ? _GEN_6159 : _GEN_5903; // @[executor.scala 473:84]
  wire [7:0] _GEN_6164 = mask_6[0] ? byte_1536 : _GEN_5904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6165 = mask_6[1] ? byte_1537 : _GEN_5905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6166 = mask_6[2] ? byte_1538 : _GEN_5906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6167 = mask_6[3] ? byte_1539 : _GEN_5907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6168 = _GEN_8850 == 8'h1 ? _GEN_6164 : _GEN_5904; // @[executor.scala 473:84]
  wire [7:0] _GEN_6169 = _GEN_8850 == 8'h1 ? _GEN_6165 : _GEN_5905; // @[executor.scala 473:84]
  wire [7:0] _GEN_6170 = _GEN_8850 == 8'h1 ? _GEN_6166 : _GEN_5906; // @[executor.scala 473:84]
  wire [7:0] _GEN_6171 = _GEN_8850 == 8'h1 ? _GEN_6167 : _GEN_5907; // @[executor.scala 473:84]
  wire [7:0] _GEN_6172 = mask_6[0] ? byte_1536 : _GEN_5908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6173 = mask_6[1] ? byte_1537 : _GEN_5909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6174 = mask_6[2] ? byte_1538 : _GEN_5910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6175 = mask_6[3] ? byte_1539 : _GEN_5911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6176 = _GEN_8850 == 8'h2 ? _GEN_6172 : _GEN_5908; // @[executor.scala 473:84]
  wire [7:0] _GEN_6177 = _GEN_8850 == 8'h2 ? _GEN_6173 : _GEN_5909; // @[executor.scala 473:84]
  wire [7:0] _GEN_6178 = _GEN_8850 == 8'h2 ? _GEN_6174 : _GEN_5910; // @[executor.scala 473:84]
  wire [7:0] _GEN_6179 = _GEN_8850 == 8'h2 ? _GEN_6175 : _GEN_5911; // @[executor.scala 473:84]
  wire [7:0] _GEN_6180 = mask_6[0] ? byte_1536 : _GEN_5912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6181 = mask_6[1] ? byte_1537 : _GEN_5913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6182 = mask_6[2] ? byte_1538 : _GEN_5914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6183 = mask_6[3] ? byte_1539 : _GEN_5915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6184 = _GEN_8850 == 8'h3 ? _GEN_6180 : _GEN_5912; // @[executor.scala 473:84]
  wire [7:0] _GEN_6185 = _GEN_8850 == 8'h3 ? _GEN_6181 : _GEN_5913; // @[executor.scala 473:84]
  wire [7:0] _GEN_6186 = _GEN_8850 == 8'h3 ? _GEN_6182 : _GEN_5914; // @[executor.scala 473:84]
  wire [7:0] _GEN_6187 = _GEN_8850 == 8'h3 ? _GEN_6183 : _GEN_5915; // @[executor.scala 473:84]
  wire [7:0] _GEN_6188 = mask_6[0] ? byte_1536 : _GEN_5916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6189 = mask_6[1] ? byte_1537 : _GEN_5917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6190 = mask_6[2] ? byte_1538 : _GEN_5918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6191 = mask_6[3] ? byte_1539 : _GEN_5919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6192 = _GEN_8850 == 8'h4 ? _GEN_6188 : _GEN_5916; // @[executor.scala 473:84]
  wire [7:0] _GEN_6193 = _GEN_8850 == 8'h4 ? _GEN_6189 : _GEN_5917; // @[executor.scala 473:84]
  wire [7:0] _GEN_6194 = _GEN_8850 == 8'h4 ? _GEN_6190 : _GEN_5918; // @[executor.scala 473:84]
  wire [7:0] _GEN_6195 = _GEN_8850 == 8'h4 ? _GEN_6191 : _GEN_5919; // @[executor.scala 473:84]
  wire [7:0] _GEN_6196 = mask_6[0] ? byte_1536 : _GEN_5920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6197 = mask_6[1] ? byte_1537 : _GEN_5921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6198 = mask_6[2] ? byte_1538 : _GEN_5922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6199 = mask_6[3] ? byte_1539 : _GEN_5923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6200 = _GEN_8850 == 8'h5 ? _GEN_6196 : _GEN_5920; // @[executor.scala 473:84]
  wire [7:0] _GEN_6201 = _GEN_8850 == 8'h5 ? _GEN_6197 : _GEN_5921; // @[executor.scala 473:84]
  wire [7:0] _GEN_6202 = _GEN_8850 == 8'h5 ? _GEN_6198 : _GEN_5922; // @[executor.scala 473:84]
  wire [7:0] _GEN_6203 = _GEN_8850 == 8'h5 ? _GEN_6199 : _GEN_5923; // @[executor.scala 473:84]
  wire [7:0] _GEN_6204 = mask_6[0] ? byte_1536 : _GEN_5924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6205 = mask_6[1] ? byte_1537 : _GEN_5925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6206 = mask_6[2] ? byte_1538 : _GEN_5926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6207 = mask_6[3] ? byte_1539 : _GEN_5927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6208 = _GEN_8850 == 8'h6 ? _GEN_6204 : _GEN_5924; // @[executor.scala 473:84]
  wire [7:0] _GEN_6209 = _GEN_8850 == 8'h6 ? _GEN_6205 : _GEN_5925; // @[executor.scala 473:84]
  wire [7:0] _GEN_6210 = _GEN_8850 == 8'h6 ? _GEN_6206 : _GEN_5926; // @[executor.scala 473:84]
  wire [7:0] _GEN_6211 = _GEN_8850 == 8'h6 ? _GEN_6207 : _GEN_5927; // @[executor.scala 473:84]
  wire [7:0] _GEN_6212 = mask_6[0] ? byte_1536 : _GEN_5928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6213 = mask_6[1] ? byte_1537 : _GEN_5929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6214 = mask_6[2] ? byte_1538 : _GEN_5930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6215 = mask_6[3] ? byte_1539 : _GEN_5931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6216 = _GEN_8850 == 8'h7 ? _GEN_6212 : _GEN_5928; // @[executor.scala 473:84]
  wire [7:0] _GEN_6217 = _GEN_8850 == 8'h7 ? _GEN_6213 : _GEN_5929; // @[executor.scala 473:84]
  wire [7:0] _GEN_6218 = _GEN_8850 == 8'h7 ? _GEN_6214 : _GEN_5930; // @[executor.scala 473:84]
  wire [7:0] _GEN_6219 = _GEN_8850 == 8'h7 ? _GEN_6215 : _GEN_5931; // @[executor.scala 473:84]
  wire [7:0] _GEN_6220 = mask_6[0] ? byte_1536 : _GEN_5932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6221 = mask_6[1] ? byte_1537 : _GEN_5933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6222 = mask_6[2] ? byte_1538 : _GEN_5934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6223 = mask_6[3] ? byte_1539 : _GEN_5935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6224 = _GEN_8850 == 8'h8 ? _GEN_6220 : _GEN_5932; // @[executor.scala 473:84]
  wire [7:0] _GEN_6225 = _GEN_8850 == 8'h8 ? _GEN_6221 : _GEN_5933; // @[executor.scala 473:84]
  wire [7:0] _GEN_6226 = _GEN_8850 == 8'h8 ? _GEN_6222 : _GEN_5934; // @[executor.scala 473:84]
  wire [7:0] _GEN_6227 = _GEN_8850 == 8'h8 ? _GEN_6223 : _GEN_5935; // @[executor.scala 473:84]
  wire [7:0] _GEN_6228 = mask_6[0] ? byte_1536 : _GEN_5936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6229 = mask_6[1] ? byte_1537 : _GEN_5937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6230 = mask_6[2] ? byte_1538 : _GEN_5938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6231 = mask_6[3] ? byte_1539 : _GEN_5939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6232 = _GEN_8850 == 8'h9 ? _GEN_6228 : _GEN_5936; // @[executor.scala 473:84]
  wire [7:0] _GEN_6233 = _GEN_8850 == 8'h9 ? _GEN_6229 : _GEN_5937; // @[executor.scala 473:84]
  wire [7:0] _GEN_6234 = _GEN_8850 == 8'h9 ? _GEN_6230 : _GEN_5938; // @[executor.scala 473:84]
  wire [7:0] _GEN_6235 = _GEN_8850 == 8'h9 ? _GEN_6231 : _GEN_5939; // @[executor.scala 473:84]
  wire [7:0] _GEN_6236 = mask_6[0] ? byte_1536 : _GEN_5940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6237 = mask_6[1] ? byte_1537 : _GEN_5941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6238 = mask_6[2] ? byte_1538 : _GEN_5942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6239 = mask_6[3] ? byte_1539 : _GEN_5943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6240 = _GEN_8850 == 8'ha ? _GEN_6236 : _GEN_5940; // @[executor.scala 473:84]
  wire [7:0] _GEN_6241 = _GEN_8850 == 8'ha ? _GEN_6237 : _GEN_5941; // @[executor.scala 473:84]
  wire [7:0] _GEN_6242 = _GEN_8850 == 8'ha ? _GEN_6238 : _GEN_5942; // @[executor.scala 473:84]
  wire [7:0] _GEN_6243 = _GEN_8850 == 8'ha ? _GEN_6239 : _GEN_5943; // @[executor.scala 473:84]
  wire [7:0] _GEN_6244 = mask_6[0] ? byte_1536 : _GEN_5944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6245 = mask_6[1] ? byte_1537 : _GEN_5945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6246 = mask_6[2] ? byte_1538 : _GEN_5946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6247 = mask_6[3] ? byte_1539 : _GEN_5947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6248 = _GEN_8850 == 8'hb ? _GEN_6244 : _GEN_5944; // @[executor.scala 473:84]
  wire [7:0] _GEN_6249 = _GEN_8850 == 8'hb ? _GEN_6245 : _GEN_5945; // @[executor.scala 473:84]
  wire [7:0] _GEN_6250 = _GEN_8850 == 8'hb ? _GEN_6246 : _GEN_5946; // @[executor.scala 473:84]
  wire [7:0] _GEN_6251 = _GEN_8850 == 8'hb ? _GEN_6247 : _GEN_5947; // @[executor.scala 473:84]
  wire [7:0] _GEN_6252 = mask_6[0] ? byte_1536 : _GEN_5948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6253 = mask_6[1] ? byte_1537 : _GEN_5949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6254 = mask_6[2] ? byte_1538 : _GEN_5950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6255 = mask_6[3] ? byte_1539 : _GEN_5951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6256 = _GEN_8850 == 8'hc ? _GEN_6252 : _GEN_5948; // @[executor.scala 473:84]
  wire [7:0] _GEN_6257 = _GEN_8850 == 8'hc ? _GEN_6253 : _GEN_5949; // @[executor.scala 473:84]
  wire [7:0] _GEN_6258 = _GEN_8850 == 8'hc ? _GEN_6254 : _GEN_5950; // @[executor.scala 473:84]
  wire [7:0] _GEN_6259 = _GEN_8850 == 8'hc ? _GEN_6255 : _GEN_5951; // @[executor.scala 473:84]
  wire [7:0] _GEN_6260 = mask_6[0] ? byte_1536 : _GEN_5952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6261 = mask_6[1] ? byte_1537 : _GEN_5953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6262 = mask_6[2] ? byte_1538 : _GEN_5954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6263 = mask_6[3] ? byte_1539 : _GEN_5955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6264 = _GEN_8850 == 8'hd ? _GEN_6260 : _GEN_5952; // @[executor.scala 473:84]
  wire [7:0] _GEN_6265 = _GEN_8850 == 8'hd ? _GEN_6261 : _GEN_5953; // @[executor.scala 473:84]
  wire [7:0] _GEN_6266 = _GEN_8850 == 8'hd ? _GEN_6262 : _GEN_5954; // @[executor.scala 473:84]
  wire [7:0] _GEN_6267 = _GEN_8850 == 8'hd ? _GEN_6263 : _GEN_5955; // @[executor.scala 473:84]
  wire [7:0] _GEN_6268 = mask_6[0] ? byte_1536 : _GEN_5956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6269 = mask_6[1] ? byte_1537 : _GEN_5957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6270 = mask_6[2] ? byte_1538 : _GEN_5958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6271 = mask_6[3] ? byte_1539 : _GEN_5959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6272 = _GEN_8850 == 8'he ? _GEN_6268 : _GEN_5956; // @[executor.scala 473:84]
  wire [7:0] _GEN_6273 = _GEN_8850 == 8'he ? _GEN_6269 : _GEN_5957; // @[executor.scala 473:84]
  wire [7:0] _GEN_6274 = _GEN_8850 == 8'he ? _GEN_6270 : _GEN_5958; // @[executor.scala 473:84]
  wire [7:0] _GEN_6275 = _GEN_8850 == 8'he ? _GEN_6271 : _GEN_5959; // @[executor.scala 473:84]
  wire [7:0] _GEN_6276 = mask_6[0] ? byte_1536 : _GEN_5960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6277 = mask_6[1] ? byte_1537 : _GEN_5961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6278 = mask_6[2] ? byte_1538 : _GEN_5962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6279 = mask_6[3] ? byte_1539 : _GEN_5963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6280 = _GEN_8850 == 8'hf ? _GEN_6276 : _GEN_5960; // @[executor.scala 473:84]
  wire [7:0] _GEN_6281 = _GEN_8850 == 8'hf ? _GEN_6277 : _GEN_5961; // @[executor.scala 473:84]
  wire [7:0] _GEN_6282 = _GEN_8850 == 8'hf ? _GEN_6278 : _GEN_5962; // @[executor.scala 473:84]
  wire [7:0] _GEN_6283 = _GEN_8850 == 8'hf ? _GEN_6279 : _GEN_5963; // @[executor.scala 473:84]
  wire [7:0] _GEN_6284 = mask_6[0] ? byte_1536 : _GEN_5964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6285 = mask_6[1] ? byte_1537 : _GEN_5965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6286 = mask_6[2] ? byte_1538 : _GEN_5966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6287 = mask_6[3] ? byte_1539 : _GEN_5967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6288 = _GEN_8850 == 8'h10 ? _GEN_6284 : _GEN_5964; // @[executor.scala 473:84]
  wire [7:0] _GEN_6289 = _GEN_8850 == 8'h10 ? _GEN_6285 : _GEN_5965; // @[executor.scala 473:84]
  wire [7:0] _GEN_6290 = _GEN_8850 == 8'h10 ? _GEN_6286 : _GEN_5966; // @[executor.scala 473:84]
  wire [7:0] _GEN_6291 = _GEN_8850 == 8'h10 ? _GEN_6287 : _GEN_5967; // @[executor.scala 473:84]
  wire [7:0] _GEN_6292 = mask_6[0] ? byte_1536 : _GEN_5968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6293 = mask_6[1] ? byte_1537 : _GEN_5969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6294 = mask_6[2] ? byte_1538 : _GEN_5970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6295 = mask_6[3] ? byte_1539 : _GEN_5971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6296 = _GEN_8850 == 8'h11 ? _GEN_6292 : _GEN_5968; // @[executor.scala 473:84]
  wire [7:0] _GEN_6297 = _GEN_8850 == 8'h11 ? _GEN_6293 : _GEN_5969; // @[executor.scala 473:84]
  wire [7:0] _GEN_6298 = _GEN_8850 == 8'h11 ? _GEN_6294 : _GEN_5970; // @[executor.scala 473:84]
  wire [7:0] _GEN_6299 = _GEN_8850 == 8'h11 ? _GEN_6295 : _GEN_5971; // @[executor.scala 473:84]
  wire [7:0] _GEN_6300 = mask_6[0] ? byte_1536 : _GEN_5972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6301 = mask_6[1] ? byte_1537 : _GEN_5973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6302 = mask_6[2] ? byte_1538 : _GEN_5974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6303 = mask_6[3] ? byte_1539 : _GEN_5975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6304 = _GEN_8850 == 8'h12 ? _GEN_6300 : _GEN_5972; // @[executor.scala 473:84]
  wire [7:0] _GEN_6305 = _GEN_8850 == 8'h12 ? _GEN_6301 : _GEN_5973; // @[executor.scala 473:84]
  wire [7:0] _GEN_6306 = _GEN_8850 == 8'h12 ? _GEN_6302 : _GEN_5974; // @[executor.scala 473:84]
  wire [7:0] _GEN_6307 = _GEN_8850 == 8'h12 ? _GEN_6303 : _GEN_5975; // @[executor.scala 473:84]
  wire [7:0] _GEN_6308 = mask_6[0] ? byte_1536 : _GEN_5976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6309 = mask_6[1] ? byte_1537 : _GEN_5977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6310 = mask_6[2] ? byte_1538 : _GEN_5978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6311 = mask_6[3] ? byte_1539 : _GEN_5979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6312 = _GEN_8850 == 8'h13 ? _GEN_6308 : _GEN_5976; // @[executor.scala 473:84]
  wire [7:0] _GEN_6313 = _GEN_8850 == 8'h13 ? _GEN_6309 : _GEN_5977; // @[executor.scala 473:84]
  wire [7:0] _GEN_6314 = _GEN_8850 == 8'h13 ? _GEN_6310 : _GEN_5978; // @[executor.scala 473:84]
  wire [7:0] _GEN_6315 = _GEN_8850 == 8'h13 ? _GEN_6311 : _GEN_5979; // @[executor.scala 473:84]
  wire [7:0] _GEN_6316 = mask_6[0] ? byte_1536 : _GEN_5980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6317 = mask_6[1] ? byte_1537 : _GEN_5981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6318 = mask_6[2] ? byte_1538 : _GEN_5982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6319 = mask_6[3] ? byte_1539 : _GEN_5983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6320 = _GEN_8850 == 8'h14 ? _GEN_6316 : _GEN_5980; // @[executor.scala 473:84]
  wire [7:0] _GEN_6321 = _GEN_8850 == 8'h14 ? _GEN_6317 : _GEN_5981; // @[executor.scala 473:84]
  wire [7:0] _GEN_6322 = _GEN_8850 == 8'h14 ? _GEN_6318 : _GEN_5982; // @[executor.scala 473:84]
  wire [7:0] _GEN_6323 = _GEN_8850 == 8'h14 ? _GEN_6319 : _GEN_5983; // @[executor.scala 473:84]
  wire [7:0] _GEN_6324 = mask_6[0] ? byte_1536 : _GEN_5984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6325 = mask_6[1] ? byte_1537 : _GEN_5985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6326 = mask_6[2] ? byte_1538 : _GEN_5986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6327 = mask_6[3] ? byte_1539 : _GEN_5987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6328 = _GEN_8850 == 8'h15 ? _GEN_6324 : _GEN_5984; // @[executor.scala 473:84]
  wire [7:0] _GEN_6329 = _GEN_8850 == 8'h15 ? _GEN_6325 : _GEN_5985; // @[executor.scala 473:84]
  wire [7:0] _GEN_6330 = _GEN_8850 == 8'h15 ? _GEN_6326 : _GEN_5986; // @[executor.scala 473:84]
  wire [7:0] _GEN_6331 = _GEN_8850 == 8'h15 ? _GEN_6327 : _GEN_5987; // @[executor.scala 473:84]
  wire [7:0] _GEN_6332 = mask_6[0] ? byte_1536 : _GEN_5988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6333 = mask_6[1] ? byte_1537 : _GEN_5989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6334 = mask_6[2] ? byte_1538 : _GEN_5990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6335 = mask_6[3] ? byte_1539 : _GEN_5991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6336 = _GEN_8850 == 8'h16 ? _GEN_6332 : _GEN_5988; // @[executor.scala 473:84]
  wire [7:0] _GEN_6337 = _GEN_8850 == 8'h16 ? _GEN_6333 : _GEN_5989; // @[executor.scala 473:84]
  wire [7:0] _GEN_6338 = _GEN_8850 == 8'h16 ? _GEN_6334 : _GEN_5990; // @[executor.scala 473:84]
  wire [7:0] _GEN_6339 = _GEN_8850 == 8'h16 ? _GEN_6335 : _GEN_5991; // @[executor.scala 473:84]
  wire [7:0] _GEN_6340 = mask_6[0] ? byte_1536 : _GEN_5992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6341 = mask_6[1] ? byte_1537 : _GEN_5993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6342 = mask_6[2] ? byte_1538 : _GEN_5994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6343 = mask_6[3] ? byte_1539 : _GEN_5995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6344 = _GEN_8850 == 8'h17 ? _GEN_6340 : _GEN_5992; // @[executor.scala 473:84]
  wire [7:0] _GEN_6345 = _GEN_8850 == 8'h17 ? _GEN_6341 : _GEN_5993; // @[executor.scala 473:84]
  wire [7:0] _GEN_6346 = _GEN_8850 == 8'h17 ? _GEN_6342 : _GEN_5994; // @[executor.scala 473:84]
  wire [7:0] _GEN_6347 = _GEN_8850 == 8'h17 ? _GEN_6343 : _GEN_5995; // @[executor.scala 473:84]
  wire [7:0] _GEN_6348 = mask_6[0] ? byte_1536 : _GEN_5996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6349 = mask_6[1] ? byte_1537 : _GEN_5997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6350 = mask_6[2] ? byte_1538 : _GEN_5998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6351 = mask_6[3] ? byte_1539 : _GEN_5999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6352 = _GEN_8850 == 8'h18 ? _GEN_6348 : _GEN_5996; // @[executor.scala 473:84]
  wire [7:0] _GEN_6353 = _GEN_8850 == 8'h18 ? _GEN_6349 : _GEN_5997; // @[executor.scala 473:84]
  wire [7:0] _GEN_6354 = _GEN_8850 == 8'h18 ? _GEN_6350 : _GEN_5998; // @[executor.scala 473:84]
  wire [7:0] _GEN_6355 = _GEN_8850 == 8'h18 ? _GEN_6351 : _GEN_5999; // @[executor.scala 473:84]
  wire [7:0] _GEN_6356 = mask_6[0] ? byte_1536 : _GEN_6000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6357 = mask_6[1] ? byte_1537 : _GEN_6001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6358 = mask_6[2] ? byte_1538 : _GEN_6002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6359 = mask_6[3] ? byte_1539 : _GEN_6003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6360 = _GEN_8850 == 8'h19 ? _GEN_6356 : _GEN_6000; // @[executor.scala 473:84]
  wire [7:0] _GEN_6361 = _GEN_8850 == 8'h19 ? _GEN_6357 : _GEN_6001; // @[executor.scala 473:84]
  wire [7:0] _GEN_6362 = _GEN_8850 == 8'h19 ? _GEN_6358 : _GEN_6002; // @[executor.scala 473:84]
  wire [7:0] _GEN_6363 = _GEN_8850 == 8'h19 ? _GEN_6359 : _GEN_6003; // @[executor.scala 473:84]
  wire [7:0] _GEN_6364 = mask_6[0] ? byte_1536 : _GEN_6004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6365 = mask_6[1] ? byte_1537 : _GEN_6005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6366 = mask_6[2] ? byte_1538 : _GEN_6006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6367 = mask_6[3] ? byte_1539 : _GEN_6007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6368 = _GEN_8850 == 8'h1a ? _GEN_6364 : _GEN_6004; // @[executor.scala 473:84]
  wire [7:0] _GEN_6369 = _GEN_8850 == 8'h1a ? _GEN_6365 : _GEN_6005; // @[executor.scala 473:84]
  wire [7:0] _GEN_6370 = _GEN_8850 == 8'h1a ? _GEN_6366 : _GEN_6006; // @[executor.scala 473:84]
  wire [7:0] _GEN_6371 = _GEN_8850 == 8'h1a ? _GEN_6367 : _GEN_6007; // @[executor.scala 473:84]
  wire [7:0] _GEN_6372 = mask_6[0] ? byte_1536 : _GEN_6008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6373 = mask_6[1] ? byte_1537 : _GEN_6009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6374 = mask_6[2] ? byte_1538 : _GEN_6010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6375 = mask_6[3] ? byte_1539 : _GEN_6011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6376 = _GEN_8850 == 8'h1b ? _GEN_6372 : _GEN_6008; // @[executor.scala 473:84]
  wire [7:0] _GEN_6377 = _GEN_8850 == 8'h1b ? _GEN_6373 : _GEN_6009; // @[executor.scala 473:84]
  wire [7:0] _GEN_6378 = _GEN_8850 == 8'h1b ? _GEN_6374 : _GEN_6010; // @[executor.scala 473:84]
  wire [7:0] _GEN_6379 = _GEN_8850 == 8'h1b ? _GEN_6375 : _GEN_6011; // @[executor.scala 473:84]
  wire [7:0] _GEN_6380 = mask_6[0] ? byte_1536 : _GEN_6012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6381 = mask_6[1] ? byte_1537 : _GEN_6013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6382 = mask_6[2] ? byte_1538 : _GEN_6014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6383 = mask_6[3] ? byte_1539 : _GEN_6015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6384 = _GEN_8850 == 8'h1c ? _GEN_6380 : _GEN_6012; // @[executor.scala 473:84]
  wire [7:0] _GEN_6385 = _GEN_8850 == 8'h1c ? _GEN_6381 : _GEN_6013; // @[executor.scala 473:84]
  wire [7:0] _GEN_6386 = _GEN_8850 == 8'h1c ? _GEN_6382 : _GEN_6014; // @[executor.scala 473:84]
  wire [7:0] _GEN_6387 = _GEN_8850 == 8'h1c ? _GEN_6383 : _GEN_6015; // @[executor.scala 473:84]
  wire [7:0] _GEN_6388 = mask_6[0] ? byte_1536 : _GEN_6016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6389 = mask_6[1] ? byte_1537 : _GEN_6017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6390 = mask_6[2] ? byte_1538 : _GEN_6018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6391 = mask_6[3] ? byte_1539 : _GEN_6019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6392 = _GEN_8850 == 8'h1d ? _GEN_6388 : _GEN_6016; // @[executor.scala 473:84]
  wire [7:0] _GEN_6393 = _GEN_8850 == 8'h1d ? _GEN_6389 : _GEN_6017; // @[executor.scala 473:84]
  wire [7:0] _GEN_6394 = _GEN_8850 == 8'h1d ? _GEN_6390 : _GEN_6018; // @[executor.scala 473:84]
  wire [7:0] _GEN_6395 = _GEN_8850 == 8'h1d ? _GEN_6391 : _GEN_6019; // @[executor.scala 473:84]
  wire [7:0] _GEN_6396 = mask_6[0] ? byte_1536 : _GEN_6020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6397 = mask_6[1] ? byte_1537 : _GEN_6021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6398 = mask_6[2] ? byte_1538 : _GEN_6022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6399 = mask_6[3] ? byte_1539 : _GEN_6023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6400 = _GEN_8850 == 8'h1e ? _GEN_6396 : _GEN_6020; // @[executor.scala 473:84]
  wire [7:0] _GEN_6401 = _GEN_8850 == 8'h1e ? _GEN_6397 : _GEN_6021; // @[executor.scala 473:84]
  wire [7:0] _GEN_6402 = _GEN_8850 == 8'h1e ? _GEN_6398 : _GEN_6022; // @[executor.scala 473:84]
  wire [7:0] _GEN_6403 = _GEN_8850 == 8'h1e ? _GEN_6399 : _GEN_6023; // @[executor.scala 473:84]
  wire [7:0] _GEN_6404 = mask_6[0] ? byte_1536 : _GEN_6024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6405 = mask_6[1] ? byte_1537 : _GEN_6025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6406 = mask_6[2] ? byte_1538 : _GEN_6026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6407 = mask_6[3] ? byte_1539 : _GEN_6027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6408 = _GEN_8850 == 8'h1f ? _GEN_6404 : _GEN_6024; // @[executor.scala 473:84]
  wire [7:0] _GEN_6409 = _GEN_8850 == 8'h1f ? _GEN_6405 : _GEN_6025; // @[executor.scala 473:84]
  wire [7:0] _GEN_6410 = _GEN_8850 == 8'h1f ? _GEN_6406 : _GEN_6026; // @[executor.scala 473:84]
  wire [7:0] _GEN_6411 = _GEN_8850 == 8'h1f ? _GEN_6407 : _GEN_6027; // @[executor.scala 473:84]
  wire [7:0] _GEN_6412 = mask_6[0] ? byte_1536 : _GEN_6028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6413 = mask_6[1] ? byte_1537 : _GEN_6029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6414 = mask_6[2] ? byte_1538 : _GEN_6030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6415 = mask_6[3] ? byte_1539 : _GEN_6031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6416 = _GEN_8850 == 8'h20 ? _GEN_6412 : _GEN_6028; // @[executor.scala 473:84]
  wire [7:0] _GEN_6417 = _GEN_8850 == 8'h20 ? _GEN_6413 : _GEN_6029; // @[executor.scala 473:84]
  wire [7:0] _GEN_6418 = _GEN_8850 == 8'h20 ? _GEN_6414 : _GEN_6030; // @[executor.scala 473:84]
  wire [7:0] _GEN_6419 = _GEN_8850 == 8'h20 ? _GEN_6415 : _GEN_6031; // @[executor.scala 473:84]
  wire [7:0] _GEN_6420 = mask_6[0] ? byte_1536 : _GEN_6032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6421 = mask_6[1] ? byte_1537 : _GEN_6033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6422 = mask_6[2] ? byte_1538 : _GEN_6034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6423 = mask_6[3] ? byte_1539 : _GEN_6035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6424 = _GEN_8850 == 8'h21 ? _GEN_6420 : _GEN_6032; // @[executor.scala 473:84]
  wire [7:0] _GEN_6425 = _GEN_8850 == 8'h21 ? _GEN_6421 : _GEN_6033; // @[executor.scala 473:84]
  wire [7:0] _GEN_6426 = _GEN_8850 == 8'h21 ? _GEN_6422 : _GEN_6034; // @[executor.scala 473:84]
  wire [7:0] _GEN_6427 = _GEN_8850 == 8'h21 ? _GEN_6423 : _GEN_6035; // @[executor.scala 473:84]
  wire [7:0] _GEN_6428 = mask_6[0] ? byte_1536 : _GEN_6036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6429 = mask_6[1] ? byte_1537 : _GEN_6037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6430 = mask_6[2] ? byte_1538 : _GEN_6038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6431 = mask_6[3] ? byte_1539 : _GEN_6039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6432 = _GEN_8850 == 8'h22 ? _GEN_6428 : _GEN_6036; // @[executor.scala 473:84]
  wire [7:0] _GEN_6433 = _GEN_8850 == 8'h22 ? _GEN_6429 : _GEN_6037; // @[executor.scala 473:84]
  wire [7:0] _GEN_6434 = _GEN_8850 == 8'h22 ? _GEN_6430 : _GEN_6038; // @[executor.scala 473:84]
  wire [7:0] _GEN_6435 = _GEN_8850 == 8'h22 ? _GEN_6431 : _GEN_6039; // @[executor.scala 473:84]
  wire [7:0] _GEN_6436 = mask_6[0] ? byte_1536 : _GEN_6040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6437 = mask_6[1] ? byte_1537 : _GEN_6041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6438 = mask_6[2] ? byte_1538 : _GEN_6042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6439 = mask_6[3] ? byte_1539 : _GEN_6043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6440 = _GEN_8850 == 8'h23 ? _GEN_6436 : _GEN_6040; // @[executor.scala 473:84]
  wire [7:0] _GEN_6441 = _GEN_8850 == 8'h23 ? _GEN_6437 : _GEN_6041; // @[executor.scala 473:84]
  wire [7:0] _GEN_6442 = _GEN_8850 == 8'h23 ? _GEN_6438 : _GEN_6042; // @[executor.scala 473:84]
  wire [7:0] _GEN_6443 = _GEN_8850 == 8'h23 ? _GEN_6439 : _GEN_6043; // @[executor.scala 473:84]
  wire [7:0] _GEN_6444 = mask_6[0] ? byte_1536 : _GEN_6044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6445 = mask_6[1] ? byte_1537 : _GEN_6045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6446 = mask_6[2] ? byte_1538 : _GEN_6046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6447 = mask_6[3] ? byte_1539 : _GEN_6047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6448 = _GEN_8850 == 8'h24 ? _GEN_6444 : _GEN_6044; // @[executor.scala 473:84]
  wire [7:0] _GEN_6449 = _GEN_8850 == 8'h24 ? _GEN_6445 : _GEN_6045; // @[executor.scala 473:84]
  wire [7:0] _GEN_6450 = _GEN_8850 == 8'h24 ? _GEN_6446 : _GEN_6046; // @[executor.scala 473:84]
  wire [7:0] _GEN_6451 = _GEN_8850 == 8'h24 ? _GEN_6447 : _GEN_6047; // @[executor.scala 473:84]
  wire [7:0] _GEN_6452 = mask_6[0] ? byte_1536 : _GEN_6048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6453 = mask_6[1] ? byte_1537 : _GEN_6049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6454 = mask_6[2] ? byte_1538 : _GEN_6050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6455 = mask_6[3] ? byte_1539 : _GEN_6051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6456 = _GEN_8850 == 8'h25 ? _GEN_6452 : _GEN_6048; // @[executor.scala 473:84]
  wire [7:0] _GEN_6457 = _GEN_8850 == 8'h25 ? _GEN_6453 : _GEN_6049; // @[executor.scala 473:84]
  wire [7:0] _GEN_6458 = _GEN_8850 == 8'h25 ? _GEN_6454 : _GEN_6050; // @[executor.scala 473:84]
  wire [7:0] _GEN_6459 = _GEN_8850 == 8'h25 ? _GEN_6455 : _GEN_6051; // @[executor.scala 473:84]
  wire [7:0] _GEN_6460 = mask_6[0] ? byte_1536 : _GEN_6052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6461 = mask_6[1] ? byte_1537 : _GEN_6053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6462 = mask_6[2] ? byte_1538 : _GEN_6054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6463 = mask_6[3] ? byte_1539 : _GEN_6055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6464 = _GEN_8850 == 8'h26 ? _GEN_6460 : _GEN_6052; // @[executor.scala 473:84]
  wire [7:0] _GEN_6465 = _GEN_8850 == 8'h26 ? _GEN_6461 : _GEN_6053; // @[executor.scala 473:84]
  wire [7:0] _GEN_6466 = _GEN_8850 == 8'h26 ? _GEN_6462 : _GEN_6054; // @[executor.scala 473:84]
  wire [7:0] _GEN_6467 = _GEN_8850 == 8'h26 ? _GEN_6463 : _GEN_6055; // @[executor.scala 473:84]
  wire [7:0] _GEN_6468 = mask_6[0] ? byte_1536 : _GEN_6056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6469 = mask_6[1] ? byte_1537 : _GEN_6057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6470 = mask_6[2] ? byte_1538 : _GEN_6058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6471 = mask_6[3] ? byte_1539 : _GEN_6059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6472 = _GEN_8850 == 8'h27 ? _GEN_6468 : _GEN_6056; // @[executor.scala 473:84]
  wire [7:0] _GEN_6473 = _GEN_8850 == 8'h27 ? _GEN_6469 : _GEN_6057; // @[executor.scala 473:84]
  wire [7:0] _GEN_6474 = _GEN_8850 == 8'h27 ? _GEN_6470 : _GEN_6058; // @[executor.scala 473:84]
  wire [7:0] _GEN_6475 = _GEN_8850 == 8'h27 ? _GEN_6471 : _GEN_6059; // @[executor.scala 473:84]
  wire [7:0] _GEN_6476 = mask_6[0] ? byte_1536 : _GEN_6060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6477 = mask_6[1] ? byte_1537 : _GEN_6061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6478 = mask_6[2] ? byte_1538 : _GEN_6062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6479 = mask_6[3] ? byte_1539 : _GEN_6063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6480 = _GEN_8850 == 8'h28 ? _GEN_6476 : _GEN_6060; // @[executor.scala 473:84]
  wire [7:0] _GEN_6481 = _GEN_8850 == 8'h28 ? _GEN_6477 : _GEN_6061; // @[executor.scala 473:84]
  wire [7:0] _GEN_6482 = _GEN_8850 == 8'h28 ? _GEN_6478 : _GEN_6062; // @[executor.scala 473:84]
  wire [7:0] _GEN_6483 = _GEN_8850 == 8'h28 ? _GEN_6479 : _GEN_6063; // @[executor.scala 473:84]
  wire [7:0] _GEN_6484 = mask_6[0] ? byte_1536 : _GEN_6064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6485 = mask_6[1] ? byte_1537 : _GEN_6065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6486 = mask_6[2] ? byte_1538 : _GEN_6066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6487 = mask_6[3] ? byte_1539 : _GEN_6067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6488 = _GEN_8850 == 8'h29 ? _GEN_6484 : _GEN_6064; // @[executor.scala 473:84]
  wire [7:0] _GEN_6489 = _GEN_8850 == 8'h29 ? _GEN_6485 : _GEN_6065; // @[executor.scala 473:84]
  wire [7:0] _GEN_6490 = _GEN_8850 == 8'h29 ? _GEN_6486 : _GEN_6066; // @[executor.scala 473:84]
  wire [7:0] _GEN_6491 = _GEN_8850 == 8'h29 ? _GEN_6487 : _GEN_6067; // @[executor.scala 473:84]
  wire [7:0] _GEN_6492 = mask_6[0] ? byte_1536 : _GEN_6068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6493 = mask_6[1] ? byte_1537 : _GEN_6069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6494 = mask_6[2] ? byte_1538 : _GEN_6070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6495 = mask_6[3] ? byte_1539 : _GEN_6071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6496 = _GEN_8850 == 8'h2a ? _GEN_6492 : _GEN_6068; // @[executor.scala 473:84]
  wire [7:0] _GEN_6497 = _GEN_8850 == 8'h2a ? _GEN_6493 : _GEN_6069; // @[executor.scala 473:84]
  wire [7:0] _GEN_6498 = _GEN_8850 == 8'h2a ? _GEN_6494 : _GEN_6070; // @[executor.scala 473:84]
  wire [7:0] _GEN_6499 = _GEN_8850 == 8'h2a ? _GEN_6495 : _GEN_6071; // @[executor.scala 473:84]
  wire [7:0] _GEN_6500 = mask_6[0] ? byte_1536 : _GEN_6072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6501 = mask_6[1] ? byte_1537 : _GEN_6073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6502 = mask_6[2] ? byte_1538 : _GEN_6074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6503 = mask_6[3] ? byte_1539 : _GEN_6075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6504 = _GEN_8850 == 8'h2b ? _GEN_6500 : _GEN_6072; // @[executor.scala 473:84]
  wire [7:0] _GEN_6505 = _GEN_8850 == 8'h2b ? _GEN_6501 : _GEN_6073; // @[executor.scala 473:84]
  wire [7:0] _GEN_6506 = _GEN_8850 == 8'h2b ? _GEN_6502 : _GEN_6074; // @[executor.scala 473:84]
  wire [7:0] _GEN_6507 = _GEN_8850 == 8'h2b ? _GEN_6503 : _GEN_6075; // @[executor.scala 473:84]
  wire [7:0] _GEN_6508 = mask_6[0] ? byte_1536 : _GEN_6076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6509 = mask_6[1] ? byte_1537 : _GEN_6077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6510 = mask_6[2] ? byte_1538 : _GEN_6078; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6511 = mask_6[3] ? byte_1539 : _GEN_6079; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6512 = _GEN_8850 == 8'h2c ? _GEN_6508 : _GEN_6076; // @[executor.scala 473:84]
  wire [7:0] _GEN_6513 = _GEN_8850 == 8'h2c ? _GEN_6509 : _GEN_6077; // @[executor.scala 473:84]
  wire [7:0] _GEN_6514 = _GEN_8850 == 8'h2c ? _GEN_6510 : _GEN_6078; // @[executor.scala 473:84]
  wire [7:0] _GEN_6515 = _GEN_8850 == 8'h2c ? _GEN_6511 : _GEN_6079; // @[executor.scala 473:84]
  wire [7:0] _GEN_6516 = mask_6[0] ? byte_1536 : _GEN_6080; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6517 = mask_6[1] ? byte_1537 : _GEN_6081; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6518 = mask_6[2] ? byte_1538 : _GEN_6082; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6519 = mask_6[3] ? byte_1539 : _GEN_6083; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6520 = _GEN_8850 == 8'h2d ? _GEN_6516 : _GEN_6080; // @[executor.scala 473:84]
  wire [7:0] _GEN_6521 = _GEN_8850 == 8'h2d ? _GEN_6517 : _GEN_6081; // @[executor.scala 473:84]
  wire [7:0] _GEN_6522 = _GEN_8850 == 8'h2d ? _GEN_6518 : _GEN_6082; // @[executor.scala 473:84]
  wire [7:0] _GEN_6523 = _GEN_8850 == 8'h2d ? _GEN_6519 : _GEN_6083; // @[executor.scala 473:84]
  wire [7:0] _GEN_6524 = mask_6[0] ? byte_1536 : _GEN_6084; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6525 = mask_6[1] ? byte_1537 : _GEN_6085; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6526 = mask_6[2] ? byte_1538 : _GEN_6086; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6527 = mask_6[3] ? byte_1539 : _GEN_6087; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6528 = _GEN_8850 == 8'h2e ? _GEN_6524 : _GEN_6084; // @[executor.scala 473:84]
  wire [7:0] _GEN_6529 = _GEN_8850 == 8'h2e ? _GEN_6525 : _GEN_6085; // @[executor.scala 473:84]
  wire [7:0] _GEN_6530 = _GEN_8850 == 8'h2e ? _GEN_6526 : _GEN_6086; // @[executor.scala 473:84]
  wire [7:0] _GEN_6531 = _GEN_8850 == 8'h2e ? _GEN_6527 : _GEN_6087; // @[executor.scala 473:84]
  wire [7:0] _GEN_6532 = mask_6[0] ? byte_1536 : _GEN_6088; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6533 = mask_6[1] ? byte_1537 : _GEN_6089; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6534 = mask_6[2] ? byte_1538 : _GEN_6090; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6535 = mask_6[3] ? byte_1539 : _GEN_6091; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6536 = _GEN_8850 == 8'h2f ? _GEN_6532 : _GEN_6088; // @[executor.scala 473:84]
  wire [7:0] _GEN_6537 = _GEN_8850 == 8'h2f ? _GEN_6533 : _GEN_6089; // @[executor.scala 473:84]
  wire [7:0] _GEN_6538 = _GEN_8850 == 8'h2f ? _GEN_6534 : _GEN_6090; // @[executor.scala 473:84]
  wire [7:0] _GEN_6539 = _GEN_8850 == 8'h2f ? _GEN_6535 : _GEN_6091; // @[executor.scala 473:84]
  wire [7:0] _GEN_6540 = mask_6[0] ? byte_1536 : _GEN_6092; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6541 = mask_6[1] ? byte_1537 : _GEN_6093; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6542 = mask_6[2] ? byte_1538 : _GEN_6094; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6543 = mask_6[3] ? byte_1539 : _GEN_6095; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6544 = _GEN_8850 == 8'h30 ? _GEN_6540 : _GEN_6092; // @[executor.scala 473:84]
  wire [7:0] _GEN_6545 = _GEN_8850 == 8'h30 ? _GEN_6541 : _GEN_6093; // @[executor.scala 473:84]
  wire [7:0] _GEN_6546 = _GEN_8850 == 8'h30 ? _GEN_6542 : _GEN_6094; // @[executor.scala 473:84]
  wire [7:0] _GEN_6547 = _GEN_8850 == 8'h30 ? _GEN_6543 : _GEN_6095; // @[executor.scala 473:84]
  wire [7:0] _GEN_6548 = mask_6[0] ? byte_1536 : _GEN_6096; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6549 = mask_6[1] ? byte_1537 : _GEN_6097; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6550 = mask_6[2] ? byte_1538 : _GEN_6098; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6551 = mask_6[3] ? byte_1539 : _GEN_6099; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6552 = _GEN_8850 == 8'h31 ? _GEN_6548 : _GEN_6096; // @[executor.scala 473:84]
  wire [7:0] _GEN_6553 = _GEN_8850 == 8'h31 ? _GEN_6549 : _GEN_6097; // @[executor.scala 473:84]
  wire [7:0] _GEN_6554 = _GEN_8850 == 8'h31 ? _GEN_6550 : _GEN_6098; // @[executor.scala 473:84]
  wire [7:0] _GEN_6555 = _GEN_8850 == 8'h31 ? _GEN_6551 : _GEN_6099; // @[executor.scala 473:84]
  wire [7:0] _GEN_6556 = mask_6[0] ? byte_1536 : _GEN_6100; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6557 = mask_6[1] ? byte_1537 : _GEN_6101; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6558 = mask_6[2] ? byte_1538 : _GEN_6102; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6559 = mask_6[3] ? byte_1539 : _GEN_6103; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6560 = _GEN_8850 == 8'h32 ? _GEN_6556 : _GEN_6100; // @[executor.scala 473:84]
  wire [7:0] _GEN_6561 = _GEN_8850 == 8'h32 ? _GEN_6557 : _GEN_6101; // @[executor.scala 473:84]
  wire [7:0] _GEN_6562 = _GEN_8850 == 8'h32 ? _GEN_6558 : _GEN_6102; // @[executor.scala 473:84]
  wire [7:0] _GEN_6563 = _GEN_8850 == 8'h32 ? _GEN_6559 : _GEN_6103; // @[executor.scala 473:84]
  wire [7:0] _GEN_6564 = mask_6[0] ? byte_1536 : _GEN_6104; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6565 = mask_6[1] ? byte_1537 : _GEN_6105; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6566 = mask_6[2] ? byte_1538 : _GEN_6106; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6567 = mask_6[3] ? byte_1539 : _GEN_6107; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6568 = _GEN_8850 == 8'h33 ? _GEN_6564 : _GEN_6104; // @[executor.scala 473:84]
  wire [7:0] _GEN_6569 = _GEN_8850 == 8'h33 ? _GEN_6565 : _GEN_6105; // @[executor.scala 473:84]
  wire [7:0] _GEN_6570 = _GEN_8850 == 8'h33 ? _GEN_6566 : _GEN_6106; // @[executor.scala 473:84]
  wire [7:0] _GEN_6571 = _GEN_8850 == 8'h33 ? _GEN_6567 : _GEN_6107; // @[executor.scala 473:84]
  wire [7:0] _GEN_6572 = mask_6[0] ? byte_1536 : _GEN_6108; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6573 = mask_6[1] ? byte_1537 : _GEN_6109; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6574 = mask_6[2] ? byte_1538 : _GEN_6110; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6575 = mask_6[3] ? byte_1539 : _GEN_6111; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6576 = _GEN_8850 == 8'h34 ? _GEN_6572 : _GEN_6108; // @[executor.scala 473:84]
  wire [7:0] _GEN_6577 = _GEN_8850 == 8'h34 ? _GEN_6573 : _GEN_6109; // @[executor.scala 473:84]
  wire [7:0] _GEN_6578 = _GEN_8850 == 8'h34 ? _GEN_6574 : _GEN_6110; // @[executor.scala 473:84]
  wire [7:0] _GEN_6579 = _GEN_8850 == 8'h34 ? _GEN_6575 : _GEN_6111; // @[executor.scala 473:84]
  wire [7:0] _GEN_6580 = mask_6[0] ? byte_1536 : _GEN_6112; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6581 = mask_6[1] ? byte_1537 : _GEN_6113; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6582 = mask_6[2] ? byte_1538 : _GEN_6114; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6583 = mask_6[3] ? byte_1539 : _GEN_6115; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6584 = _GEN_8850 == 8'h35 ? _GEN_6580 : _GEN_6112; // @[executor.scala 473:84]
  wire [7:0] _GEN_6585 = _GEN_8850 == 8'h35 ? _GEN_6581 : _GEN_6113; // @[executor.scala 473:84]
  wire [7:0] _GEN_6586 = _GEN_8850 == 8'h35 ? _GEN_6582 : _GEN_6114; // @[executor.scala 473:84]
  wire [7:0] _GEN_6587 = _GEN_8850 == 8'h35 ? _GEN_6583 : _GEN_6115; // @[executor.scala 473:84]
  wire [7:0] _GEN_6588 = mask_6[0] ? byte_1536 : _GEN_6116; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6589 = mask_6[1] ? byte_1537 : _GEN_6117; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6590 = mask_6[2] ? byte_1538 : _GEN_6118; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6591 = mask_6[3] ? byte_1539 : _GEN_6119; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6592 = _GEN_8850 == 8'h36 ? _GEN_6588 : _GEN_6116; // @[executor.scala 473:84]
  wire [7:0] _GEN_6593 = _GEN_8850 == 8'h36 ? _GEN_6589 : _GEN_6117; // @[executor.scala 473:84]
  wire [7:0] _GEN_6594 = _GEN_8850 == 8'h36 ? _GEN_6590 : _GEN_6118; // @[executor.scala 473:84]
  wire [7:0] _GEN_6595 = _GEN_8850 == 8'h36 ? _GEN_6591 : _GEN_6119; // @[executor.scala 473:84]
  wire [7:0] _GEN_6596 = mask_6[0] ? byte_1536 : _GEN_6120; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6597 = mask_6[1] ? byte_1537 : _GEN_6121; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6598 = mask_6[2] ? byte_1538 : _GEN_6122; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6599 = mask_6[3] ? byte_1539 : _GEN_6123; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6600 = _GEN_8850 == 8'h37 ? _GEN_6596 : _GEN_6120; // @[executor.scala 473:84]
  wire [7:0] _GEN_6601 = _GEN_8850 == 8'h37 ? _GEN_6597 : _GEN_6121; // @[executor.scala 473:84]
  wire [7:0] _GEN_6602 = _GEN_8850 == 8'h37 ? _GEN_6598 : _GEN_6122; // @[executor.scala 473:84]
  wire [7:0] _GEN_6603 = _GEN_8850 == 8'h37 ? _GEN_6599 : _GEN_6123; // @[executor.scala 473:84]
  wire [7:0] _GEN_6604 = mask_6[0] ? byte_1536 : _GEN_6124; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6605 = mask_6[1] ? byte_1537 : _GEN_6125; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6606 = mask_6[2] ? byte_1538 : _GEN_6126; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6607 = mask_6[3] ? byte_1539 : _GEN_6127; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6608 = _GEN_8850 == 8'h38 ? _GEN_6604 : _GEN_6124; // @[executor.scala 473:84]
  wire [7:0] _GEN_6609 = _GEN_8850 == 8'h38 ? _GEN_6605 : _GEN_6125; // @[executor.scala 473:84]
  wire [7:0] _GEN_6610 = _GEN_8850 == 8'h38 ? _GEN_6606 : _GEN_6126; // @[executor.scala 473:84]
  wire [7:0] _GEN_6611 = _GEN_8850 == 8'h38 ? _GEN_6607 : _GEN_6127; // @[executor.scala 473:84]
  wire [7:0] _GEN_6612 = mask_6[0] ? byte_1536 : _GEN_6128; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6613 = mask_6[1] ? byte_1537 : _GEN_6129; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6614 = mask_6[2] ? byte_1538 : _GEN_6130; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6615 = mask_6[3] ? byte_1539 : _GEN_6131; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6616 = _GEN_8850 == 8'h39 ? _GEN_6612 : _GEN_6128; // @[executor.scala 473:84]
  wire [7:0] _GEN_6617 = _GEN_8850 == 8'h39 ? _GEN_6613 : _GEN_6129; // @[executor.scala 473:84]
  wire [7:0] _GEN_6618 = _GEN_8850 == 8'h39 ? _GEN_6614 : _GEN_6130; // @[executor.scala 473:84]
  wire [7:0] _GEN_6619 = _GEN_8850 == 8'h39 ? _GEN_6615 : _GEN_6131; // @[executor.scala 473:84]
  wire [7:0] _GEN_6620 = mask_6[0] ? byte_1536 : _GEN_6132; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6621 = mask_6[1] ? byte_1537 : _GEN_6133; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6622 = mask_6[2] ? byte_1538 : _GEN_6134; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6623 = mask_6[3] ? byte_1539 : _GEN_6135; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6624 = _GEN_8850 == 8'h3a ? _GEN_6620 : _GEN_6132; // @[executor.scala 473:84]
  wire [7:0] _GEN_6625 = _GEN_8850 == 8'h3a ? _GEN_6621 : _GEN_6133; // @[executor.scala 473:84]
  wire [7:0] _GEN_6626 = _GEN_8850 == 8'h3a ? _GEN_6622 : _GEN_6134; // @[executor.scala 473:84]
  wire [7:0] _GEN_6627 = _GEN_8850 == 8'h3a ? _GEN_6623 : _GEN_6135; // @[executor.scala 473:84]
  wire [7:0] _GEN_6628 = mask_6[0] ? byte_1536 : _GEN_6136; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6629 = mask_6[1] ? byte_1537 : _GEN_6137; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6630 = mask_6[2] ? byte_1538 : _GEN_6138; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6631 = mask_6[3] ? byte_1539 : _GEN_6139; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6632 = _GEN_8850 == 8'h3b ? _GEN_6628 : _GEN_6136; // @[executor.scala 473:84]
  wire [7:0] _GEN_6633 = _GEN_8850 == 8'h3b ? _GEN_6629 : _GEN_6137; // @[executor.scala 473:84]
  wire [7:0] _GEN_6634 = _GEN_8850 == 8'h3b ? _GEN_6630 : _GEN_6138; // @[executor.scala 473:84]
  wire [7:0] _GEN_6635 = _GEN_8850 == 8'h3b ? _GEN_6631 : _GEN_6139; // @[executor.scala 473:84]
  wire [7:0] _GEN_6636 = mask_6[0] ? byte_1536 : _GEN_6140; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6637 = mask_6[1] ? byte_1537 : _GEN_6141; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6638 = mask_6[2] ? byte_1538 : _GEN_6142; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6639 = mask_6[3] ? byte_1539 : _GEN_6143; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6640 = _GEN_8850 == 8'h3c ? _GEN_6636 : _GEN_6140; // @[executor.scala 473:84]
  wire [7:0] _GEN_6641 = _GEN_8850 == 8'h3c ? _GEN_6637 : _GEN_6141; // @[executor.scala 473:84]
  wire [7:0] _GEN_6642 = _GEN_8850 == 8'h3c ? _GEN_6638 : _GEN_6142; // @[executor.scala 473:84]
  wire [7:0] _GEN_6643 = _GEN_8850 == 8'h3c ? _GEN_6639 : _GEN_6143; // @[executor.scala 473:84]
  wire [7:0] _GEN_6644 = mask_6[0] ? byte_1536 : _GEN_6144; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6645 = mask_6[1] ? byte_1537 : _GEN_6145; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6646 = mask_6[2] ? byte_1538 : _GEN_6146; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6647 = mask_6[3] ? byte_1539 : _GEN_6147; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6648 = _GEN_8850 == 8'h3d ? _GEN_6644 : _GEN_6144; // @[executor.scala 473:84]
  wire [7:0] _GEN_6649 = _GEN_8850 == 8'h3d ? _GEN_6645 : _GEN_6145; // @[executor.scala 473:84]
  wire [7:0] _GEN_6650 = _GEN_8850 == 8'h3d ? _GEN_6646 : _GEN_6146; // @[executor.scala 473:84]
  wire [7:0] _GEN_6651 = _GEN_8850 == 8'h3d ? _GEN_6647 : _GEN_6147; // @[executor.scala 473:84]
  wire [7:0] _GEN_6652 = mask_6[0] ? byte_1536 : _GEN_6148; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6653 = mask_6[1] ? byte_1537 : _GEN_6149; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6654 = mask_6[2] ? byte_1538 : _GEN_6150; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6655 = mask_6[3] ? byte_1539 : _GEN_6151; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6656 = _GEN_8850 == 8'h3e ? _GEN_6652 : _GEN_6148; // @[executor.scala 473:84]
  wire [7:0] _GEN_6657 = _GEN_8850 == 8'h3e ? _GEN_6653 : _GEN_6149; // @[executor.scala 473:84]
  wire [7:0] _GEN_6658 = _GEN_8850 == 8'h3e ? _GEN_6654 : _GEN_6150; // @[executor.scala 473:84]
  wire [7:0] _GEN_6659 = _GEN_8850 == 8'h3e ? _GEN_6655 : _GEN_6151; // @[executor.scala 473:84]
  wire [7:0] _GEN_6660 = mask_6[0] ? byte_1536 : _GEN_6152; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6661 = mask_6[1] ? byte_1537 : _GEN_6153; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6662 = mask_6[2] ? byte_1538 : _GEN_6154; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6663 = mask_6[3] ? byte_1539 : _GEN_6155; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6664 = _GEN_8850 == 8'h3f ? _GEN_6660 : _GEN_6152; // @[executor.scala 473:84]
  wire [7:0] _GEN_6665 = _GEN_8850 == 8'h3f ? _GEN_6661 : _GEN_6153; // @[executor.scala 473:84]
  wire [7:0] _GEN_6666 = _GEN_8850 == 8'h3f ? _GEN_6662 : _GEN_6154; // @[executor.scala 473:84]
  wire [7:0] _GEN_6667 = _GEN_8850 == 8'h3f ? _GEN_6663 : _GEN_6155; // @[executor.scala 473:84]
  wire [7:0] _GEN_6668 = opcode_6 != 4'h0 ? _GEN_6160 : _GEN_5900; // @[executor.scala 470:55]
  wire [7:0] _GEN_6669 = opcode_6 != 4'h0 ? _GEN_6161 : _GEN_5901; // @[executor.scala 470:55]
  wire [7:0] _GEN_6670 = opcode_6 != 4'h0 ? _GEN_6162 : _GEN_5902; // @[executor.scala 470:55]
  wire [7:0] _GEN_6671 = opcode_6 != 4'h0 ? _GEN_6163 : _GEN_5903; // @[executor.scala 470:55]
  wire [7:0] _GEN_6672 = opcode_6 != 4'h0 ? _GEN_6168 : _GEN_5904; // @[executor.scala 470:55]
  wire [7:0] _GEN_6673 = opcode_6 != 4'h0 ? _GEN_6169 : _GEN_5905; // @[executor.scala 470:55]
  wire [7:0] _GEN_6674 = opcode_6 != 4'h0 ? _GEN_6170 : _GEN_5906; // @[executor.scala 470:55]
  wire [7:0] _GEN_6675 = opcode_6 != 4'h0 ? _GEN_6171 : _GEN_5907; // @[executor.scala 470:55]
  wire [7:0] _GEN_6676 = opcode_6 != 4'h0 ? _GEN_6176 : _GEN_5908; // @[executor.scala 470:55]
  wire [7:0] _GEN_6677 = opcode_6 != 4'h0 ? _GEN_6177 : _GEN_5909; // @[executor.scala 470:55]
  wire [7:0] _GEN_6678 = opcode_6 != 4'h0 ? _GEN_6178 : _GEN_5910; // @[executor.scala 470:55]
  wire [7:0] _GEN_6679 = opcode_6 != 4'h0 ? _GEN_6179 : _GEN_5911; // @[executor.scala 470:55]
  wire [7:0] _GEN_6680 = opcode_6 != 4'h0 ? _GEN_6184 : _GEN_5912; // @[executor.scala 470:55]
  wire [7:0] _GEN_6681 = opcode_6 != 4'h0 ? _GEN_6185 : _GEN_5913; // @[executor.scala 470:55]
  wire [7:0] _GEN_6682 = opcode_6 != 4'h0 ? _GEN_6186 : _GEN_5914; // @[executor.scala 470:55]
  wire [7:0] _GEN_6683 = opcode_6 != 4'h0 ? _GEN_6187 : _GEN_5915; // @[executor.scala 470:55]
  wire [7:0] _GEN_6684 = opcode_6 != 4'h0 ? _GEN_6192 : _GEN_5916; // @[executor.scala 470:55]
  wire [7:0] _GEN_6685 = opcode_6 != 4'h0 ? _GEN_6193 : _GEN_5917; // @[executor.scala 470:55]
  wire [7:0] _GEN_6686 = opcode_6 != 4'h0 ? _GEN_6194 : _GEN_5918; // @[executor.scala 470:55]
  wire [7:0] _GEN_6687 = opcode_6 != 4'h0 ? _GEN_6195 : _GEN_5919; // @[executor.scala 470:55]
  wire [7:0] _GEN_6688 = opcode_6 != 4'h0 ? _GEN_6200 : _GEN_5920; // @[executor.scala 470:55]
  wire [7:0] _GEN_6689 = opcode_6 != 4'h0 ? _GEN_6201 : _GEN_5921; // @[executor.scala 470:55]
  wire [7:0] _GEN_6690 = opcode_6 != 4'h0 ? _GEN_6202 : _GEN_5922; // @[executor.scala 470:55]
  wire [7:0] _GEN_6691 = opcode_6 != 4'h0 ? _GEN_6203 : _GEN_5923; // @[executor.scala 470:55]
  wire [7:0] _GEN_6692 = opcode_6 != 4'h0 ? _GEN_6208 : _GEN_5924; // @[executor.scala 470:55]
  wire [7:0] _GEN_6693 = opcode_6 != 4'h0 ? _GEN_6209 : _GEN_5925; // @[executor.scala 470:55]
  wire [7:0] _GEN_6694 = opcode_6 != 4'h0 ? _GEN_6210 : _GEN_5926; // @[executor.scala 470:55]
  wire [7:0] _GEN_6695 = opcode_6 != 4'h0 ? _GEN_6211 : _GEN_5927; // @[executor.scala 470:55]
  wire [7:0] _GEN_6696 = opcode_6 != 4'h0 ? _GEN_6216 : _GEN_5928; // @[executor.scala 470:55]
  wire [7:0] _GEN_6697 = opcode_6 != 4'h0 ? _GEN_6217 : _GEN_5929; // @[executor.scala 470:55]
  wire [7:0] _GEN_6698 = opcode_6 != 4'h0 ? _GEN_6218 : _GEN_5930; // @[executor.scala 470:55]
  wire [7:0] _GEN_6699 = opcode_6 != 4'h0 ? _GEN_6219 : _GEN_5931; // @[executor.scala 470:55]
  wire [7:0] _GEN_6700 = opcode_6 != 4'h0 ? _GEN_6224 : _GEN_5932; // @[executor.scala 470:55]
  wire [7:0] _GEN_6701 = opcode_6 != 4'h0 ? _GEN_6225 : _GEN_5933; // @[executor.scala 470:55]
  wire [7:0] _GEN_6702 = opcode_6 != 4'h0 ? _GEN_6226 : _GEN_5934; // @[executor.scala 470:55]
  wire [7:0] _GEN_6703 = opcode_6 != 4'h0 ? _GEN_6227 : _GEN_5935; // @[executor.scala 470:55]
  wire [7:0] _GEN_6704 = opcode_6 != 4'h0 ? _GEN_6232 : _GEN_5936; // @[executor.scala 470:55]
  wire [7:0] _GEN_6705 = opcode_6 != 4'h0 ? _GEN_6233 : _GEN_5937; // @[executor.scala 470:55]
  wire [7:0] _GEN_6706 = opcode_6 != 4'h0 ? _GEN_6234 : _GEN_5938; // @[executor.scala 470:55]
  wire [7:0] _GEN_6707 = opcode_6 != 4'h0 ? _GEN_6235 : _GEN_5939; // @[executor.scala 470:55]
  wire [7:0] _GEN_6708 = opcode_6 != 4'h0 ? _GEN_6240 : _GEN_5940; // @[executor.scala 470:55]
  wire [7:0] _GEN_6709 = opcode_6 != 4'h0 ? _GEN_6241 : _GEN_5941; // @[executor.scala 470:55]
  wire [7:0] _GEN_6710 = opcode_6 != 4'h0 ? _GEN_6242 : _GEN_5942; // @[executor.scala 470:55]
  wire [7:0] _GEN_6711 = opcode_6 != 4'h0 ? _GEN_6243 : _GEN_5943; // @[executor.scala 470:55]
  wire [7:0] _GEN_6712 = opcode_6 != 4'h0 ? _GEN_6248 : _GEN_5944; // @[executor.scala 470:55]
  wire [7:0] _GEN_6713 = opcode_6 != 4'h0 ? _GEN_6249 : _GEN_5945; // @[executor.scala 470:55]
  wire [7:0] _GEN_6714 = opcode_6 != 4'h0 ? _GEN_6250 : _GEN_5946; // @[executor.scala 470:55]
  wire [7:0] _GEN_6715 = opcode_6 != 4'h0 ? _GEN_6251 : _GEN_5947; // @[executor.scala 470:55]
  wire [7:0] _GEN_6716 = opcode_6 != 4'h0 ? _GEN_6256 : _GEN_5948; // @[executor.scala 470:55]
  wire [7:0] _GEN_6717 = opcode_6 != 4'h0 ? _GEN_6257 : _GEN_5949; // @[executor.scala 470:55]
  wire [7:0] _GEN_6718 = opcode_6 != 4'h0 ? _GEN_6258 : _GEN_5950; // @[executor.scala 470:55]
  wire [7:0] _GEN_6719 = opcode_6 != 4'h0 ? _GEN_6259 : _GEN_5951; // @[executor.scala 470:55]
  wire [7:0] _GEN_6720 = opcode_6 != 4'h0 ? _GEN_6264 : _GEN_5952; // @[executor.scala 470:55]
  wire [7:0] _GEN_6721 = opcode_6 != 4'h0 ? _GEN_6265 : _GEN_5953; // @[executor.scala 470:55]
  wire [7:0] _GEN_6722 = opcode_6 != 4'h0 ? _GEN_6266 : _GEN_5954; // @[executor.scala 470:55]
  wire [7:0] _GEN_6723 = opcode_6 != 4'h0 ? _GEN_6267 : _GEN_5955; // @[executor.scala 470:55]
  wire [7:0] _GEN_6724 = opcode_6 != 4'h0 ? _GEN_6272 : _GEN_5956; // @[executor.scala 470:55]
  wire [7:0] _GEN_6725 = opcode_6 != 4'h0 ? _GEN_6273 : _GEN_5957; // @[executor.scala 470:55]
  wire [7:0] _GEN_6726 = opcode_6 != 4'h0 ? _GEN_6274 : _GEN_5958; // @[executor.scala 470:55]
  wire [7:0] _GEN_6727 = opcode_6 != 4'h0 ? _GEN_6275 : _GEN_5959; // @[executor.scala 470:55]
  wire [7:0] _GEN_6728 = opcode_6 != 4'h0 ? _GEN_6280 : _GEN_5960; // @[executor.scala 470:55]
  wire [7:0] _GEN_6729 = opcode_6 != 4'h0 ? _GEN_6281 : _GEN_5961; // @[executor.scala 470:55]
  wire [7:0] _GEN_6730 = opcode_6 != 4'h0 ? _GEN_6282 : _GEN_5962; // @[executor.scala 470:55]
  wire [7:0] _GEN_6731 = opcode_6 != 4'h0 ? _GEN_6283 : _GEN_5963; // @[executor.scala 470:55]
  wire [7:0] _GEN_6732 = opcode_6 != 4'h0 ? _GEN_6288 : _GEN_5964; // @[executor.scala 470:55]
  wire [7:0] _GEN_6733 = opcode_6 != 4'h0 ? _GEN_6289 : _GEN_5965; // @[executor.scala 470:55]
  wire [7:0] _GEN_6734 = opcode_6 != 4'h0 ? _GEN_6290 : _GEN_5966; // @[executor.scala 470:55]
  wire [7:0] _GEN_6735 = opcode_6 != 4'h0 ? _GEN_6291 : _GEN_5967; // @[executor.scala 470:55]
  wire [7:0] _GEN_6736 = opcode_6 != 4'h0 ? _GEN_6296 : _GEN_5968; // @[executor.scala 470:55]
  wire [7:0] _GEN_6737 = opcode_6 != 4'h0 ? _GEN_6297 : _GEN_5969; // @[executor.scala 470:55]
  wire [7:0] _GEN_6738 = opcode_6 != 4'h0 ? _GEN_6298 : _GEN_5970; // @[executor.scala 470:55]
  wire [7:0] _GEN_6739 = opcode_6 != 4'h0 ? _GEN_6299 : _GEN_5971; // @[executor.scala 470:55]
  wire [7:0] _GEN_6740 = opcode_6 != 4'h0 ? _GEN_6304 : _GEN_5972; // @[executor.scala 470:55]
  wire [7:0] _GEN_6741 = opcode_6 != 4'h0 ? _GEN_6305 : _GEN_5973; // @[executor.scala 470:55]
  wire [7:0] _GEN_6742 = opcode_6 != 4'h0 ? _GEN_6306 : _GEN_5974; // @[executor.scala 470:55]
  wire [7:0] _GEN_6743 = opcode_6 != 4'h0 ? _GEN_6307 : _GEN_5975; // @[executor.scala 470:55]
  wire [7:0] _GEN_6744 = opcode_6 != 4'h0 ? _GEN_6312 : _GEN_5976; // @[executor.scala 470:55]
  wire [7:0] _GEN_6745 = opcode_6 != 4'h0 ? _GEN_6313 : _GEN_5977; // @[executor.scala 470:55]
  wire [7:0] _GEN_6746 = opcode_6 != 4'h0 ? _GEN_6314 : _GEN_5978; // @[executor.scala 470:55]
  wire [7:0] _GEN_6747 = opcode_6 != 4'h0 ? _GEN_6315 : _GEN_5979; // @[executor.scala 470:55]
  wire [7:0] _GEN_6748 = opcode_6 != 4'h0 ? _GEN_6320 : _GEN_5980; // @[executor.scala 470:55]
  wire [7:0] _GEN_6749 = opcode_6 != 4'h0 ? _GEN_6321 : _GEN_5981; // @[executor.scala 470:55]
  wire [7:0] _GEN_6750 = opcode_6 != 4'h0 ? _GEN_6322 : _GEN_5982; // @[executor.scala 470:55]
  wire [7:0] _GEN_6751 = opcode_6 != 4'h0 ? _GEN_6323 : _GEN_5983; // @[executor.scala 470:55]
  wire [7:0] _GEN_6752 = opcode_6 != 4'h0 ? _GEN_6328 : _GEN_5984; // @[executor.scala 470:55]
  wire [7:0] _GEN_6753 = opcode_6 != 4'h0 ? _GEN_6329 : _GEN_5985; // @[executor.scala 470:55]
  wire [7:0] _GEN_6754 = opcode_6 != 4'h0 ? _GEN_6330 : _GEN_5986; // @[executor.scala 470:55]
  wire [7:0] _GEN_6755 = opcode_6 != 4'h0 ? _GEN_6331 : _GEN_5987; // @[executor.scala 470:55]
  wire [7:0] _GEN_6756 = opcode_6 != 4'h0 ? _GEN_6336 : _GEN_5988; // @[executor.scala 470:55]
  wire [7:0] _GEN_6757 = opcode_6 != 4'h0 ? _GEN_6337 : _GEN_5989; // @[executor.scala 470:55]
  wire [7:0] _GEN_6758 = opcode_6 != 4'h0 ? _GEN_6338 : _GEN_5990; // @[executor.scala 470:55]
  wire [7:0] _GEN_6759 = opcode_6 != 4'h0 ? _GEN_6339 : _GEN_5991; // @[executor.scala 470:55]
  wire [7:0] _GEN_6760 = opcode_6 != 4'h0 ? _GEN_6344 : _GEN_5992; // @[executor.scala 470:55]
  wire [7:0] _GEN_6761 = opcode_6 != 4'h0 ? _GEN_6345 : _GEN_5993; // @[executor.scala 470:55]
  wire [7:0] _GEN_6762 = opcode_6 != 4'h0 ? _GEN_6346 : _GEN_5994; // @[executor.scala 470:55]
  wire [7:0] _GEN_6763 = opcode_6 != 4'h0 ? _GEN_6347 : _GEN_5995; // @[executor.scala 470:55]
  wire [7:0] _GEN_6764 = opcode_6 != 4'h0 ? _GEN_6352 : _GEN_5996; // @[executor.scala 470:55]
  wire [7:0] _GEN_6765 = opcode_6 != 4'h0 ? _GEN_6353 : _GEN_5997; // @[executor.scala 470:55]
  wire [7:0] _GEN_6766 = opcode_6 != 4'h0 ? _GEN_6354 : _GEN_5998; // @[executor.scala 470:55]
  wire [7:0] _GEN_6767 = opcode_6 != 4'h0 ? _GEN_6355 : _GEN_5999; // @[executor.scala 470:55]
  wire [7:0] _GEN_6768 = opcode_6 != 4'h0 ? _GEN_6360 : _GEN_6000; // @[executor.scala 470:55]
  wire [7:0] _GEN_6769 = opcode_6 != 4'h0 ? _GEN_6361 : _GEN_6001; // @[executor.scala 470:55]
  wire [7:0] _GEN_6770 = opcode_6 != 4'h0 ? _GEN_6362 : _GEN_6002; // @[executor.scala 470:55]
  wire [7:0] _GEN_6771 = opcode_6 != 4'h0 ? _GEN_6363 : _GEN_6003; // @[executor.scala 470:55]
  wire [7:0] _GEN_6772 = opcode_6 != 4'h0 ? _GEN_6368 : _GEN_6004; // @[executor.scala 470:55]
  wire [7:0] _GEN_6773 = opcode_6 != 4'h0 ? _GEN_6369 : _GEN_6005; // @[executor.scala 470:55]
  wire [7:0] _GEN_6774 = opcode_6 != 4'h0 ? _GEN_6370 : _GEN_6006; // @[executor.scala 470:55]
  wire [7:0] _GEN_6775 = opcode_6 != 4'h0 ? _GEN_6371 : _GEN_6007; // @[executor.scala 470:55]
  wire [7:0] _GEN_6776 = opcode_6 != 4'h0 ? _GEN_6376 : _GEN_6008; // @[executor.scala 470:55]
  wire [7:0] _GEN_6777 = opcode_6 != 4'h0 ? _GEN_6377 : _GEN_6009; // @[executor.scala 470:55]
  wire [7:0] _GEN_6778 = opcode_6 != 4'h0 ? _GEN_6378 : _GEN_6010; // @[executor.scala 470:55]
  wire [7:0] _GEN_6779 = opcode_6 != 4'h0 ? _GEN_6379 : _GEN_6011; // @[executor.scala 470:55]
  wire [7:0] _GEN_6780 = opcode_6 != 4'h0 ? _GEN_6384 : _GEN_6012; // @[executor.scala 470:55]
  wire [7:0] _GEN_6781 = opcode_6 != 4'h0 ? _GEN_6385 : _GEN_6013; // @[executor.scala 470:55]
  wire [7:0] _GEN_6782 = opcode_6 != 4'h0 ? _GEN_6386 : _GEN_6014; // @[executor.scala 470:55]
  wire [7:0] _GEN_6783 = opcode_6 != 4'h0 ? _GEN_6387 : _GEN_6015; // @[executor.scala 470:55]
  wire [7:0] _GEN_6784 = opcode_6 != 4'h0 ? _GEN_6392 : _GEN_6016; // @[executor.scala 470:55]
  wire [7:0] _GEN_6785 = opcode_6 != 4'h0 ? _GEN_6393 : _GEN_6017; // @[executor.scala 470:55]
  wire [7:0] _GEN_6786 = opcode_6 != 4'h0 ? _GEN_6394 : _GEN_6018; // @[executor.scala 470:55]
  wire [7:0] _GEN_6787 = opcode_6 != 4'h0 ? _GEN_6395 : _GEN_6019; // @[executor.scala 470:55]
  wire [7:0] _GEN_6788 = opcode_6 != 4'h0 ? _GEN_6400 : _GEN_6020; // @[executor.scala 470:55]
  wire [7:0] _GEN_6789 = opcode_6 != 4'h0 ? _GEN_6401 : _GEN_6021; // @[executor.scala 470:55]
  wire [7:0] _GEN_6790 = opcode_6 != 4'h0 ? _GEN_6402 : _GEN_6022; // @[executor.scala 470:55]
  wire [7:0] _GEN_6791 = opcode_6 != 4'h0 ? _GEN_6403 : _GEN_6023; // @[executor.scala 470:55]
  wire [7:0] _GEN_6792 = opcode_6 != 4'h0 ? _GEN_6408 : _GEN_6024; // @[executor.scala 470:55]
  wire [7:0] _GEN_6793 = opcode_6 != 4'h0 ? _GEN_6409 : _GEN_6025; // @[executor.scala 470:55]
  wire [7:0] _GEN_6794 = opcode_6 != 4'h0 ? _GEN_6410 : _GEN_6026; // @[executor.scala 470:55]
  wire [7:0] _GEN_6795 = opcode_6 != 4'h0 ? _GEN_6411 : _GEN_6027; // @[executor.scala 470:55]
  wire [7:0] _GEN_6796 = opcode_6 != 4'h0 ? _GEN_6416 : _GEN_6028; // @[executor.scala 470:55]
  wire [7:0] _GEN_6797 = opcode_6 != 4'h0 ? _GEN_6417 : _GEN_6029; // @[executor.scala 470:55]
  wire [7:0] _GEN_6798 = opcode_6 != 4'h0 ? _GEN_6418 : _GEN_6030; // @[executor.scala 470:55]
  wire [7:0] _GEN_6799 = opcode_6 != 4'h0 ? _GEN_6419 : _GEN_6031; // @[executor.scala 470:55]
  wire [7:0] _GEN_6800 = opcode_6 != 4'h0 ? _GEN_6424 : _GEN_6032; // @[executor.scala 470:55]
  wire [7:0] _GEN_6801 = opcode_6 != 4'h0 ? _GEN_6425 : _GEN_6033; // @[executor.scala 470:55]
  wire [7:0] _GEN_6802 = opcode_6 != 4'h0 ? _GEN_6426 : _GEN_6034; // @[executor.scala 470:55]
  wire [7:0] _GEN_6803 = opcode_6 != 4'h0 ? _GEN_6427 : _GEN_6035; // @[executor.scala 470:55]
  wire [7:0] _GEN_6804 = opcode_6 != 4'h0 ? _GEN_6432 : _GEN_6036; // @[executor.scala 470:55]
  wire [7:0] _GEN_6805 = opcode_6 != 4'h0 ? _GEN_6433 : _GEN_6037; // @[executor.scala 470:55]
  wire [7:0] _GEN_6806 = opcode_6 != 4'h0 ? _GEN_6434 : _GEN_6038; // @[executor.scala 470:55]
  wire [7:0] _GEN_6807 = opcode_6 != 4'h0 ? _GEN_6435 : _GEN_6039; // @[executor.scala 470:55]
  wire [7:0] _GEN_6808 = opcode_6 != 4'h0 ? _GEN_6440 : _GEN_6040; // @[executor.scala 470:55]
  wire [7:0] _GEN_6809 = opcode_6 != 4'h0 ? _GEN_6441 : _GEN_6041; // @[executor.scala 470:55]
  wire [7:0] _GEN_6810 = opcode_6 != 4'h0 ? _GEN_6442 : _GEN_6042; // @[executor.scala 470:55]
  wire [7:0] _GEN_6811 = opcode_6 != 4'h0 ? _GEN_6443 : _GEN_6043; // @[executor.scala 470:55]
  wire [7:0] _GEN_6812 = opcode_6 != 4'h0 ? _GEN_6448 : _GEN_6044; // @[executor.scala 470:55]
  wire [7:0] _GEN_6813 = opcode_6 != 4'h0 ? _GEN_6449 : _GEN_6045; // @[executor.scala 470:55]
  wire [7:0] _GEN_6814 = opcode_6 != 4'h0 ? _GEN_6450 : _GEN_6046; // @[executor.scala 470:55]
  wire [7:0] _GEN_6815 = opcode_6 != 4'h0 ? _GEN_6451 : _GEN_6047; // @[executor.scala 470:55]
  wire [7:0] _GEN_6816 = opcode_6 != 4'h0 ? _GEN_6456 : _GEN_6048; // @[executor.scala 470:55]
  wire [7:0] _GEN_6817 = opcode_6 != 4'h0 ? _GEN_6457 : _GEN_6049; // @[executor.scala 470:55]
  wire [7:0] _GEN_6818 = opcode_6 != 4'h0 ? _GEN_6458 : _GEN_6050; // @[executor.scala 470:55]
  wire [7:0] _GEN_6819 = opcode_6 != 4'h0 ? _GEN_6459 : _GEN_6051; // @[executor.scala 470:55]
  wire [7:0] _GEN_6820 = opcode_6 != 4'h0 ? _GEN_6464 : _GEN_6052; // @[executor.scala 470:55]
  wire [7:0] _GEN_6821 = opcode_6 != 4'h0 ? _GEN_6465 : _GEN_6053; // @[executor.scala 470:55]
  wire [7:0] _GEN_6822 = opcode_6 != 4'h0 ? _GEN_6466 : _GEN_6054; // @[executor.scala 470:55]
  wire [7:0] _GEN_6823 = opcode_6 != 4'h0 ? _GEN_6467 : _GEN_6055; // @[executor.scala 470:55]
  wire [7:0] _GEN_6824 = opcode_6 != 4'h0 ? _GEN_6472 : _GEN_6056; // @[executor.scala 470:55]
  wire [7:0] _GEN_6825 = opcode_6 != 4'h0 ? _GEN_6473 : _GEN_6057; // @[executor.scala 470:55]
  wire [7:0] _GEN_6826 = opcode_6 != 4'h0 ? _GEN_6474 : _GEN_6058; // @[executor.scala 470:55]
  wire [7:0] _GEN_6827 = opcode_6 != 4'h0 ? _GEN_6475 : _GEN_6059; // @[executor.scala 470:55]
  wire [7:0] _GEN_6828 = opcode_6 != 4'h0 ? _GEN_6480 : _GEN_6060; // @[executor.scala 470:55]
  wire [7:0] _GEN_6829 = opcode_6 != 4'h0 ? _GEN_6481 : _GEN_6061; // @[executor.scala 470:55]
  wire [7:0] _GEN_6830 = opcode_6 != 4'h0 ? _GEN_6482 : _GEN_6062; // @[executor.scala 470:55]
  wire [7:0] _GEN_6831 = opcode_6 != 4'h0 ? _GEN_6483 : _GEN_6063; // @[executor.scala 470:55]
  wire [7:0] _GEN_6832 = opcode_6 != 4'h0 ? _GEN_6488 : _GEN_6064; // @[executor.scala 470:55]
  wire [7:0] _GEN_6833 = opcode_6 != 4'h0 ? _GEN_6489 : _GEN_6065; // @[executor.scala 470:55]
  wire [7:0] _GEN_6834 = opcode_6 != 4'h0 ? _GEN_6490 : _GEN_6066; // @[executor.scala 470:55]
  wire [7:0] _GEN_6835 = opcode_6 != 4'h0 ? _GEN_6491 : _GEN_6067; // @[executor.scala 470:55]
  wire [7:0] _GEN_6836 = opcode_6 != 4'h0 ? _GEN_6496 : _GEN_6068; // @[executor.scala 470:55]
  wire [7:0] _GEN_6837 = opcode_6 != 4'h0 ? _GEN_6497 : _GEN_6069; // @[executor.scala 470:55]
  wire [7:0] _GEN_6838 = opcode_6 != 4'h0 ? _GEN_6498 : _GEN_6070; // @[executor.scala 470:55]
  wire [7:0] _GEN_6839 = opcode_6 != 4'h0 ? _GEN_6499 : _GEN_6071; // @[executor.scala 470:55]
  wire [7:0] _GEN_6840 = opcode_6 != 4'h0 ? _GEN_6504 : _GEN_6072; // @[executor.scala 470:55]
  wire [7:0] _GEN_6841 = opcode_6 != 4'h0 ? _GEN_6505 : _GEN_6073; // @[executor.scala 470:55]
  wire [7:0] _GEN_6842 = opcode_6 != 4'h0 ? _GEN_6506 : _GEN_6074; // @[executor.scala 470:55]
  wire [7:0] _GEN_6843 = opcode_6 != 4'h0 ? _GEN_6507 : _GEN_6075; // @[executor.scala 470:55]
  wire [7:0] _GEN_6844 = opcode_6 != 4'h0 ? _GEN_6512 : _GEN_6076; // @[executor.scala 470:55]
  wire [7:0] _GEN_6845 = opcode_6 != 4'h0 ? _GEN_6513 : _GEN_6077; // @[executor.scala 470:55]
  wire [7:0] _GEN_6846 = opcode_6 != 4'h0 ? _GEN_6514 : _GEN_6078; // @[executor.scala 470:55]
  wire [7:0] _GEN_6847 = opcode_6 != 4'h0 ? _GEN_6515 : _GEN_6079; // @[executor.scala 470:55]
  wire [7:0] _GEN_6848 = opcode_6 != 4'h0 ? _GEN_6520 : _GEN_6080; // @[executor.scala 470:55]
  wire [7:0] _GEN_6849 = opcode_6 != 4'h0 ? _GEN_6521 : _GEN_6081; // @[executor.scala 470:55]
  wire [7:0] _GEN_6850 = opcode_6 != 4'h0 ? _GEN_6522 : _GEN_6082; // @[executor.scala 470:55]
  wire [7:0] _GEN_6851 = opcode_6 != 4'h0 ? _GEN_6523 : _GEN_6083; // @[executor.scala 470:55]
  wire [7:0] _GEN_6852 = opcode_6 != 4'h0 ? _GEN_6528 : _GEN_6084; // @[executor.scala 470:55]
  wire [7:0] _GEN_6853 = opcode_6 != 4'h0 ? _GEN_6529 : _GEN_6085; // @[executor.scala 470:55]
  wire [7:0] _GEN_6854 = opcode_6 != 4'h0 ? _GEN_6530 : _GEN_6086; // @[executor.scala 470:55]
  wire [7:0] _GEN_6855 = opcode_6 != 4'h0 ? _GEN_6531 : _GEN_6087; // @[executor.scala 470:55]
  wire [7:0] _GEN_6856 = opcode_6 != 4'h0 ? _GEN_6536 : _GEN_6088; // @[executor.scala 470:55]
  wire [7:0] _GEN_6857 = opcode_6 != 4'h0 ? _GEN_6537 : _GEN_6089; // @[executor.scala 470:55]
  wire [7:0] _GEN_6858 = opcode_6 != 4'h0 ? _GEN_6538 : _GEN_6090; // @[executor.scala 470:55]
  wire [7:0] _GEN_6859 = opcode_6 != 4'h0 ? _GEN_6539 : _GEN_6091; // @[executor.scala 470:55]
  wire [7:0] _GEN_6860 = opcode_6 != 4'h0 ? _GEN_6544 : _GEN_6092; // @[executor.scala 470:55]
  wire [7:0] _GEN_6861 = opcode_6 != 4'h0 ? _GEN_6545 : _GEN_6093; // @[executor.scala 470:55]
  wire [7:0] _GEN_6862 = opcode_6 != 4'h0 ? _GEN_6546 : _GEN_6094; // @[executor.scala 470:55]
  wire [7:0] _GEN_6863 = opcode_6 != 4'h0 ? _GEN_6547 : _GEN_6095; // @[executor.scala 470:55]
  wire [7:0] _GEN_6864 = opcode_6 != 4'h0 ? _GEN_6552 : _GEN_6096; // @[executor.scala 470:55]
  wire [7:0] _GEN_6865 = opcode_6 != 4'h0 ? _GEN_6553 : _GEN_6097; // @[executor.scala 470:55]
  wire [7:0] _GEN_6866 = opcode_6 != 4'h0 ? _GEN_6554 : _GEN_6098; // @[executor.scala 470:55]
  wire [7:0] _GEN_6867 = opcode_6 != 4'h0 ? _GEN_6555 : _GEN_6099; // @[executor.scala 470:55]
  wire [7:0] _GEN_6868 = opcode_6 != 4'h0 ? _GEN_6560 : _GEN_6100; // @[executor.scala 470:55]
  wire [7:0] _GEN_6869 = opcode_6 != 4'h0 ? _GEN_6561 : _GEN_6101; // @[executor.scala 470:55]
  wire [7:0] _GEN_6870 = opcode_6 != 4'h0 ? _GEN_6562 : _GEN_6102; // @[executor.scala 470:55]
  wire [7:0] _GEN_6871 = opcode_6 != 4'h0 ? _GEN_6563 : _GEN_6103; // @[executor.scala 470:55]
  wire [7:0] _GEN_6872 = opcode_6 != 4'h0 ? _GEN_6568 : _GEN_6104; // @[executor.scala 470:55]
  wire [7:0] _GEN_6873 = opcode_6 != 4'h0 ? _GEN_6569 : _GEN_6105; // @[executor.scala 470:55]
  wire [7:0] _GEN_6874 = opcode_6 != 4'h0 ? _GEN_6570 : _GEN_6106; // @[executor.scala 470:55]
  wire [7:0] _GEN_6875 = opcode_6 != 4'h0 ? _GEN_6571 : _GEN_6107; // @[executor.scala 470:55]
  wire [7:0] _GEN_6876 = opcode_6 != 4'h0 ? _GEN_6576 : _GEN_6108; // @[executor.scala 470:55]
  wire [7:0] _GEN_6877 = opcode_6 != 4'h0 ? _GEN_6577 : _GEN_6109; // @[executor.scala 470:55]
  wire [7:0] _GEN_6878 = opcode_6 != 4'h0 ? _GEN_6578 : _GEN_6110; // @[executor.scala 470:55]
  wire [7:0] _GEN_6879 = opcode_6 != 4'h0 ? _GEN_6579 : _GEN_6111; // @[executor.scala 470:55]
  wire [7:0] _GEN_6880 = opcode_6 != 4'h0 ? _GEN_6584 : _GEN_6112; // @[executor.scala 470:55]
  wire [7:0] _GEN_6881 = opcode_6 != 4'h0 ? _GEN_6585 : _GEN_6113; // @[executor.scala 470:55]
  wire [7:0] _GEN_6882 = opcode_6 != 4'h0 ? _GEN_6586 : _GEN_6114; // @[executor.scala 470:55]
  wire [7:0] _GEN_6883 = opcode_6 != 4'h0 ? _GEN_6587 : _GEN_6115; // @[executor.scala 470:55]
  wire [7:0] _GEN_6884 = opcode_6 != 4'h0 ? _GEN_6592 : _GEN_6116; // @[executor.scala 470:55]
  wire [7:0] _GEN_6885 = opcode_6 != 4'h0 ? _GEN_6593 : _GEN_6117; // @[executor.scala 470:55]
  wire [7:0] _GEN_6886 = opcode_6 != 4'h0 ? _GEN_6594 : _GEN_6118; // @[executor.scala 470:55]
  wire [7:0] _GEN_6887 = opcode_6 != 4'h0 ? _GEN_6595 : _GEN_6119; // @[executor.scala 470:55]
  wire [7:0] _GEN_6888 = opcode_6 != 4'h0 ? _GEN_6600 : _GEN_6120; // @[executor.scala 470:55]
  wire [7:0] _GEN_6889 = opcode_6 != 4'h0 ? _GEN_6601 : _GEN_6121; // @[executor.scala 470:55]
  wire [7:0] _GEN_6890 = opcode_6 != 4'h0 ? _GEN_6602 : _GEN_6122; // @[executor.scala 470:55]
  wire [7:0] _GEN_6891 = opcode_6 != 4'h0 ? _GEN_6603 : _GEN_6123; // @[executor.scala 470:55]
  wire [7:0] _GEN_6892 = opcode_6 != 4'h0 ? _GEN_6608 : _GEN_6124; // @[executor.scala 470:55]
  wire [7:0] _GEN_6893 = opcode_6 != 4'h0 ? _GEN_6609 : _GEN_6125; // @[executor.scala 470:55]
  wire [7:0] _GEN_6894 = opcode_6 != 4'h0 ? _GEN_6610 : _GEN_6126; // @[executor.scala 470:55]
  wire [7:0] _GEN_6895 = opcode_6 != 4'h0 ? _GEN_6611 : _GEN_6127; // @[executor.scala 470:55]
  wire [7:0] _GEN_6896 = opcode_6 != 4'h0 ? _GEN_6616 : _GEN_6128; // @[executor.scala 470:55]
  wire [7:0] _GEN_6897 = opcode_6 != 4'h0 ? _GEN_6617 : _GEN_6129; // @[executor.scala 470:55]
  wire [7:0] _GEN_6898 = opcode_6 != 4'h0 ? _GEN_6618 : _GEN_6130; // @[executor.scala 470:55]
  wire [7:0] _GEN_6899 = opcode_6 != 4'h0 ? _GEN_6619 : _GEN_6131; // @[executor.scala 470:55]
  wire [7:0] _GEN_6900 = opcode_6 != 4'h0 ? _GEN_6624 : _GEN_6132; // @[executor.scala 470:55]
  wire [7:0] _GEN_6901 = opcode_6 != 4'h0 ? _GEN_6625 : _GEN_6133; // @[executor.scala 470:55]
  wire [7:0] _GEN_6902 = opcode_6 != 4'h0 ? _GEN_6626 : _GEN_6134; // @[executor.scala 470:55]
  wire [7:0] _GEN_6903 = opcode_6 != 4'h0 ? _GEN_6627 : _GEN_6135; // @[executor.scala 470:55]
  wire [7:0] _GEN_6904 = opcode_6 != 4'h0 ? _GEN_6632 : _GEN_6136; // @[executor.scala 470:55]
  wire [7:0] _GEN_6905 = opcode_6 != 4'h0 ? _GEN_6633 : _GEN_6137; // @[executor.scala 470:55]
  wire [7:0] _GEN_6906 = opcode_6 != 4'h0 ? _GEN_6634 : _GEN_6138; // @[executor.scala 470:55]
  wire [7:0] _GEN_6907 = opcode_6 != 4'h0 ? _GEN_6635 : _GEN_6139; // @[executor.scala 470:55]
  wire [7:0] _GEN_6908 = opcode_6 != 4'h0 ? _GEN_6640 : _GEN_6140; // @[executor.scala 470:55]
  wire [7:0] _GEN_6909 = opcode_6 != 4'h0 ? _GEN_6641 : _GEN_6141; // @[executor.scala 470:55]
  wire [7:0] _GEN_6910 = opcode_6 != 4'h0 ? _GEN_6642 : _GEN_6142; // @[executor.scala 470:55]
  wire [7:0] _GEN_6911 = opcode_6 != 4'h0 ? _GEN_6643 : _GEN_6143; // @[executor.scala 470:55]
  wire [7:0] _GEN_6912 = opcode_6 != 4'h0 ? _GEN_6648 : _GEN_6144; // @[executor.scala 470:55]
  wire [7:0] _GEN_6913 = opcode_6 != 4'h0 ? _GEN_6649 : _GEN_6145; // @[executor.scala 470:55]
  wire [7:0] _GEN_6914 = opcode_6 != 4'h0 ? _GEN_6650 : _GEN_6146; // @[executor.scala 470:55]
  wire [7:0] _GEN_6915 = opcode_6 != 4'h0 ? _GEN_6651 : _GEN_6147; // @[executor.scala 470:55]
  wire [7:0] _GEN_6916 = opcode_6 != 4'h0 ? _GEN_6656 : _GEN_6148; // @[executor.scala 470:55]
  wire [7:0] _GEN_6917 = opcode_6 != 4'h0 ? _GEN_6657 : _GEN_6149; // @[executor.scala 470:55]
  wire [7:0] _GEN_6918 = opcode_6 != 4'h0 ? _GEN_6658 : _GEN_6150; // @[executor.scala 470:55]
  wire [7:0] _GEN_6919 = opcode_6 != 4'h0 ? _GEN_6659 : _GEN_6151; // @[executor.scala 470:55]
  wire [7:0] _GEN_6920 = opcode_6 != 4'h0 ? _GEN_6664 : _GEN_6152; // @[executor.scala 470:55]
  wire [7:0] _GEN_6921 = opcode_6 != 4'h0 ? _GEN_6665 : _GEN_6153; // @[executor.scala 470:55]
  wire [7:0] _GEN_6922 = opcode_6 != 4'h0 ? _GEN_6666 : _GEN_6154; // @[executor.scala 470:55]
  wire [7:0] _GEN_6923 = opcode_6 != 4'h0 ? _GEN_6667 : _GEN_6155; // @[executor.scala 470:55]
  wire [3:0] _GEN_6924 = opcode_6 == 4'hf ? parameter_2_6[13:10] : _GEN_5898; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_6925 = opcode_6 == 4'hf ? parameter_2_6[0] : _GEN_5899; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_6926 = opcode_6 == 4'hf ? _GEN_5900 : _GEN_6668; // @[executor.scala 466:52]
  wire [7:0] _GEN_6927 = opcode_6 == 4'hf ? _GEN_5901 : _GEN_6669; // @[executor.scala 466:52]
  wire [7:0] _GEN_6928 = opcode_6 == 4'hf ? _GEN_5902 : _GEN_6670; // @[executor.scala 466:52]
  wire [7:0] _GEN_6929 = opcode_6 == 4'hf ? _GEN_5903 : _GEN_6671; // @[executor.scala 466:52]
  wire [7:0] _GEN_6930 = opcode_6 == 4'hf ? _GEN_5904 : _GEN_6672; // @[executor.scala 466:52]
  wire [7:0] _GEN_6931 = opcode_6 == 4'hf ? _GEN_5905 : _GEN_6673; // @[executor.scala 466:52]
  wire [7:0] _GEN_6932 = opcode_6 == 4'hf ? _GEN_5906 : _GEN_6674; // @[executor.scala 466:52]
  wire [7:0] _GEN_6933 = opcode_6 == 4'hf ? _GEN_5907 : _GEN_6675; // @[executor.scala 466:52]
  wire [7:0] _GEN_6934 = opcode_6 == 4'hf ? _GEN_5908 : _GEN_6676; // @[executor.scala 466:52]
  wire [7:0] _GEN_6935 = opcode_6 == 4'hf ? _GEN_5909 : _GEN_6677; // @[executor.scala 466:52]
  wire [7:0] _GEN_6936 = opcode_6 == 4'hf ? _GEN_5910 : _GEN_6678; // @[executor.scala 466:52]
  wire [7:0] _GEN_6937 = opcode_6 == 4'hf ? _GEN_5911 : _GEN_6679; // @[executor.scala 466:52]
  wire [7:0] _GEN_6938 = opcode_6 == 4'hf ? _GEN_5912 : _GEN_6680; // @[executor.scala 466:52]
  wire [7:0] _GEN_6939 = opcode_6 == 4'hf ? _GEN_5913 : _GEN_6681; // @[executor.scala 466:52]
  wire [7:0] _GEN_6940 = opcode_6 == 4'hf ? _GEN_5914 : _GEN_6682; // @[executor.scala 466:52]
  wire [7:0] _GEN_6941 = opcode_6 == 4'hf ? _GEN_5915 : _GEN_6683; // @[executor.scala 466:52]
  wire [7:0] _GEN_6942 = opcode_6 == 4'hf ? _GEN_5916 : _GEN_6684; // @[executor.scala 466:52]
  wire [7:0] _GEN_6943 = opcode_6 == 4'hf ? _GEN_5917 : _GEN_6685; // @[executor.scala 466:52]
  wire [7:0] _GEN_6944 = opcode_6 == 4'hf ? _GEN_5918 : _GEN_6686; // @[executor.scala 466:52]
  wire [7:0] _GEN_6945 = opcode_6 == 4'hf ? _GEN_5919 : _GEN_6687; // @[executor.scala 466:52]
  wire [7:0] _GEN_6946 = opcode_6 == 4'hf ? _GEN_5920 : _GEN_6688; // @[executor.scala 466:52]
  wire [7:0] _GEN_6947 = opcode_6 == 4'hf ? _GEN_5921 : _GEN_6689; // @[executor.scala 466:52]
  wire [7:0] _GEN_6948 = opcode_6 == 4'hf ? _GEN_5922 : _GEN_6690; // @[executor.scala 466:52]
  wire [7:0] _GEN_6949 = opcode_6 == 4'hf ? _GEN_5923 : _GEN_6691; // @[executor.scala 466:52]
  wire [7:0] _GEN_6950 = opcode_6 == 4'hf ? _GEN_5924 : _GEN_6692; // @[executor.scala 466:52]
  wire [7:0] _GEN_6951 = opcode_6 == 4'hf ? _GEN_5925 : _GEN_6693; // @[executor.scala 466:52]
  wire [7:0] _GEN_6952 = opcode_6 == 4'hf ? _GEN_5926 : _GEN_6694; // @[executor.scala 466:52]
  wire [7:0] _GEN_6953 = opcode_6 == 4'hf ? _GEN_5927 : _GEN_6695; // @[executor.scala 466:52]
  wire [7:0] _GEN_6954 = opcode_6 == 4'hf ? _GEN_5928 : _GEN_6696; // @[executor.scala 466:52]
  wire [7:0] _GEN_6955 = opcode_6 == 4'hf ? _GEN_5929 : _GEN_6697; // @[executor.scala 466:52]
  wire [7:0] _GEN_6956 = opcode_6 == 4'hf ? _GEN_5930 : _GEN_6698; // @[executor.scala 466:52]
  wire [7:0] _GEN_6957 = opcode_6 == 4'hf ? _GEN_5931 : _GEN_6699; // @[executor.scala 466:52]
  wire [7:0] _GEN_6958 = opcode_6 == 4'hf ? _GEN_5932 : _GEN_6700; // @[executor.scala 466:52]
  wire [7:0] _GEN_6959 = opcode_6 == 4'hf ? _GEN_5933 : _GEN_6701; // @[executor.scala 466:52]
  wire [7:0] _GEN_6960 = opcode_6 == 4'hf ? _GEN_5934 : _GEN_6702; // @[executor.scala 466:52]
  wire [7:0] _GEN_6961 = opcode_6 == 4'hf ? _GEN_5935 : _GEN_6703; // @[executor.scala 466:52]
  wire [7:0] _GEN_6962 = opcode_6 == 4'hf ? _GEN_5936 : _GEN_6704; // @[executor.scala 466:52]
  wire [7:0] _GEN_6963 = opcode_6 == 4'hf ? _GEN_5937 : _GEN_6705; // @[executor.scala 466:52]
  wire [7:0] _GEN_6964 = opcode_6 == 4'hf ? _GEN_5938 : _GEN_6706; // @[executor.scala 466:52]
  wire [7:0] _GEN_6965 = opcode_6 == 4'hf ? _GEN_5939 : _GEN_6707; // @[executor.scala 466:52]
  wire [7:0] _GEN_6966 = opcode_6 == 4'hf ? _GEN_5940 : _GEN_6708; // @[executor.scala 466:52]
  wire [7:0] _GEN_6967 = opcode_6 == 4'hf ? _GEN_5941 : _GEN_6709; // @[executor.scala 466:52]
  wire [7:0] _GEN_6968 = opcode_6 == 4'hf ? _GEN_5942 : _GEN_6710; // @[executor.scala 466:52]
  wire [7:0] _GEN_6969 = opcode_6 == 4'hf ? _GEN_5943 : _GEN_6711; // @[executor.scala 466:52]
  wire [7:0] _GEN_6970 = opcode_6 == 4'hf ? _GEN_5944 : _GEN_6712; // @[executor.scala 466:52]
  wire [7:0] _GEN_6971 = opcode_6 == 4'hf ? _GEN_5945 : _GEN_6713; // @[executor.scala 466:52]
  wire [7:0] _GEN_6972 = opcode_6 == 4'hf ? _GEN_5946 : _GEN_6714; // @[executor.scala 466:52]
  wire [7:0] _GEN_6973 = opcode_6 == 4'hf ? _GEN_5947 : _GEN_6715; // @[executor.scala 466:52]
  wire [7:0] _GEN_6974 = opcode_6 == 4'hf ? _GEN_5948 : _GEN_6716; // @[executor.scala 466:52]
  wire [7:0] _GEN_6975 = opcode_6 == 4'hf ? _GEN_5949 : _GEN_6717; // @[executor.scala 466:52]
  wire [7:0] _GEN_6976 = opcode_6 == 4'hf ? _GEN_5950 : _GEN_6718; // @[executor.scala 466:52]
  wire [7:0] _GEN_6977 = opcode_6 == 4'hf ? _GEN_5951 : _GEN_6719; // @[executor.scala 466:52]
  wire [7:0] _GEN_6978 = opcode_6 == 4'hf ? _GEN_5952 : _GEN_6720; // @[executor.scala 466:52]
  wire [7:0] _GEN_6979 = opcode_6 == 4'hf ? _GEN_5953 : _GEN_6721; // @[executor.scala 466:52]
  wire [7:0] _GEN_6980 = opcode_6 == 4'hf ? _GEN_5954 : _GEN_6722; // @[executor.scala 466:52]
  wire [7:0] _GEN_6981 = opcode_6 == 4'hf ? _GEN_5955 : _GEN_6723; // @[executor.scala 466:52]
  wire [7:0] _GEN_6982 = opcode_6 == 4'hf ? _GEN_5956 : _GEN_6724; // @[executor.scala 466:52]
  wire [7:0] _GEN_6983 = opcode_6 == 4'hf ? _GEN_5957 : _GEN_6725; // @[executor.scala 466:52]
  wire [7:0] _GEN_6984 = opcode_6 == 4'hf ? _GEN_5958 : _GEN_6726; // @[executor.scala 466:52]
  wire [7:0] _GEN_6985 = opcode_6 == 4'hf ? _GEN_5959 : _GEN_6727; // @[executor.scala 466:52]
  wire [7:0] _GEN_6986 = opcode_6 == 4'hf ? _GEN_5960 : _GEN_6728; // @[executor.scala 466:52]
  wire [7:0] _GEN_6987 = opcode_6 == 4'hf ? _GEN_5961 : _GEN_6729; // @[executor.scala 466:52]
  wire [7:0] _GEN_6988 = opcode_6 == 4'hf ? _GEN_5962 : _GEN_6730; // @[executor.scala 466:52]
  wire [7:0] _GEN_6989 = opcode_6 == 4'hf ? _GEN_5963 : _GEN_6731; // @[executor.scala 466:52]
  wire [7:0] _GEN_6990 = opcode_6 == 4'hf ? _GEN_5964 : _GEN_6732; // @[executor.scala 466:52]
  wire [7:0] _GEN_6991 = opcode_6 == 4'hf ? _GEN_5965 : _GEN_6733; // @[executor.scala 466:52]
  wire [7:0] _GEN_6992 = opcode_6 == 4'hf ? _GEN_5966 : _GEN_6734; // @[executor.scala 466:52]
  wire [7:0] _GEN_6993 = opcode_6 == 4'hf ? _GEN_5967 : _GEN_6735; // @[executor.scala 466:52]
  wire [7:0] _GEN_6994 = opcode_6 == 4'hf ? _GEN_5968 : _GEN_6736; // @[executor.scala 466:52]
  wire [7:0] _GEN_6995 = opcode_6 == 4'hf ? _GEN_5969 : _GEN_6737; // @[executor.scala 466:52]
  wire [7:0] _GEN_6996 = opcode_6 == 4'hf ? _GEN_5970 : _GEN_6738; // @[executor.scala 466:52]
  wire [7:0] _GEN_6997 = opcode_6 == 4'hf ? _GEN_5971 : _GEN_6739; // @[executor.scala 466:52]
  wire [7:0] _GEN_6998 = opcode_6 == 4'hf ? _GEN_5972 : _GEN_6740; // @[executor.scala 466:52]
  wire [7:0] _GEN_6999 = opcode_6 == 4'hf ? _GEN_5973 : _GEN_6741; // @[executor.scala 466:52]
  wire [7:0] _GEN_7000 = opcode_6 == 4'hf ? _GEN_5974 : _GEN_6742; // @[executor.scala 466:52]
  wire [7:0] _GEN_7001 = opcode_6 == 4'hf ? _GEN_5975 : _GEN_6743; // @[executor.scala 466:52]
  wire [7:0] _GEN_7002 = opcode_6 == 4'hf ? _GEN_5976 : _GEN_6744; // @[executor.scala 466:52]
  wire [7:0] _GEN_7003 = opcode_6 == 4'hf ? _GEN_5977 : _GEN_6745; // @[executor.scala 466:52]
  wire [7:0] _GEN_7004 = opcode_6 == 4'hf ? _GEN_5978 : _GEN_6746; // @[executor.scala 466:52]
  wire [7:0] _GEN_7005 = opcode_6 == 4'hf ? _GEN_5979 : _GEN_6747; // @[executor.scala 466:52]
  wire [7:0] _GEN_7006 = opcode_6 == 4'hf ? _GEN_5980 : _GEN_6748; // @[executor.scala 466:52]
  wire [7:0] _GEN_7007 = opcode_6 == 4'hf ? _GEN_5981 : _GEN_6749; // @[executor.scala 466:52]
  wire [7:0] _GEN_7008 = opcode_6 == 4'hf ? _GEN_5982 : _GEN_6750; // @[executor.scala 466:52]
  wire [7:0] _GEN_7009 = opcode_6 == 4'hf ? _GEN_5983 : _GEN_6751; // @[executor.scala 466:52]
  wire [7:0] _GEN_7010 = opcode_6 == 4'hf ? _GEN_5984 : _GEN_6752; // @[executor.scala 466:52]
  wire [7:0] _GEN_7011 = opcode_6 == 4'hf ? _GEN_5985 : _GEN_6753; // @[executor.scala 466:52]
  wire [7:0] _GEN_7012 = opcode_6 == 4'hf ? _GEN_5986 : _GEN_6754; // @[executor.scala 466:52]
  wire [7:0] _GEN_7013 = opcode_6 == 4'hf ? _GEN_5987 : _GEN_6755; // @[executor.scala 466:52]
  wire [7:0] _GEN_7014 = opcode_6 == 4'hf ? _GEN_5988 : _GEN_6756; // @[executor.scala 466:52]
  wire [7:0] _GEN_7015 = opcode_6 == 4'hf ? _GEN_5989 : _GEN_6757; // @[executor.scala 466:52]
  wire [7:0] _GEN_7016 = opcode_6 == 4'hf ? _GEN_5990 : _GEN_6758; // @[executor.scala 466:52]
  wire [7:0] _GEN_7017 = opcode_6 == 4'hf ? _GEN_5991 : _GEN_6759; // @[executor.scala 466:52]
  wire [7:0] _GEN_7018 = opcode_6 == 4'hf ? _GEN_5992 : _GEN_6760; // @[executor.scala 466:52]
  wire [7:0] _GEN_7019 = opcode_6 == 4'hf ? _GEN_5993 : _GEN_6761; // @[executor.scala 466:52]
  wire [7:0] _GEN_7020 = opcode_6 == 4'hf ? _GEN_5994 : _GEN_6762; // @[executor.scala 466:52]
  wire [7:0] _GEN_7021 = opcode_6 == 4'hf ? _GEN_5995 : _GEN_6763; // @[executor.scala 466:52]
  wire [7:0] _GEN_7022 = opcode_6 == 4'hf ? _GEN_5996 : _GEN_6764; // @[executor.scala 466:52]
  wire [7:0] _GEN_7023 = opcode_6 == 4'hf ? _GEN_5997 : _GEN_6765; // @[executor.scala 466:52]
  wire [7:0] _GEN_7024 = opcode_6 == 4'hf ? _GEN_5998 : _GEN_6766; // @[executor.scala 466:52]
  wire [7:0] _GEN_7025 = opcode_6 == 4'hf ? _GEN_5999 : _GEN_6767; // @[executor.scala 466:52]
  wire [7:0] _GEN_7026 = opcode_6 == 4'hf ? _GEN_6000 : _GEN_6768; // @[executor.scala 466:52]
  wire [7:0] _GEN_7027 = opcode_6 == 4'hf ? _GEN_6001 : _GEN_6769; // @[executor.scala 466:52]
  wire [7:0] _GEN_7028 = opcode_6 == 4'hf ? _GEN_6002 : _GEN_6770; // @[executor.scala 466:52]
  wire [7:0] _GEN_7029 = opcode_6 == 4'hf ? _GEN_6003 : _GEN_6771; // @[executor.scala 466:52]
  wire [7:0] _GEN_7030 = opcode_6 == 4'hf ? _GEN_6004 : _GEN_6772; // @[executor.scala 466:52]
  wire [7:0] _GEN_7031 = opcode_6 == 4'hf ? _GEN_6005 : _GEN_6773; // @[executor.scala 466:52]
  wire [7:0] _GEN_7032 = opcode_6 == 4'hf ? _GEN_6006 : _GEN_6774; // @[executor.scala 466:52]
  wire [7:0] _GEN_7033 = opcode_6 == 4'hf ? _GEN_6007 : _GEN_6775; // @[executor.scala 466:52]
  wire [7:0] _GEN_7034 = opcode_6 == 4'hf ? _GEN_6008 : _GEN_6776; // @[executor.scala 466:52]
  wire [7:0] _GEN_7035 = opcode_6 == 4'hf ? _GEN_6009 : _GEN_6777; // @[executor.scala 466:52]
  wire [7:0] _GEN_7036 = opcode_6 == 4'hf ? _GEN_6010 : _GEN_6778; // @[executor.scala 466:52]
  wire [7:0] _GEN_7037 = opcode_6 == 4'hf ? _GEN_6011 : _GEN_6779; // @[executor.scala 466:52]
  wire [7:0] _GEN_7038 = opcode_6 == 4'hf ? _GEN_6012 : _GEN_6780; // @[executor.scala 466:52]
  wire [7:0] _GEN_7039 = opcode_6 == 4'hf ? _GEN_6013 : _GEN_6781; // @[executor.scala 466:52]
  wire [7:0] _GEN_7040 = opcode_6 == 4'hf ? _GEN_6014 : _GEN_6782; // @[executor.scala 466:52]
  wire [7:0] _GEN_7041 = opcode_6 == 4'hf ? _GEN_6015 : _GEN_6783; // @[executor.scala 466:52]
  wire [7:0] _GEN_7042 = opcode_6 == 4'hf ? _GEN_6016 : _GEN_6784; // @[executor.scala 466:52]
  wire [7:0] _GEN_7043 = opcode_6 == 4'hf ? _GEN_6017 : _GEN_6785; // @[executor.scala 466:52]
  wire [7:0] _GEN_7044 = opcode_6 == 4'hf ? _GEN_6018 : _GEN_6786; // @[executor.scala 466:52]
  wire [7:0] _GEN_7045 = opcode_6 == 4'hf ? _GEN_6019 : _GEN_6787; // @[executor.scala 466:52]
  wire [7:0] _GEN_7046 = opcode_6 == 4'hf ? _GEN_6020 : _GEN_6788; // @[executor.scala 466:52]
  wire [7:0] _GEN_7047 = opcode_6 == 4'hf ? _GEN_6021 : _GEN_6789; // @[executor.scala 466:52]
  wire [7:0] _GEN_7048 = opcode_6 == 4'hf ? _GEN_6022 : _GEN_6790; // @[executor.scala 466:52]
  wire [7:0] _GEN_7049 = opcode_6 == 4'hf ? _GEN_6023 : _GEN_6791; // @[executor.scala 466:52]
  wire [7:0] _GEN_7050 = opcode_6 == 4'hf ? _GEN_6024 : _GEN_6792; // @[executor.scala 466:52]
  wire [7:0] _GEN_7051 = opcode_6 == 4'hf ? _GEN_6025 : _GEN_6793; // @[executor.scala 466:52]
  wire [7:0] _GEN_7052 = opcode_6 == 4'hf ? _GEN_6026 : _GEN_6794; // @[executor.scala 466:52]
  wire [7:0] _GEN_7053 = opcode_6 == 4'hf ? _GEN_6027 : _GEN_6795; // @[executor.scala 466:52]
  wire [7:0] _GEN_7054 = opcode_6 == 4'hf ? _GEN_6028 : _GEN_6796; // @[executor.scala 466:52]
  wire [7:0] _GEN_7055 = opcode_6 == 4'hf ? _GEN_6029 : _GEN_6797; // @[executor.scala 466:52]
  wire [7:0] _GEN_7056 = opcode_6 == 4'hf ? _GEN_6030 : _GEN_6798; // @[executor.scala 466:52]
  wire [7:0] _GEN_7057 = opcode_6 == 4'hf ? _GEN_6031 : _GEN_6799; // @[executor.scala 466:52]
  wire [7:0] _GEN_7058 = opcode_6 == 4'hf ? _GEN_6032 : _GEN_6800; // @[executor.scala 466:52]
  wire [7:0] _GEN_7059 = opcode_6 == 4'hf ? _GEN_6033 : _GEN_6801; // @[executor.scala 466:52]
  wire [7:0] _GEN_7060 = opcode_6 == 4'hf ? _GEN_6034 : _GEN_6802; // @[executor.scala 466:52]
  wire [7:0] _GEN_7061 = opcode_6 == 4'hf ? _GEN_6035 : _GEN_6803; // @[executor.scala 466:52]
  wire [7:0] _GEN_7062 = opcode_6 == 4'hf ? _GEN_6036 : _GEN_6804; // @[executor.scala 466:52]
  wire [7:0] _GEN_7063 = opcode_6 == 4'hf ? _GEN_6037 : _GEN_6805; // @[executor.scala 466:52]
  wire [7:0] _GEN_7064 = opcode_6 == 4'hf ? _GEN_6038 : _GEN_6806; // @[executor.scala 466:52]
  wire [7:0] _GEN_7065 = opcode_6 == 4'hf ? _GEN_6039 : _GEN_6807; // @[executor.scala 466:52]
  wire [7:0] _GEN_7066 = opcode_6 == 4'hf ? _GEN_6040 : _GEN_6808; // @[executor.scala 466:52]
  wire [7:0] _GEN_7067 = opcode_6 == 4'hf ? _GEN_6041 : _GEN_6809; // @[executor.scala 466:52]
  wire [7:0] _GEN_7068 = opcode_6 == 4'hf ? _GEN_6042 : _GEN_6810; // @[executor.scala 466:52]
  wire [7:0] _GEN_7069 = opcode_6 == 4'hf ? _GEN_6043 : _GEN_6811; // @[executor.scala 466:52]
  wire [7:0] _GEN_7070 = opcode_6 == 4'hf ? _GEN_6044 : _GEN_6812; // @[executor.scala 466:52]
  wire [7:0] _GEN_7071 = opcode_6 == 4'hf ? _GEN_6045 : _GEN_6813; // @[executor.scala 466:52]
  wire [7:0] _GEN_7072 = opcode_6 == 4'hf ? _GEN_6046 : _GEN_6814; // @[executor.scala 466:52]
  wire [7:0] _GEN_7073 = opcode_6 == 4'hf ? _GEN_6047 : _GEN_6815; // @[executor.scala 466:52]
  wire [7:0] _GEN_7074 = opcode_6 == 4'hf ? _GEN_6048 : _GEN_6816; // @[executor.scala 466:52]
  wire [7:0] _GEN_7075 = opcode_6 == 4'hf ? _GEN_6049 : _GEN_6817; // @[executor.scala 466:52]
  wire [7:0] _GEN_7076 = opcode_6 == 4'hf ? _GEN_6050 : _GEN_6818; // @[executor.scala 466:52]
  wire [7:0] _GEN_7077 = opcode_6 == 4'hf ? _GEN_6051 : _GEN_6819; // @[executor.scala 466:52]
  wire [7:0] _GEN_7078 = opcode_6 == 4'hf ? _GEN_6052 : _GEN_6820; // @[executor.scala 466:52]
  wire [7:0] _GEN_7079 = opcode_6 == 4'hf ? _GEN_6053 : _GEN_6821; // @[executor.scala 466:52]
  wire [7:0] _GEN_7080 = opcode_6 == 4'hf ? _GEN_6054 : _GEN_6822; // @[executor.scala 466:52]
  wire [7:0] _GEN_7081 = opcode_6 == 4'hf ? _GEN_6055 : _GEN_6823; // @[executor.scala 466:52]
  wire [7:0] _GEN_7082 = opcode_6 == 4'hf ? _GEN_6056 : _GEN_6824; // @[executor.scala 466:52]
  wire [7:0] _GEN_7083 = opcode_6 == 4'hf ? _GEN_6057 : _GEN_6825; // @[executor.scala 466:52]
  wire [7:0] _GEN_7084 = opcode_6 == 4'hf ? _GEN_6058 : _GEN_6826; // @[executor.scala 466:52]
  wire [7:0] _GEN_7085 = opcode_6 == 4'hf ? _GEN_6059 : _GEN_6827; // @[executor.scala 466:52]
  wire [7:0] _GEN_7086 = opcode_6 == 4'hf ? _GEN_6060 : _GEN_6828; // @[executor.scala 466:52]
  wire [7:0] _GEN_7087 = opcode_6 == 4'hf ? _GEN_6061 : _GEN_6829; // @[executor.scala 466:52]
  wire [7:0] _GEN_7088 = opcode_6 == 4'hf ? _GEN_6062 : _GEN_6830; // @[executor.scala 466:52]
  wire [7:0] _GEN_7089 = opcode_6 == 4'hf ? _GEN_6063 : _GEN_6831; // @[executor.scala 466:52]
  wire [7:0] _GEN_7090 = opcode_6 == 4'hf ? _GEN_6064 : _GEN_6832; // @[executor.scala 466:52]
  wire [7:0] _GEN_7091 = opcode_6 == 4'hf ? _GEN_6065 : _GEN_6833; // @[executor.scala 466:52]
  wire [7:0] _GEN_7092 = opcode_6 == 4'hf ? _GEN_6066 : _GEN_6834; // @[executor.scala 466:52]
  wire [7:0] _GEN_7093 = opcode_6 == 4'hf ? _GEN_6067 : _GEN_6835; // @[executor.scala 466:52]
  wire [7:0] _GEN_7094 = opcode_6 == 4'hf ? _GEN_6068 : _GEN_6836; // @[executor.scala 466:52]
  wire [7:0] _GEN_7095 = opcode_6 == 4'hf ? _GEN_6069 : _GEN_6837; // @[executor.scala 466:52]
  wire [7:0] _GEN_7096 = opcode_6 == 4'hf ? _GEN_6070 : _GEN_6838; // @[executor.scala 466:52]
  wire [7:0] _GEN_7097 = opcode_6 == 4'hf ? _GEN_6071 : _GEN_6839; // @[executor.scala 466:52]
  wire [7:0] _GEN_7098 = opcode_6 == 4'hf ? _GEN_6072 : _GEN_6840; // @[executor.scala 466:52]
  wire [7:0] _GEN_7099 = opcode_6 == 4'hf ? _GEN_6073 : _GEN_6841; // @[executor.scala 466:52]
  wire [7:0] _GEN_7100 = opcode_6 == 4'hf ? _GEN_6074 : _GEN_6842; // @[executor.scala 466:52]
  wire [7:0] _GEN_7101 = opcode_6 == 4'hf ? _GEN_6075 : _GEN_6843; // @[executor.scala 466:52]
  wire [7:0] _GEN_7102 = opcode_6 == 4'hf ? _GEN_6076 : _GEN_6844; // @[executor.scala 466:52]
  wire [7:0] _GEN_7103 = opcode_6 == 4'hf ? _GEN_6077 : _GEN_6845; // @[executor.scala 466:52]
  wire [7:0] _GEN_7104 = opcode_6 == 4'hf ? _GEN_6078 : _GEN_6846; // @[executor.scala 466:52]
  wire [7:0] _GEN_7105 = opcode_6 == 4'hf ? _GEN_6079 : _GEN_6847; // @[executor.scala 466:52]
  wire [7:0] _GEN_7106 = opcode_6 == 4'hf ? _GEN_6080 : _GEN_6848; // @[executor.scala 466:52]
  wire [7:0] _GEN_7107 = opcode_6 == 4'hf ? _GEN_6081 : _GEN_6849; // @[executor.scala 466:52]
  wire [7:0] _GEN_7108 = opcode_6 == 4'hf ? _GEN_6082 : _GEN_6850; // @[executor.scala 466:52]
  wire [7:0] _GEN_7109 = opcode_6 == 4'hf ? _GEN_6083 : _GEN_6851; // @[executor.scala 466:52]
  wire [7:0] _GEN_7110 = opcode_6 == 4'hf ? _GEN_6084 : _GEN_6852; // @[executor.scala 466:52]
  wire [7:0] _GEN_7111 = opcode_6 == 4'hf ? _GEN_6085 : _GEN_6853; // @[executor.scala 466:52]
  wire [7:0] _GEN_7112 = opcode_6 == 4'hf ? _GEN_6086 : _GEN_6854; // @[executor.scala 466:52]
  wire [7:0] _GEN_7113 = opcode_6 == 4'hf ? _GEN_6087 : _GEN_6855; // @[executor.scala 466:52]
  wire [7:0] _GEN_7114 = opcode_6 == 4'hf ? _GEN_6088 : _GEN_6856; // @[executor.scala 466:52]
  wire [7:0] _GEN_7115 = opcode_6 == 4'hf ? _GEN_6089 : _GEN_6857; // @[executor.scala 466:52]
  wire [7:0] _GEN_7116 = opcode_6 == 4'hf ? _GEN_6090 : _GEN_6858; // @[executor.scala 466:52]
  wire [7:0] _GEN_7117 = opcode_6 == 4'hf ? _GEN_6091 : _GEN_6859; // @[executor.scala 466:52]
  wire [7:0] _GEN_7118 = opcode_6 == 4'hf ? _GEN_6092 : _GEN_6860; // @[executor.scala 466:52]
  wire [7:0] _GEN_7119 = opcode_6 == 4'hf ? _GEN_6093 : _GEN_6861; // @[executor.scala 466:52]
  wire [7:0] _GEN_7120 = opcode_6 == 4'hf ? _GEN_6094 : _GEN_6862; // @[executor.scala 466:52]
  wire [7:0] _GEN_7121 = opcode_6 == 4'hf ? _GEN_6095 : _GEN_6863; // @[executor.scala 466:52]
  wire [7:0] _GEN_7122 = opcode_6 == 4'hf ? _GEN_6096 : _GEN_6864; // @[executor.scala 466:52]
  wire [7:0] _GEN_7123 = opcode_6 == 4'hf ? _GEN_6097 : _GEN_6865; // @[executor.scala 466:52]
  wire [7:0] _GEN_7124 = opcode_6 == 4'hf ? _GEN_6098 : _GEN_6866; // @[executor.scala 466:52]
  wire [7:0] _GEN_7125 = opcode_6 == 4'hf ? _GEN_6099 : _GEN_6867; // @[executor.scala 466:52]
  wire [7:0] _GEN_7126 = opcode_6 == 4'hf ? _GEN_6100 : _GEN_6868; // @[executor.scala 466:52]
  wire [7:0] _GEN_7127 = opcode_6 == 4'hf ? _GEN_6101 : _GEN_6869; // @[executor.scala 466:52]
  wire [7:0] _GEN_7128 = opcode_6 == 4'hf ? _GEN_6102 : _GEN_6870; // @[executor.scala 466:52]
  wire [7:0] _GEN_7129 = opcode_6 == 4'hf ? _GEN_6103 : _GEN_6871; // @[executor.scala 466:52]
  wire [7:0] _GEN_7130 = opcode_6 == 4'hf ? _GEN_6104 : _GEN_6872; // @[executor.scala 466:52]
  wire [7:0] _GEN_7131 = opcode_6 == 4'hf ? _GEN_6105 : _GEN_6873; // @[executor.scala 466:52]
  wire [7:0] _GEN_7132 = opcode_6 == 4'hf ? _GEN_6106 : _GEN_6874; // @[executor.scala 466:52]
  wire [7:0] _GEN_7133 = opcode_6 == 4'hf ? _GEN_6107 : _GEN_6875; // @[executor.scala 466:52]
  wire [7:0] _GEN_7134 = opcode_6 == 4'hf ? _GEN_6108 : _GEN_6876; // @[executor.scala 466:52]
  wire [7:0] _GEN_7135 = opcode_6 == 4'hf ? _GEN_6109 : _GEN_6877; // @[executor.scala 466:52]
  wire [7:0] _GEN_7136 = opcode_6 == 4'hf ? _GEN_6110 : _GEN_6878; // @[executor.scala 466:52]
  wire [7:0] _GEN_7137 = opcode_6 == 4'hf ? _GEN_6111 : _GEN_6879; // @[executor.scala 466:52]
  wire [7:0] _GEN_7138 = opcode_6 == 4'hf ? _GEN_6112 : _GEN_6880; // @[executor.scala 466:52]
  wire [7:0] _GEN_7139 = opcode_6 == 4'hf ? _GEN_6113 : _GEN_6881; // @[executor.scala 466:52]
  wire [7:0] _GEN_7140 = opcode_6 == 4'hf ? _GEN_6114 : _GEN_6882; // @[executor.scala 466:52]
  wire [7:0] _GEN_7141 = opcode_6 == 4'hf ? _GEN_6115 : _GEN_6883; // @[executor.scala 466:52]
  wire [7:0] _GEN_7142 = opcode_6 == 4'hf ? _GEN_6116 : _GEN_6884; // @[executor.scala 466:52]
  wire [7:0] _GEN_7143 = opcode_6 == 4'hf ? _GEN_6117 : _GEN_6885; // @[executor.scala 466:52]
  wire [7:0] _GEN_7144 = opcode_6 == 4'hf ? _GEN_6118 : _GEN_6886; // @[executor.scala 466:52]
  wire [7:0] _GEN_7145 = opcode_6 == 4'hf ? _GEN_6119 : _GEN_6887; // @[executor.scala 466:52]
  wire [7:0] _GEN_7146 = opcode_6 == 4'hf ? _GEN_6120 : _GEN_6888; // @[executor.scala 466:52]
  wire [7:0] _GEN_7147 = opcode_6 == 4'hf ? _GEN_6121 : _GEN_6889; // @[executor.scala 466:52]
  wire [7:0] _GEN_7148 = opcode_6 == 4'hf ? _GEN_6122 : _GEN_6890; // @[executor.scala 466:52]
  wire [7:0] _GEN_7149 = opcode_6 == 4'hf ? _GEN_6123 : _GEN_6891; // @[executor.scala 466:52]
  wire [7:0] _GEN_7150 = opcode_6 == 4'hf ? _GEN_6124 : _GEN_6892; // @[executor.scala 466:52]
  wire [7:0] _GEN_7151 = opcode_6 == 4'hf ? _GEN_6125 : _GEN_6893; // @[executor.scala 466:52]
  wire [7:0] _GEN_7152 = opcode_6 == 4'hf ? _GEN_6126 : _GEN_6894; // @[executor.scala 466:52]
  wire [7:0] _GEN_7153 = opcode_6 == 4'hf ? _GEN_6127 : _GEN_6895; // @[executor.scala 466:52]
  wire [7:0] _GEN_7154 = opcode_6 == 4'hf ? _GEN_6128 : _GEN_6896; // @[executor.scala 466:52]
  wire [7:0] _GEN_7155 = opcode_6 == 4'hf ? _GEN_6129 : _GEN_6897; // @[executor.scala 466:52]
  wire [7:0] _GEN_7156 = opcode_6 == 4'hf ? _GEN_6130 : _GEN_6898; // @[executor.scala 466:52]
  wire [7:0] _GEN_7157 = opcode_6 == 4'hf ? _GEN_6131 : _GEN_6899; // @[executor.scala 466:52]
  wire [7:0] _GEN_7158 = opcode_6 == 4'hf ? _GEN_6132 : _GEN_6900; // @[executor.scala 466:52]
  wire [7:0] _GEN_7159 = opcode_6 == 4'hf ? _GEN_6133 : _GEN_6901; // @[executor.scala 466:52]
  wire [7:0] _GEN_7160 = opcode_6 == 4'hf ? _GEN_6134 : _GEN_6902; // @[executor.scala 466:52]
  wire [7:0] _GEN_7161 = opcode_6 == 4'hf ? _GEN_6135 : _GEN_6903; // @[executor.scala 466:52]
  wire [7:0] _GEN_7162 = opcode_6 == 4'hf ? _GEN_6136 : _GEN_6904; // @[executor.scala 466:52]
  wire [7:0] _GEN_7163 = opcode_6 == 4'hf ? _GEN_6137 : _GEN_6905; // @[executor.scala 466:52]
  wire [7:0] _GEN_7164 = opcode_6 == 4'hf ? _GEN_6138 : _GEN_6906; // @[executor.scala 466:52]
  wire [7:0] _GEN_7165 = opcode_6 == 4'hf ? _GEN_6139 : _GEN_6907; // @[executor.scala 466:52]
  wire [7:0] _GEN_7166 = opcode_6 == 4'hf ? _GEN_6140 : _GEN_6908; // @[executor.scala 466:52]
  wire [7:0] _GEN_7167 = opcode_6 == 4'hf ? _GEN_6141 : _GEN_6909; // @[executor.scala 466:52]
  wire [7:0] _GEN_7168 = opcode_6 == 4'hf ? _GEN_6142 : _GEN_6910; // @[executor.scala 466:52]
  wire [7:0] _GEN_7169 = opcode_6 == 4'hf ? _GEN_6143 : _GEN_6911; // @[executor.scala 466:52]
  wire [7:0] _GEN_7170 = opcode_6 == 4'hf ? _GEN_6144 : _GEN_6912; // @[executor.scala 466:52]
  wire [7:0] _GEN_7171 = opcode_6 == 4'hf ? _GEN_6145 : _GEN_6913; // @[executor.scala 466:52]
  wire [7:0] _GEN_7172 = opcode_6 == 4'hf ? _GEN_6146 : _GEN_6914; // @[executor.scala 466:52]
  wire [7:0] _GEN_7173 = opcode_6 == 4'hf ? _GEN_6147 : _GEN_6915; // @[executor.scala 466:52]
  wire [7:0] _GEN_7174 = opcode_6 == 4'hf ? _GEN_6148 : _GEN_6916; // @[executor.scala 466:52]
  wire [7:0] _GEN_7175 = opcode_6 == 4'hf ? _GEN_6149 : _GEN_6917; // @[executor.scala 466:52]
  wire [7:0] _GEN_7176 = opcode_6 == 4'hf ? _GEN_6150 : _GEN_6918; // @[executor.scala 466:52]
  wire [7:0] _GEN_7177 = opcode_6 == 4'hf ? _GEN_6151 : _GEN_6919; // @[executor.scala 466:52]
  wire [7:0] _GEN_7178 = opcode_6 == 4'hf ? _GEN_6152 : _GEN_6920; // @[executor.scala 466:52]
  wire [7:0] _GEN_7179 = opcode_6 == 4'hf ? _GEN_6153 : _GEN_6921; // @[executor.scala 466:52]
  wire [7:0] _GEN_7180 = opcode_6 == 4'hf ? _GEN_6154 : _GEN_6922; // @[executor.scala 466:52]
  wire [7:0] _GEN_7181 = opcode_6 == 4'hf ? _GEN_6155 : _GEN_6923; // @[executor.scala 466:52]
  wire [3:0] opcode_7 = vliw_7[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_7 = vliw_7[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8914 = {{2'd0}, dst_offset_7}; // @[executor.scala 473:49]
  wire [7:0] byte_1792 = field_7[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_7182 = mask_7[0] ? byte_1792 : _GEN_6926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1793 = field_7[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_7183 = mask_7[1] ? byte_1793 : _GEN_6927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1794 = field_7[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_7184 = mask_7[2] ? byte_1794 : _GEN_6928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1795 = field_7[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_7185 = mask_7[3] ? byte_1795 : _GEN_6929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7186 = _GEN_8914 == 8'h0 ? _GEN_7182 : _GEN_6926; // @[executor.scala 473:84]
  wire [7:0] _GEN_7187 = _GEN_8914 == 8'h0 ? _GEN_7183 : _GEN_6927; // @[executor.scala 473:84]
  wire [7:0] _GEN_7188 = _GEN_8914 == 8'h0 ? _GEN_7184 : _GEN_6928; // @[executor.scala 473:84]
  wire [7:0] _GEN_7189 = _GEN_8914 == 8'h0 ? _GEN_7185 : _GEN_6929; // @[executor.scala 473:84]
  wire [7:0] _GEN_7190 = mask_7[0] ? byte_1792 : _GEN_6930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7191 = mask_7[1] ? byte_1793 : _GEN_6931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7192 = mask_7[2] ? byte_1794 : _GEN_6932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7193 = mask_7[3] ? byte_1795 : _GEN_6933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7194 = _GEN_8914 == 8'h1 ? _GEN_7190 : _GEN_6930; // @[executor.scala 473:84]
  wire [7:0] _GEN_7195 = _GEN_8914 == 8'h1 ? _GEN_7191 : _GEN_6931; // @[executor.scala 473:84]
  wire [7:0] _GEN_7196 = _GEN_8914 == 8'h1 ? _GEN_7192 : _GEN_6932; // @[executor.scala 473:84]
  wire [7:0] _GEN_7197 = _GEN_8914 == 8'h1 ? _GEN_7193 : _GEN_6933; // @[executor.scala 473:84]
  wire [7:0] _GEN_7198 = mask_7[0] ? byte_1792 : _GEN_6934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7199 = mask_7[1] ? byte_1793 : _GEN_6935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7200 = mask_7[2] ? byte_1794 : _GEN_6936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7201 = mask_7[3] ? byte_1795 : _GEN_6937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7202 = _GEN_8914 == 8'h2 ? _GEN_7198 : _GEN_6934; // @[executor.scala 473:84]
  wire [7:0] _GEN_7203 = _GEN_8914 == 8'h2 ? _GEN_7199 : _GEN_6935; // @[executor.scala 473:84]
  wire [7:0] _GEN_7204 = _GEN_8914 == 8'h2 ? _GEN_7200 : _GEN_6936; // @[executor.scala 473:84]
  wire [7:0] _GEN_7205 = _GEN_8914 == 8'h2 ? _GEN_7201 : _GEN_6937; // @[executor.scala 473:84]
  wire [7:0] _GEN_7206 = mask_7[0] ? byte_1792 : _GEN_6938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7207 = mask_7[1] ? byte_1793 : _GEN_6939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7208 = mask_7[2] ? byte_1794 : _GEN_6940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7209 = mask_7[3] ? byte_1795 : _GEN_6941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7210 = _GEN_8914 == 8'h3 ? _GEN_7206 : _GEN_6938; // @[executor.scala 473:84]
  wire [7:0] _GEN_7211 = _GEN_8914 == 8'h3 ? _GEN_7207 : _GEN_6939; // @[executor.scala 473:84]
  wire [7:0] _GEN_7212 = _GEN_8914 == 8'h3 ? _GEN_7208 : _GEN_6940; // @[executor.scala 473:84]
  wire [7:0] _GEN_7213 = _GEN_8914 == 8'h3 ? _GEN_7209 : _GEN_6941; // @[executor.scala 473:84]
  wire [7:0] _GEN_7214 = mask_7[0] ? byte_1792 : _GEN_6942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7215 = mask_7[1] ? byte_1793 : _GEN_6943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7216 = mask_7[2] ? byte_1794 : _GEN_6944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7217 = mask_7[3] ? byte_1795 : _GEN_6945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7218 = _GEN_8914 == 8'h4 ? _GEN_7214 : _GEN_6942; // @[executor.scala 473:84]
  wire [7:0] _GEN_7219 = _GEN_8914 == 8'h4 ? _GEN_7215 : _GEN_6943; // @[executor.scala 473:84]
  wire [7:0] _GEN_7220 = _GEN_8914 == 8'h4 ? _GEN_7216 : _GEN_6944; // @[executor.scala 473:84]
  wire [7:0] _GEN_7221 = _GEN_8914 == 8'h4 ? _GEN_7217 : _GEN_6945; // @[executor.scala 473:84]
  wire [7:0] _GEN_7222 = mask_7[0] ? byte_1792 : _GEN_6946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7223 = mask_7[1] ? byte_1793 : _GEN_6947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7224 = mask_7[2] ? byte_1794 : _GEN_6948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7225 = mask_7[3] ? byte_1795 : _GEN_6949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7226 = _GEN_8914 == 8'h5 ? _GEN_7222 : _GEN_6946; // @[executor.scala 473:84]
  wire [7:0] _GEN_7227 = _GEN_8914 == 8'h5 ? _GEN_7223 : _GEN_6947; // @[executor.scala 473:84]
  wire [7:0] _GEN_7228 = _GEN_8914 == 8'h5 ? _GEN_7224 : _GEN_6948; // @[executor.scala 473:84]
  wire [7:0] _GEN_7229 = _GEN_8914 == 8'h5 ? _GEN_7225 : _GEN_6949; // @[executor.scala 473:84]
  wire [7:0] _GEN_7230 = mask_7[0] ? byte_1792 : _GEN_6950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7231 = mask_7[1] ? byte_1793 : _GEN_6951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7232 = mask_7[2] ? byte_1794 : _GEN_6952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7233 = mask_7[3] ? byte_1795 : _GEN_6953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7234 = _GEN_8914 == 8'h6 ? _GEN_7230 : _GEN_6950; // @[executor.scala 473:84]
  wire [7:0] _GEN_7235 = _GEN_8914 == 8'h6 ? _GEN_7231 : _GEN_6951; // @[executor.scala 473:84]
  wire [7:0] _GEN_7236 = _GEN_8914 == 8'h6 ? _GEN_7232 : _GEN_6952; // @[executor.scala 473:84]
  wire [7:0] _GEN_7237 = _GEN_8914 == 8'h6 ? _GEN_7233 : _GEN_6953; // @[executor.scala 473:84]
  wire [7:0] _GEN_7238 = mask_7[0] ? byte_1792 : _GEN_6954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7239 = mask_7[1] ? byte_1793 : _GEN_6955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7240 = mask_7[2] ? byte_1794 : _GEN_6956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7241 = mask_7[3] ? byte_1795 : _GEN_6957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7242 = _GEN_8914 == 8'h7 ? _GEN_7238 : _GEN_6954; // @[executor.scala 473:84]
  wire [7:0] _GEN_7243 = _GEN_8914 == 8'h7 ? _GEN_7239 : _GEN_6955; // @[executor.scala 473:84]
  wire [7:0] _GEN_7244 = _GEN_8914 == 8'h7 ? _GEN_7240 : _GEN_6956; // @[executor.scala 473:84]
  wire [7:0] _GEN_7245 = _GEN_8914 == 8'h7 ? _GEN_7241 : _GEN_6957; // @[executor.scala 473:84]
  wire [7:0] _GEN_7246 = mask_7[0] ? byte_1792 : _GEN_6958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7247 = mask_7[1] ? byte_1793 : _GEN_6959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7248 = mask_7[2] ? byte_1794 : _GEN_6960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7249 = mask_7[3] ? byte_1795 : _GEN_6961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7250 = _GEN_8914 == 8'h8 ? _GEN_7246 : _GEN_6958; // @[executor.scala 473:84]
  wire [7:0] _GEN_7251 = _GEN_8914 == 8'h8 ? _GEN_7247 : _GEN_6959; // @[executor.scala 473:84]
  wire [7:0] _GEN_7252 = _GEN_8914 == 8'h8 ? _GEN_7248 : _GEN_6960; // @[executor.scala 473:84]
  wire [7:0] _GEN_7253 = _GEN_8914 == 8'h8 ? _GEN_7249 : _GEN_6961; // @[executor.scala 473:84]
  wire [7:0] _GEN_7254 = mask_7[0] ? byte_1792 : _GEN_6962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7255 = mask_7[1] ? byte_1793 : _GEN_6963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7256 = mask_7[2] ? byte_1794 : _GEN_6964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7257 = mask_7[3] ? byte_1795 : _GEN_6965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7258 = _GEN_8914 == 8'h9 ? _GEN_7254 : _GEN_6962; // @[executor.scala 473:84]
  wire [7:0] _GEN_7259 = _GEN_8914 == 8'h9 ? _GEN_7255 : _GEN_6963; // @[executor.scala 473:84]
  wire [7:0] _GEN_7260 = _GEN_8914 == 8'h9 ? _GEN_7256 : _GEN_6964; // @[executor.scala 473:84]
  wire [7:0] _GEN_7261 = _GEN_8914 == 8'h9 ? _GEN_7257 : _GEN_6965; // @[executor.scala 473:84]
  wire [7:0] _GEN_7262 = mask_7[0] ? byte_1792 : _GEN_6966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7263 = mask_7[1] ? byte_1793 : _GEN_6967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7264 = mask_7[2] ? byte_1794 : _GEN_6968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7265 = mask_7[3] ? byte_1795 : _GEN_6969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7266 = _GEN_8914 == 8'ha ? _GEN_7262 : _GEN_6966; // @[executor.scala 473:84]
  wire [7:0] _GEN_7267 = _GEN_8914 == 8'ha ? _GEN_7263 : _GEN_6967; // @[executor.scala 473:84]
  wire [7:0] _GEN_7268 = _GEN_8914 == 8'ha ? _GEN_7264 : _GEN_6968; // @[executor.scala 473:84]
  wire [7:0] _GEN_7269 = _GEN_8914 == 8'ha ? _GEN_7265 : _GEN_6969; // @[executor.scala 473:84]
  wire [7:0] _GEN_7270 = mask_7[0] ? byte_1792 : _GEN_6970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7271 = mask_7[1] ? byte_1793 : _GEN_6971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7272 = mask_7[2] ? byte_1794 : _GEN_6972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7273 = mask_7[3] ? byte_1795 : _GEN_6973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7274 = _GEN_8914 == 8'hb ? _GEN_7270 : _GEN_6970; // @[executor.scala 473:84]
  wire [7:0] _GEN_7275 = _GEN_8914 == 8'hb ? _GEN_7271 : _GEN_6971; // @[executor.scala 473:84]
  wire [7:0] _GEN_7276 = _GEN_8914 == 8'hb ? _GEN_7272 : _GEN_6972; // @[executor.scala 473:84]
  wire [7:0] _GEN_7277 = _GEN_8914 == 8'hb ? _GEN_7273 : _GEN_6973; // @[executor.scala 473:84]
  wire [7:0] _GEN_7278 = mask_7[0] ? byte_1792 : _GEN_6974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7279 = mask_7[1] ? byte_1793 : _GEN_6975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7280 = mask_7[2] ? byte_1794 : _GEN_6976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7281 = mask_7[3] ? byte_1795 : _GEN_6977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7282 = _GEN_8914 == 8'hc ? _GEN_7278 : _GEN_6974; // @[executor.scala 473:84]
  wire [7:0] _GEN_7283 = _GEN_8914 == 8'hc ? _GEN_7279 : _GEN_6975; // @[executor.scala 473:84]
  wire [7:0] _GEN_7284 = _GEN_8914 == 8'hc ? _GEN_7280 : _GEN_6976; // @[executor.scala 473:84]
  wire [7:0] _GEN_7285 = _GEN_8914 == 8'hc ? _GEN_7281 : _GEN_6977; // @[executor.scala 473:84]
  wire [7:0] _GEN_7286 = mask_7[0] ? byte_1792 : _GEN_6978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7287 = mask_7[1] ? byte_1793 : _GEN_6979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7288 = mask_7[2] ? byte_1794 : _GEN_6980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7289 = mask_7[3] ? byte_1795 : _GEN_6981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7290 = _GEN_8914 == 8'hd ? _GEN_7286 : _GEN_6978; // @[executor.scala 473:84]
  wire [7:0] _GEN_7291 = _GEN_8914 == 8'hd ? _GEN_7287 : _GEN_6979; // @[executor.scala 473:84]
  wire [7:0] _GEN_7292 = _GEN_8914 == 8'hd ? _GEN_7288 : _GEN_6980; // @[executor.scala 473:84]
  wire [7:0] _GEN_7293 = _GEN_8914 == 8'hd ? _GEN_7289 : _GEN_6981; // @[executor.scala 473:84]
  wire [7:0] _GEN_7294 = mask_7[0] ? byte_1792 : _GEN_6982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7295 = mask_7[1] ? byte_1793 : _GEN_6983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7296 = mask_7[2] ? byte_1794 : _GEN_6984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7297 = mask_7[3] ? byte_1795 : _GEN_6985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7298 = _GEN_8914 == 8'he ? _GEN_7294 : _GEN_6982; // @[executor.scala 473:84]
  wire [7:0] _GEN_7299 = _GEN_8914 == 8'he ? _GEN_7295 : _GEN_6983; // @[executor.scala 473:84]
  wire [7:0] _GEN_7300 = _GEN_8914 == 8'he ? _GEN_7296 : _GEN_6984; // @[executor.scala 473:84]
  wire [7:0] _GEN_7301 = _GEN_8914 == 8'he ? _GEN_7297 : _GEN_6985; // @[executor.scala 473:84]
  wire [7:0] _GEN_7302 = mask_7[0] ? byte_1792 : _GEN_6986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7303 = mask_7[1] ? byte_1793 : _GEN_6987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7304 = mask_7[2] ? byte_1794 : _GEN_6988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7305 = mask_7[3] ? byte_1795 : _GEN_6989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7306 = _GEN_8914 == 8'hf ? _GEN_7302 : _GEN_6986; // @[executor.scala 473:84]
  wire [7:0] _GEN_7307 = _GEN_8914 == 8'hf ? _GEN_7303 : _GEN_6987; // @[executor.scala 473:84]
  wire [7:0] _GEN_7308 = _GEN_8914 == 8'hf ? _GEN_7304 : _GEN_6988; // @[executor.scala 473:84]
  wire [7:0] _GEN_7309 = _GEN_8914 == 8'hf ? _GEN_7305 : _GEN_6989; // @[executor.scala 473:84]
  wire [7:0] _GEN_7310 = mask_7[0] ? byte_1792 : _GEN_6990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7311 = mask_7[1] ? byte_1793 : _GEN_6991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7312 = mask_7[2] ? byte_1794 : _GEN_6992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7313 = mask_7[3] ? byte_1795 : _GEN_6993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7314 = _GEN_8914 == 8'h10 ? _GEN_7310 : _GEN_6990; // @[executor.scala 473:84]
  wire [7:0] _GEN_7315 = _GEN_8914 == 8'h10 ? _GEN_7311 : _GEN_6991; // @[executor.scala 473:84]
  wire [7:0] _GEN_7316 = _GEN_8914 == 8'h10 ? _GEN_7312 : _GEN_6992; // @[executor.scala 473:84]
  wire [7:0] _GEN_7317 = _GEN_8914 == 8'h10 ? _GEN_7313 : _GEN_6993; // @[executor.scala 473:84]
  wire [7:0] _GEN_7318 = mask_7[0] ? byte_1792 : _GEN_6994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7319 = mask_7[1] ? byte_1793 : _GEN_6995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7320 = mask_7[2] ? byte_1794 : _GEN_6996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7321 = mask_7[3] ? byte_1795 : _GEN_6997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7322 = _GEN_8914 == 8'h11 ? _GEN_7318 : _GEN_6994; // @[executor.scala 473:84]
  wire [7:0] _GEN_7323 = _GEN_8914 == 8'h11 ? _GEN_7319 : _GEN_6995; // @[executor.scala 473:84]
  wire [7:0] _GEN_7324 = _GEN_8914 == 8'h11 ? _GEN_7320 : _GEN_6996; // @[executor.scala 473:84]
  wire [7:0] _GEN_7325 = _GEN_8914 == 8'h11 ? _GEN_7321 : _GEN_6997; // @[executor.scala 473:84]
  wire [7:0] _GEN_7326 = mask_7[0] ? byte_1792 : _GEN_6998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7327 = mask_7[1] ? byte_1793 : _GEN_6999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7328 = mask_7[2] ? byte_1794 : _GEN_7000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7329 = mask_7[3] ? byte_1795 : _GEN_7001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7330 = _GEN_8914 == 8'h12 ? _GEN_7326 : _GEN_6998; // @[executor.scala 473:84]
  wire [7:0] _GEN_7331 = _GEN_8914 == 8'h12 ? _GEN_7327 : _GEN_6999; // @[executor.scala 473:84]
  wire [7:0] _GEN_7332 = _GEN_8914 == 8'h12 ? _GEN_7328 : _GEN_7000; // @[executor.scala 473:84]
  wire [7:0] _GEN_7333 = _GEN_8914 == 8'h12 ? _GEN_7329 : _GEN_7001; // @[executor.scala 473:84]
  wire [7:0] _GEN_7334 = mask_7[0] ? byte_1792 : _GEN_7002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7335 = mask_7[1] ? byte_1793 : _GEN_7003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7336 = mask_7[2] ? byte_1794 : _GEN_7004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7337 = mask_7[3] ? byte_1795 : _GEN_7005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7338 = _GEN_8914 == 8'h13 ? _GEN_7334 : _GEN_7002; // @[executor.scala 473:84]
  wire [7:0] _GEN_7339 = _GEN_8914 == 8'h13 ? _GEN_7335 : _GEN_7003; // @[executor.scala 473:84]
  wire [7:0] _GEN_7340 = _GEN_8914 == 8'h13 ? _GEN_7336 : _GEN_7004; // @[executor.scala 473:84]
  wire [7:0] _GEN_7341 = _GEN_8914 == 8'h13 ? _GEN_7337 : _GEN_7005; // @[executor.scala 473:84]
  wire [7:0] _GEN_7342 = mask_7[0] ? byte_1792 : _GEN_7006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7343 = mask_7[1] ? byte_1793 : _GEN_7007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7344 = mask_7[2] ? byte_1794 : _GEN_7008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7345 = mask_7[3] ? byte_1795 : _GEN_7009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7346 = _GEN_8914 == 8'h14 ? _GEN_7342 : _GEN_7006; // @[executor.scala 473:84]
  wire [7:0] _GEN_7347 = _GEN_8914 == 8'h14 ? _GEN_7343 : _GEN_7007; // @[executor.scala 473:84]
  wire [7:0] _GEN_7348 = _GEN_8914 == 8'h14 ? _GEN_7344 : _GEN_7008; // @[executor.scala 473:84]
  wire [7:0] _GEN_7349 = _GEN_8914 == 8'h14 ? _GEN_7345 : _GEN_7009; // @[executor.scala 473:84]
  wire [7:0] _GEN_7350 = mask_7[0] ? byte_1792 : _GEN_7010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7351 = mask_7[1] ? byte_1793 : _GEN_7011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7352 = mask_7[2] ? byte_1794 : _GEN_7012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7353 = mask_7[3] ? byte_1795 : _GEN_7013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7354 = _GEN_8914 == 8'h15 ? _GEN_7350 : _GEN_7010; // @[executor.scala 473:84]
  wire [7:0] _GEN_7355 = _GEN_8914 == 8'h15 ? _GEN_7351 : _GEN_7011; // @[executor.scala 473:84]
  wire [7:0] _GEN_7356 = _GEN_8914 == 8'h15 ? _GEN_7352 : _GEN_7012; // @[executor.scala 473:84]
  wire [7:0] _GEN_7357 = _GEN_8914 == 8'h15 ? _GEN_7353 : _GEN_7013; // @[executor.scala 473:84]
  wire [7:0] _GEN_7358 = mask_7[0] ? byte_1792 : _GEN_7014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7359 = mask_7[1] ? byte_1793 : _GEN_7015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7360 = mask_7[2] ? byte_1794 : _GEN_7016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7361 = mask_7[3] ? byte_1795 : _GEN_7017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7362 = _GEN_8914 == 8'h16 ? _GEN_7358 : _GEN_7014; // @[executor.scala 473:84]
  wire [7:0] _GEN_7363 = _GEN_8914 == 8'h16 ? _GEN_7359 : _GEN_7015; // @[executor.scala 473:84]
  wire [7:0] _GEN_7364 = _GEN_8914 == 8'h16 ? _GEN_7360 : _GEN_7016; // @[executor.scala 473:84]
  wire [7:0] _GEN_7365 = _GEN_8914 == 8'h16 ? _GEN_7361 : _GEN_7017; // @[executor.scala 473:84]
  wire [7:0] _GEN_7366 = mask_7[0] ? byte_1792 : _GEN_7018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7367 = mask_7[1] ? byte_1793 : _GEN_7019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7368 = mask_7[2] ? byte_1794 : _GEN_7020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7369 = mask_7[3] ? byte_1795 : _GEN_7021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7370 = _GEN_8914 == 8'h17 ? _GEN_7366 : _GEN_7018; // @[executor.scala 473:84]
  wire [7:0] _GEN_7371 = _GEN_8914 == 8'h17 ? _GEN_7367 : _GEN_7019; // @[executor.scala 473:84]
  wire [7:0] _GEN_7372 = _GEN_8914 == 8'h17 ? _GEN_7368 : _GEN_7020; // @[executor.scala 473:84]
  wire [7:0] _GEN_7373 = _GEN_8914 == 8'h17 ? _GEN_7369 : _GEN_7021; // @[executor.scala 473:84]
  wire [7:0] _GEN_7374 = mask_7[0] ? byte_1792 : _GEN_7022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7375 = mask_7[1] ? byte_1793 : _GEN_7023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7376 = mask_7[2] ? byte_1794 : _GEN_7024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7377 = mask_7[3] ? byte_1795 : _GEN_7025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7378 = _GEN_8914 == 8'h18 ? _GEN_7374 : _GEN_7022; // @[executor.scala 473:84]
  wire [7:0] _GEN_7379 = _GEN_8914 == 8'h18 ? _GEN_7375 : _GEN_7023; // @[executor.scala 473:84]
  wire [7:0] _GEN_7380 = _GEN_8914 == 8'h18 ? _GEN_7376 : _GEN_7024; // @[executor.scala 473:84]
  wire [7:0] _GEN_7381 = _GEN_8914 == 8'h18 ? _GEN_7377 : _GEN_7025; // @[executor.scala 473:84]
  wire [7:0] _GEN_7382 = mask_7[0] ? byte_1792 : _GEN_7026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7383 = mask_7[1] ? byte_1793 : _GEN_7027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7384 = mask_7[2] ? byte_1794 : _GEN_7028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7385 = mask_7[3] ? byte_1795 : _GEN_7029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7386 = _GEN_8914 == 8'h19 ? _GEN_7382 : _GEN_7026; // @[executor.scala 473:84]
  wire [7:0] _GEN_7387 = _GEN_8914 == 8'h19 ? _GEN_7383 : _GEN_7027; // @[executor.scala 473:84]
  wire [7:0] _GEN_7388 = _GEN_8914 == 8'h19 ? _GEN_7384 : _GEN_7028; // @[executor.scala 473:84]
  wire [7:0] _GEN_7389 = _GEN_8914 == 8'h19 ? _GEN_7385 : _GEN_7029; // @[executor.scala 473:84]
  wire [7:0] _GEN_7390 = mask_7[0] ? byte_1792 : _GEN_7030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7391 = mask_7[1] ? byte_1793 : _GEN_7031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7392 = mask_7[2] ? byte_1794 : _GEN_7032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7393 = mask_7[3] ? byte_1795 : _GEN_7033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7394 = _GEN_8914 == 8'h1a ? _GEN_7390 : _GEN_7030; // @[executor.scala 473:84]
  wire [7:0] _GEN_7395 = _GEN_8914 == 8'h1a ? _GEN_7391 : _GEN_7031; // @[executor.scala 473:84]
  wire [7:0] _GEN_7396 = _GEN_8914 == 8'h1a ? _GEN_7392 : _GEN_7032; // @[executor.scala 473:84]
  wire [7:0] _GEN_7397 = _GEN_8914 == 8'h1a ? _GEN_7393 : _GEN_7033; // @[executor.scala 473:84]
  wire [7:0] _GEN_7398 = mask_7[0] ? byte_1792 : _GEN_7034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7399 = mask_7[1] ? byte_1793 : _GEN_7035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7400 = mask_7[2] ? byte_1794 : _GEN_7036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7401 = mask_7[3] ? byte_1795 : _GEN_7037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7402 = _GEN_8914 == 8'h1b ? _GEN_7398 : _GEN_7034; // @[executor.scala 473:84]
  wire [7:0] _GEN_7403 = _GEN_8914 == 8'h1b ? _GEN_7399 : _GEN_7035; // @[executor.scala 473:84]
  wire [7:0] _GEN_7404 = _GEN_8914 == 8'h1b ? _GEN_7400 : _GEN_7036; // @[executor.scala 473:84]
  wire [7:0] _GEN_7405 = _GEN_8914 == 8'h1b ? _GEN_7401 : _GEN_7037; // @[executor.scala 473:84]
  wire [7:0] _GEN_7406 = mask_7[0] ? byte_1792 : _GEN_7038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7407 = mask_7[1] ? byte_1793 : _GEN_7039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7408 = mask_7[2] ? byte_1794 : _GEN_7040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7409 = mask_7[3] ? byte_1795 : _GEN_7041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7410 = _GEN_8914 == 8'h1c ? _GEN_7406 : _GEN_7038; // @[executor.scala 473:84]
  wire [7:0] _GEN_7411 = _GEN_8914 == 8'h1c ? _GEN_7407 : _GEN_7039; // @[executor.scala 473:84]
  wire [7:0] _GEN_7412 = _GEN_8914 == 8'h1c ? _GEN_7408 : _GEN_7040; // @[executor.scala 473:84]
  wire [7:0] _GEN_7413 = _GEN_8914 == 8'h1c ? _GEN_7409 : _GEN_7041; // @[executor.scala 473:84]
  wire [7:0] _GEN_7414 = mask_7[0] ? byte_1792 : _GEN_7042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7415 = mask_7[1] ? byte_1793 : _GEN_7043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7416 = mask_7[2] ? byte_1794 : _GEN_7044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7417 = mask_7[3] ? byte_1795 : _GEN_7045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7418 = _GEN_8914 == 8'h1d ? _GEN_7414 : _GEN_7042; // @[executor.scala 473:84]
  wire [7:0] _GEN_7419 = _GEN_8914 == 8'h1d ? _GEN_7415 : _GEN_7043; // @[executor.scala 473:84]
  wire [7:0] _GEN_7420 = _GEN_8914 == 8'h1d ? _GEN_7416 : _GEN_7044; // @[executor.scala 473:84]
  wire [7:0] _GEN_7421 = _GEN_8914 == 8'h1d ? _GEN_7417 : _GEN_7045; // @[executor.scala 473:84]
  wire [7:0] _GEN_7422 = mask_7[0] ? byte_1792 : _GEN_7046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7423 = mask_7[1] ? byte_1793 : _GEN_7047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7424 = mask_7[2] ? byte_1794 : _GEN_7048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7425 = mask_7[3] ? byte_1795 : _GEN_7049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7426 = _GEN_8914 == 8'h1e ? _GEN_7422 : _GEN_7046; // @[executor.scala 473:84]
  wire [7:0] _GEN_7427 = _GEN_8914 == 8'h1e ? _GEN_7423 : _GEN_7047; // @[executor.scala 473:84]
  wire [7:0] _GEN_7428 = _GEN_8914 == 8'h1e ? _GEN_7424 : _GEN_7048; // @[executor.scala 473:84]
  wire [7:0] _GEN_7429 = _GEN_8914 == 8'h1e ? _GEN_7425 : _GEN_7049; // @[executor.scala 473:84]
  wire [7:0] _GEN_7430 = mask_7[0] ? byte_1792 : _GEN_7050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7431 = mask_7[1] ? byte_1793 : _GEN_7051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7432 = mask_7[2] ? byte_1794 : _GEN_7052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7433 = mask_7[3] ? byte_1795 : _GEN_7053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7434 = _GEN_8914 == 8'h1f ? _GEN_7430 : _GEN_7050; // @[executor.scala 473:84]
  wire [7:0] _GEN_7435 = _GEN_8914 == 8'h1f ? _GEN_7431 : _GEN_7051; // @[executor.scala 473:84]
  wire [7:0] _GEN_7436 = _GEN_8914 == 8'h1f ? _GEN_7432 : _GEN_7052; // @[executor.scala 473:84]
  wire [7:0] _GEN_7437 = _GEN_8914 == 8'h1f ? _GEN_7433 : _GEN_7053; // @[executor.scala 473:84]
  wire [7:0] _GEN_7438 = mask_7[0] ? byte_1792 : _GEN_7054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7439 = mask_7[1] ? byte_1793 : _GEN_7055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7440 = mask_7[2] ? byte_1794 : _GEN_7056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7441 = mask_7[3] ? byte_1795 : _GEN_7057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7442 = _GEN_8914 == 8'h20 ? _GEN_7438 : _GEN_7054; // @[executor.scala 473:84]
  wire [7:0] _GEN_7443 = _GEN_8914 == 8'h20 ? _GEN_7439 : _GEN_7055; // @[executor.scala 473:84]
  wire [7:0] _GEN_7444 = _GEN_8914 == 8'h20 ? _GEN_7440 : _GEN_7056; // @[executor.scala 473:84]
  wire [7:0] _GEN_7445 = _GEN_8914 == 8'h20 ? _GEN_7441 : _GEN_7057; // @[executor.scala 473:84]
  wire [7:0] _GEN_7446 = mask_7[0] ? byte_1792 : _GEN_7058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7447 = mask_7[1] ? byte_1793 : _GEN_7059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7448 = mask_7[2] ? byte_1794 : _GEN_7060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7449 = mask_7[3] ? byte_1795 : _GEN_7061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7450 = _GEN_8914 == 8'h21 ? _GEN_7446 : _GEN_7058; // @[executor.scala 473:84]
  wire [7:0] _GEN_7451 = _GEN_8914 == 8'h21 ? _GEN_7447 : _GEN_7059; // @[executor.scala 473:84]
  wire [7:0] _GEN_7452 = _GEN_8914 == 8'h21 ? _GEN_7448 : _GEN_7060; // @[executor.scala 473:84]
  wire [7:0] _GEN_7453 = _GEN_8914 == 8'h21 ? _GEN_7449 : _GEN_7061; // @[executor.scala 473:84]
  wire [7:0] _GEN_7454 = mask_7[0] ? byte_1792 : _GEN_7062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7455 = mask_7[1] ? byte_1793 : _GEN_7063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7456 = mask_7[2] ? byte_1794 : _GEN_7064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7457 = mask_7[3] ? byte_1795 : _GEN_7065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7458 = _GEN_8914 == 8'h22 ? _GEN_7454 : _GEN_7062; // @[executor.scala 473:84]
  wire [7:0] _GEN_7459 = _GEN_8914 == 8'h22 ? _GEN_7455 : _GEN_7063; // @[executor.scala 473:84]
  wire [7:0] _GEN_7460 = _GEN_8914 == 8'h22 ? _GEN_7456 : _GEN_7064; // @[executor.scala 473:84]
  wire [7:0] _GEN_7461 = _GEN_8914 == 8'h22 ? _GEN_7457 : _GEN_7065; // @[executor.scala 473:84]
  wire [7:0] _GEN_7462 = mask_7[0] ? byte_1792 : _GEN_7066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7463 = mask_7[1] ? byte_1793 : _GEN_7067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7464 = mask_7[2] ? byte_1794 : _GEN_7068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7465 = mask_7[3] ? byte_1795 : _GEN_7069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7466 = _GEN_8914 == 8'h23 ? _GEN_7462 : _GEN_7066; // @[executor.scala 473:84]
  wire [7:0] _GEN_7467 = _GEN_8914 == 8'h23 ? _GEN_7463 : _GEN_7067; // @[executor.scala 473:84]
  wire [7:0] _GEN_7468 = _GEN_8914 == 8'h23 ? _GEN_7464 : _GEN_7068; // @[executor.scala 473:84]
  wire [7:0] _GEN_7469 = _GEN_8914 == 8'h23 ? _GEN_7465 : _GEN_7069; // @[executor.scala 473:84]
  wire [7:0] _GEN_7470 = mask_7[0] ? byte_1792 : _GEN_7070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7471 = mask_7[1] ? byte_1793 : _GEN_7071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7472 = mask_7[2] ? byte_1794 : _GEN_7072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7473 = mask_7[3] ? byte_1795 : _GEN_7073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7474 = _GEN_8914 == 8'h24 ? _GEN_7470 : _GEN_7070; // @[executor.scala 473:84]
  wire [7:0] _GEN_7475 = _GEN_8914 == 8'h24 ? _GEN_7471 : _GEN_7071; // @[executor.scala 473:84]
  wire [7:0] _GEN_7476 = _GEN_8914 == 8'h24 ? _GEN_7472 : _GEN_7072; // @[executor.scala 473:84]
  wire [7:0] _GEN_7477 = _GEN_8914 == 8'h24 ? _GEN_7473 : _GEN_7073; // @[executor.scala 473:84]
  wire [7:0] _GEN_7478 = mask_7[0] ? byte_1792 : _GEN_7074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7479 = mask_7[1] ? byte_1793 : _GEN_7075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7480 = mask_7[2] ? byte_1794 : _GEN_7076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7481 = mask_7[3] ? byte_1795 : _GEN_7077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7482 = _GEN_8914 == 8'h25 ? _GEN_7478 : _GEN_7074; // @[executor.scala 473:84]
  wire [7:0] _GEN_7483 = _GEN_8914 == 8'h25 ? _GEN_7479 : _GEN_7075; // @[executor.scala 473:84]
  wire [7:0] _GEN_7484 = _GEN_8914 == 8'h25 ? _GEN_7480 : _GEN_7076; // @[executor.scala 473:84]
  wire [7:0] _GEN_7485 = _GEN_8914 == 8'h25 ? _GEN_7481 : _GEN_7077; // @[executor.scala 473:84]
  wire [7:0] _GEN_7486 = mask_7[0] ? byte_1792 : _GEN_7078; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7487 = mask_7[1] ? byte_1793 : _GEN_7079; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7488 = mask_7[2] ? byte_1794 : _GEN_7080; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7489 = mask_7[3] ? byte_1795 : _GEN_7081; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7490 = _GEN_8914 == 8'h26 ? _GEN_7486 : _GEN_7078; // @[executor.scala 473:84]
  wire [7:0] _GEN_7491 = _GEN_8914 == 8'h26 ? _GEN_7487 : _GEN_7079; // @[executor.scala 473:84]
  wire [7:0] _GEN_7492 = _GEN_8914 == 8'h26 ? _GEN_7488 : _GEN_7080; // @[executor.scala 473:84]
  wire [7:0] _GEN_7493 = _GEN_8914 == 8'h26 ? _GEN_7489 : _GEN_7081; // @[executor.scala 473:84]
  wire [7:0] _GEN_7494 = mask_7[0] ? byte_1792 : _GEN_7082; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7495 = mask_7[1] ? byte_1793 : _GEN_7083; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7496 = mask_7[2] ? byte_1794 : _GEN_7084; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7497 = mask_7[3] ? byte_1795 : _GEN_7085; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7498 = _GEN_8914 == 8'h27 ? _GEN_7494 : _GEN_7082; // @[executor.scala 473:84]
  wire [7:0] _GEN_7499 = _GEN_8914 == 8'h27 ? _GEN_7495 : _GEN_7083; // @[executor.scala 473:84]
  wire [7:0] _GEN_7500 = _GEN_8914 == 8'h27 ? _GEN_7496 : _GEN_7084; // @[executor.scala 473:84]
  wire [7:0] _GEN_7501 = _GEN_8914 == 8'h27 ? _GEN_7497 : _GEN_7085; // @[executor.scala 473:84]
  wire [7:0] _GEN_7502 = mask_7[0] ? byte_1792 : _GEN_7086; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7503 = mask_7[1] ? byte_1793 : _GEN_7087; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7504 = mask_7[2] ? byte_1794 : _GEN_7088; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7505 = mask_7[3] ? byte_1795 : _GEN_7089; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7506 = _GEN_8914 == 8'h28 ? _GEN_7502 : _GEN_7086; // @[executor.scala 473:84]
  wire [7:0] _GEN_7507 = _GEN_8914 == 8'h28 ? _GEN_7503 : _GEN_7087; // @[executor.scala 473:84]
  wire [7:0] _GEN_7508 = _GEN_8914 == 8'h28 ? _GEN_7504 : _GEN_7088; // @[executor.scala 473:84]
  wire [7:0] _GEN_7509 = _GEN_8914 == 8'h28 ? _GEN_7505 : _GEN_7089; // @[executor.scala 473:84]
  wire [7:0] _GEN_7510 = mask_7[0] ? byte_1792 : _GEN_7090; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7511 = mask_7[1] ? byte_1793 : _GEN_7091; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7512 = mask_7[2] ? byte_1794 : _GEN_7092; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7513 = mask_7[3] ? byte_1795 : _GEN_7093; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7514 = _GEN_8914 == 8'h29 ? _GEN_7510 : _GEN_7090; // @[executor.scala 473:84]
  wire [7:0] _GEN_7515 = _GEN_8914 == 8'h29 ? _GEN_7511 : _GEN_7091; // @[executor.scala 473:84]
  wire [7:0] _GEN_7516 = _GEN_8914 == 8'h29 ? _GEN_7512 : _GEN_7092; // @[executor.scala 473:84]
  wire [7:0] _GEN_7517 = _GEN_8914 == 8'h29 ? _GEN_7513 : _GEN_7093; // @[executor.scala 473:84]
  wire [7:0] _GEN_7518 = mask_7[0] ? byte_1792 : _GEN_7094; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7519 = mask_7[1] ? byte_1793 : _GEN_7095; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7520 = mask_7[2] ? byte_1794 : _GEN_7096; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7521 = mask_7[3] ? byte_1795 : _GEN_7097; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7522 = _GEN_8914 == 8'h2a ? _GEN_7518 : _GEN_7094; // @[executor.scala 473:84]
  wire [7:0] _GEN_7523 = _GEN_8914 == 8'h2a ? _GEN_7519 : _GEN_7095; // @[executor.scala 473:84]
  wire [7:0] _GEN_7524 = _GEN_8914 == 8'h2a ? _GEN_7520 : _GEN_7096; // @[executor.scala 473:84]
  wire [7:0] _GEN_7525 = _GEN_8914 == 8'h2a ? _GEN_7521 : _GEN_7097; // @[executor.scala 473:84]
  wire [7:0] _GEN_7526 = mask_7[0] ? byte_1792 : _GEN_7098; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7527 = mask_7[1] ? byte_1793 : _GEN_7099; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7528 = mask_7[2] ? byte_1794 : _GEN_7100; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7529 = mask_7[3] ? byte_1795 : _GEN_7101; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7530 = _GEN_8914 == 8'h2b ? _GEN_7526 : _GEN_7098; // @[executor.scala 473:84]
  wire [7:0] _GEN_7531 = _GEN_8914 == 8'h2b ? _GEN_7527 : _GEN_7099; // @[executor.scala 473:84]
  wire [7:0] _GEN_7532 = _GEN_8914 == 8'h2b ? _GEN_7528 : _GEN_7100; // @[executor.scala 473:84]
  wire [7:0] _GEN_7533 = _GEN_8914 == 8'h2b ? _GEN_7529 : _GEN_7101; // @[executor.scala 473:84]
  wire [7:0] _GEN_7534 = mask_7[0] ? byte_1792 : _GEN_7102; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7535 = mask_7[1] ? byte_1793 : _GEN_7103; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7536 = mask_7[2] ? byte_1794 : _GEN_7104; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7537 = mask_7[3] ? byte_1795 : _GEN_7105; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7538 = _GEN_8914 == 8'h2c ? _GEN_7534 : _GEN_7102; // @[executor.scala 473:84]
  wire [7:0] _GEN_7539 = _GEN_8914 == 8'h2c ? _GEN_7535 : _GEN_7103; // @[executor.scala 473:84]
  wire [7:0] _GEN_7540 = _GEN_8914 == 8'h2c ? _GEN_7536 : _GEN_7104; // @[executor.scala 473:84]
  wire [7:0] _GEN_7541 = _GEN_8914 == 8'h2c ? _GEN_7537 : _GEN_7105; // @[executor.scala 473:84]
  wire [7:0] _GEN_7542 = mask_7[0] ? byte_1792 : _GEN_7106; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7543 = mask_7[1] ? byte_1793 : _GEN_7107; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7544 = mask_7[2] ? byte_1794 : _GEN_7108; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7545 = mask_7[3] ? byte_1795 : _GEN_7109; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7546 = _GEN_8914 == 8'h2d ? _GEN_7542 : _GEN_7106; // @[executor.scala 473:84]
  wire [7:0] _GEN_7547 = _GEN_8914 == 8'h2d ? _GEN_7543 : _GEN_7107; // @[executor.scala 473:84]
  wire [7:0] _GEN_7548 = _GEN_8914 == 8'h2d ? _GEN_7544 : _GEN_7108; // @[executor.scala 473:84]
  wire [7:0] _GEN_7549 = _GEN_8914 == 8'h2d ? _GEN_7545 : _GEN_7109; // @[executor.scala 473:84]
  wire [7:0] _GEN_7550 = mask_7[0] ? byte_1792 : _GEN_7110; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7551 = mask_7[1] ? byte_1793 : _GEN_7111; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7552 = mask_7[2] ? byte_1794 : _GEN_7112; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7553 = mask_7[3] ? byte_1795 : _GEN_7113; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7554 = _GEN_8914 == 8'h2e ? _GEN_7550 : _GEN_7110; // @[executor.scala 473:84]
  wire [7:0] _GEN_7555 = _GEN_8914 == 8'h2e ? _GEN_7551 : _GEN_7111; // @[executor.scala 473:84]
  wire [7:0] _GEN_7556 = _GEN_8914 == 8'h2e ? _GEN_7552 : _GEN_7112; // @[executor.scala 473:84]
  wire [7:0] _GEN_7557 = _GEN_8914 == 8'h2e ? _GEN_7553 : _GEN_7113; // @[executor.scala 473:84]
  wire [7:0] _GEN_7558 = mask_7[0] ? byte_1792 : _GEN_7114; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7559 = mask_7[1] ? byte_1793 : _GEN_7115; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7560 = mask_7[2] ? byte_1794 : _GEN_7116; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7561 = mask_7[3] ? byte_1795 : _GEN_7117; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7562 = _GEN_8914 == 8'h2f ? _GEN_7558 : _GEN_7114; // @[executor.scala 473:84]
  wire [7:0] _GEN_7563 = _GEN_8914 == 8'h2f ? _GEN_7559 : _GEN_7115; // @[executor.scala 473:84]
  wire [7:0] _GEN_7564 = _GEN_8914 == 8'h2f ? _GEN_7560 : _GEN_7116; // @[executor.scala 473:84]
  wire [7:0] _GEN_7565 = _GEN_8914 == 8'h2f ? _GEN_7561 : _GEN_7117; // @[executor.scala 473:84]
  wire [7:0] _GEN_7566 = mask_7[0] ? byte_1792 : _GEN_7118; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7567 = mask_7[1] ? byte_1793 : _GEN_7119; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7568 = mask_7[2] ? byte_1794 : _GEN_7120; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7569 = mask_7[3] ? byte_1795 : _GEN_7121; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7570 = _GEN_8914 == 8'h30 ? _GEN_7566 : _GEN_7118; // @[executor.scala 473:84]
  wire [7:0] _GEN_7571 = _GEN_8914 == 8'h30 ? _GEN_7567 : _GEN_7119; // @[executor.scala 473:84]
  wire [7:0] _GEN_7572 = _GEN_8914 == 8'h30 ? _GEN_7568 : _GEN_7120; // @[executor.scala 473:84]
  wire [7:0] _GEN_7573 = _GEN_8914 == 8'h30 ? _GEN_7569 : _GEN_7121; // @[executor.scala 473:84]
  wire [7:0] _GEN_7574 = mask_7[0] ? byte_1792 : _GEN_7122; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7575 = mask_7[1] ? byte_1793 : _GEN_7123; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7576 = mask_7[2] ? byte_1794 : _GEN_7124; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7577 = mask_7[3] ? byte_1795 : _GEN_7125; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7578 = _GEN_8914 == 8'h31 ? _GEN_7574 : _GEN_7122; // @[executor.scala 473:84]
  wire [7:0] _GEN_7579 = _GEN_8914 == 8'h31 ? _GEN_7575 : _GEN_7123; // @[executor.scala 473:84]
  wire [7:0] _GEN_7580 = _GEN_8914 == 8'h31 ? _GEN_7576 : _GEN_7124; // @[executor.scala 473:84]
  wire [7:0] _GEN_7581 = _GEN_8914 == 8'h31 ? _GEN_7577 : _GEN_7125; // @[executor.scala 473:84]
  wire [7:0] _GEN_7582 = mask_7[0] ? byte_1792 : _GEN_7126; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7583 = mask_7[1] ? byte_1793 : _GEN_7127; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7584 = mask_7[2] ? byte_1794 : _GEN_7128; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7585 = mask_7[3] ? byte_1795 : _GEN_7129; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7586 = _GEN_8914 == 8'h32 ? _GEN_7582 : _GEN_7126; // @[executor.scala 473:84]
  wire [7:0] _GEN_7587 = _GEN_8914 == 8'h32 ? _GEN_7583 : _GEN_7127; // @[executor.scala 473:84]
  wire [7:0] _GEN_7588 = _GEN_8914 == 8'h32 ? _GEN_7584 : _GEN_7128; // @[executor.scala 473:84]
  wire [7:0] _GEN_7589 = _GEN_8914 == 8'h32 ? _GEN_7585 : _GEN_7129; // @[executor.scala 473:84]
  wire [7:0] _GEN_7590 = mask_7[0] ? byte_1792 : _GEN_7130; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7591 = mask_7[1] ? byte_1793 : _GEN_7131; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7592 = mask_7[2] ? byte_1794 : _GEN_7132; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7593 = mask_7[3] ? byte_1795 : _GEN_7133; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7594 = _GEN_8914 == 8'h33 ? _GEN_7590 : _GEN_7130; // @[executor.scala 473:84]
  wire [7:0] _GEN_7595 = _GEN_8914 == 8'h33 ? _GEN_7591 : _GEN_7131; // @[executor.scala 473:84]
  wire [7:0] _GEN_7596 = _GEN_8914 == 8'h33 ? _GEN_7592 : _GEN_7132; // @[executor.scala 473:84]
  wire [7:0] _GEN_7597 = _GEN_8914 == 8'h33 ? _GEN_7593 : _GEN_7133; // @[executor.scala 473:84]
  wire [7:0] _GEN_7598 = mask_7[0] ? byte_1792 : _GEN_7134; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7599 = mask_7[1] ? byte_1793 : _GEN_7135; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7600 = mask_7[2] ? byte_1794 : _GEN_7136; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7601 = mask_7[3] ? byte_1795 : _GEN_7137; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7602 = _GEN_8914 == 8'h34 ? _GEN_7598 : _GEN_7134; // @[executor.scala 473:84]
  wire [7:0] _GEN_7603 = _GEN_8914 == 8'h34 ? _GEN_7599 : _GEN_7135; // @[executor.scala 473:84]
  wire [7:0] _GEN_7604 = _GEN_8914 == 8'h34 ? _GEN_7600 : _GEN_7136; // @[executor.scala 473:84]
  wire [7:0] _GEN_7605 = _GEN_8914 == 8'h34 ? _GEN_7601 : _GEN_7137; // @[executor.scala 473:84]
  wire [7:0] _GEN_7606 = mask_7[0] ? byte_1792 : _GEN_7138; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7607 = mask_7[1] ? byte_1793 : _GEN_7139; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7608 = mask_7[2] ? byte_1794 : _GEN_7140; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7609 = mask_7[3] ? byte_1795 : _GEN_7141; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7610 = _GEN_8914 == 8'h35 ? _GEN_7606 : _GEN_7138; // @[executor.scala 473:84]
  wire [7:0] _GEN_7611 = _GEN_8914 == 8'h35 ? _GEN_7607 : _GEN_7139; // @[executor.scala 473:84]
  wire [7:0] _GEN_7612 = _GEN_8914 == 8'h35 ? _GEN_7608 : _GEN_7140; // @[executor.scala 473:84]
  wire [7:0] _GEN_7613 = _GEN_8914 == 8'h35 ? _GEN_7609 : _GEN_7141; // @[executor.scala 473:84]
  wire [7:0] _GEN_7614 = mask_7[0] ? byte_1792 : _GEN_7142; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7615 = mask_7[1] ? byte_1793 : _GEN_7143; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7616 = mask_7[2] ? byte_1794 : _GEN_7144; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7617 = mask_7[3] ? byte_1795 : _GEN_7145; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7618 = _GEN_8914 == 8'h36 ? _GEN_7614 : _GEN_7142; // @[executor.scala 473:84]
  wire [7:0] _GEN_7619 = _GEN_8914 == 8'h36 ? _GEN_7615 : _GEN_7143; // @[executor.scala 473:84]
  wire [7:0] _GEN_7620 = _GEN_8914 == 8'h36 ? _GEN_7616 : _GEN_7144; // @[executor.scala 473:84]
  wire [7:0] _GEN_7621 = _GEN_8914 == 8'h36 ? _GEN_7617 : _GEN_7145; // @[executor.scala 473:84]
  wire [7:0] _GEN_7622 = mask_7[0] ? byte_1792 : _GEN_7146; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7623 = mask_7[1] ? byte_1793 : _GEN_7147; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7624 = mask_7[2] ? byte_1794 : _GEN_7148; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7625 = mask_7[3] ? byte_1795 : _GEN_7149; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7626 = _GEN_8914 == 8'h37 ? _GEN_7622 : _GEN_7146; // @[executor.scala 473:84]
  wire [7:0] _GEN_7627 = _GEN_8914 == 8'h37 ? _GEN_7623 : _GEN_7147; // @[executor.scala 473:84]
  wire [7:0] _GEN_7628 = _GEN_8914 == 8'h37 ? _GEN_7624 : _GEN_7148; // @[executor.scala 473:84]
  wire [7:0] _GEN_7629 = _GEN_8914 == 8'h37 ? _GEN_7625 : _GEN_7149; // @[executor.scala 473:84]
  wire [7:0] _GEN_7630 = mask_7[0] ? byte_1792 : _GEN_7150; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7631 = mask_7[1] ? byte_1793 : _GEN_7151; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7632 = mask_7[2] ? byte_1794 : _GEN_7152; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7633 = mask_7[3] ? byte_1795 : _GEN_7153; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7634 = _GEN_8914 == 8'h38 ? _GEN_7630 : _GEN_7150; // @[executor.scala 473:84]
  wire [7:0] _GEN_7635 = _GEN_8914 == 8'h38 ? _GEN_7631 : _GEN_7151; // @[executor.scala 473:84]
  wire [7:0] _GEN_7636 = _GEN_8914 == 8'h38 ? _GEN_7632 : _GEN_7152; // @[executor.scala 473:84]
  wire [7:0] _GEN_7637 = _GEN_8914 == 8'h38 ? _GEN_7633 : _GEN_7153; // @[executor.scala 473:84]
  wire [7:0] _GEN_7638 = mask_7[0] ? byte_1792 : _GEN_7154; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7639 = mask_7[1] ? byte_1793 : _GEN_7155; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7640 = mask_7[2] ? byte_1794 : _GEN_7156; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7641 = mask_7[3] ? byte_1795 : _GEN_7157; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7642 = _GEN_8914 == 8'h39 ? _GEN_7638 : _GEN_7154; // @[executor.scala 473:84]
  wire [7:0] _GEN_7643 = _GEN_8914 == 8'h39 ? _GEN_7639 : _GEN_7155; // @[executor.scala 473:84]
  wire [7:0] _GEN_7644 = _GEN_8914 == 8'h39 ? _GEN_7640 : _GEN_7156; // @[executor.scala 473:84]
  wire [7:0] _GEN_7645 = _GEN_8914 == 8'h39 ? _GEN_7641 : _GEN_7157; // @[executor.scala 473:84]
  wire [7:0] _GEN_7646 = mask_7[0] ? byte_1792 : _GEN_7158; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7647 = mask_7[1] ? byte_1793 : _GEN_7159; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7648 = mask_7[2] ? byte_1794 : _GEN_7160; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7649 = mask_7[3] ? byte_1795 : _GEN_7161; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7650 = _GEN_8914 == 8'h3a ? _GEN_7646 : _GEN_7158; // @[executor.scala 473:84]
  wire [7:0] _GEN_7651 = _GEN_8914 == 8'h3a ? _GEN_7647 : _GEN_7159; // @[executor.scala 473:84]
  wire [7:0] _GEN_7652 = _GEN_8914 == 8'h3a ? _GEN_7648 : _GEN_7160; // @[executor.scala 473:84]
  wire [7:0] _GEN_7653 = _GEN_8914 == 8'h3a ? _GEN_7649 : _GEN_7161; // @[executor.scala 473:84]
  wire [7:0] _GEN_7654 = mask_7[0] ? byte_1792 : _GEN_7162; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7655 = mask_7[1] ? byte_1793 : _GEN_7163; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7656 = mask_7[2] ? byte_1794 : _GEN_7164; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7657 = mask_7[3] ? byte_1795 : _GEN_7165; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7658 = _GEN_8914 == 8'h3b ? _GEN_7654 : _GEN_7162; // @[executor.scala 473:84]
  wire [7:0] _GEN_7659 = _GEN_8914 == 8'h3b ? _GEN_7655 : _GEN_7163; // @[executor.scala 473:84]
  wire [7:0] _GEN_7660 = _GEN_8914 == 8'h3b ? _GEN_7656 : _GEN_7164; // @[executor.scala 473:84]
  wire [7:0] _GEN_7661 = _GEN_8914 == 8'h3b ? _GEN_7657 : _GEN_7165; // @[executor.scala 473:84]
  wire [7:0] _GEN_7662 = mask_7[0] ? byte_1792 : _GEN_7166; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7663 = mask_7[1] ? byte_1793 : _GEN_7167; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7664 = mask_7[2] ? byte_1794 : _GEN_7168; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7665 = mask_7[3] ? byte_1795 : _GEN_7169; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7666 = _GEN_8914 == 8'h3c ? _GEN_7662 : _GEN_7166; // @[executor.scala 473:84]
  wire [7:0] _GEN_7667 = _GEN_8914 == 8'h3c ? _GEN_7663 : _GEN_7167; // @[executor.scala 473:84]
  wire [7:0] _GEN_7668 = _GEN_8914 == 8'h3c ? _GEN_7664 : _GEN_7168; // @[executor.scala 473:84]
  wire [7:0] _GEN_7669 = _GEN_8914 == 8'h3c ? _GEN_7665 : _GEN_7169; // @[executor.scala 473:84]
  wire [7:0] _GEN_7670 = mask_7[0] ? byte_1792 : _GEN_7170; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7671 = mask_7[1] ? byte_1793 : _GEN_7171; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7672 = mask_7[2] ? byte_1794 : _GEN_7172; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7673 = mask_7[3] ? byte_1795 : _GEN_7173; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7674 = _GEN_8914 == 8'h3d ? _GEN_7670 : _GEN_7170; // @[executor.scala 473:84]
  wire [7:0] _GEN_7675 = _GEN_8914 == 8'h3d ? _GEN_7671 : _GEN_7171; // @[executor.scala 473:84]
  wire [7:0] _GEN_7676 = _GEN_8914 == 8'h3d ? _GEN_7672 : _GEN_7172; // @[executor.scala 473:84]
  wire [7:0] _GEN_7677 = _GEN_8914 == 8'h3d ? _GEN_7673 : _GEN_7173; // @[executor.scala 473:84]
  wire [7:0] _GEN_7678 = mask_7[0] ? byte_1792 : _GEN_7174; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7679 = mask_7[1] ? byte_1793 : _GEN_7175; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7680 = mask_7[2] ? byte_1794 : _GEN_7176; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7681 = mask_7[3] ? byte_1795 : _GEN_7177; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7682 = _GEN_8914 == 8'h3e ? _GEN_7678 : _GEN_7174; // @[executor.scala 473:84]
  wire [7:0] _GEN_7683 = _GEN_8914 == 8'h3e ? _GEN_7679 : _GEN_7175; // @[executor.scala 473:84]
  wire [7:0] _GEN_7684 = _GEN_8914 == 8'h3e ? _GEN_7680 : _GEN_7176; // @[executor.scala 473:84]
  wire [7:0] _GEN_7685 = _GEN_8914 == 8'h3e ? _GEN_7681 : _GEN_7177; // @[executor.scala 473:84]
  wire [7:0] _GEN_7686 = mask_7[0] ? byte_1792 : _GEN_7178; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7687 = mask_7[1] ? byte_1793 : _GEN_7179; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7688 = mask_7[2] ? byte_1794 : _GEN_7180; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7689 = mask_7[3] ? byte_1795 : _GEN_7181; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7690 = _GEN_8914 == 8'h3f ? _GEN_7686 : _GEN_7178; // @[executor.scala 473:84]
  wire [7:0] _GEN_7691 = _GEN_8914 == 8'h3f ? _GEN_7687 : _GEN_7179; // @[executor.scala 473:84]
  wire [7:0] _GEN_7692 = _GEN_8914 == 8'h3f ? _GEN_7688 : _GEN_7180; // @[executor.scala 473:84]
  wire [7:0] _GEN_7693 = _GEN_8914 == 8'h3f ? _GEN_7689 : _GEN_7181; // @[executor.scala 473:84]
  wire [7:0] _GEN_7694 = opcode_7 != 4'h0 ? _GEN_7186 : _GEN_6926; // @[executor.scala 470:55]
  wire [7:0] _GEN_7695 = opcode_7 != 4'h0 ? _GEN_7187 : _GEN_6927; // @[executor.scala 470:55]
  wire [7:0] _GEN_7696 = opcode_7 != 4'h0 ? _GEN_7188 : _GEN_6928; // @[executor.scala 470:55]
  wire [7:0] _GEN_7697 = opcode_7 != 4'h0 ? _GEN_7189 : _GEN_6929; // @[executor.scala 470:55]
  wire [7:0] _GEN_7698 = opcode_7 != 4'h0 ? _GEN_7194 : _GEN_6930; // @[executor.scala 470:55]
  wire [7:0] _GEN_7699 = opcode_7 != 4'h0 ? _GEN_7195 : _GEN_6931; // @[executor.scala 470:55]
  wire [7:0] _GEN_7700 = opcode_7 != 4'h0 ? _GEN_7196 : _GEN_6932; // @[executor.scala 470:55]
  wire [7:0] _GEN_7701 = opcode_7 != 4'h0 ? _GEN_7197 : _GEN_6933; // @[executor.scala 470:55]
  wire [7:0] _GEN_7702 = opcode_7 != 4'h0 ? _GEN_7202 : _GEN_6934; // @[executor.scala 470:55]
  wire [7:0] _GEN_7703 = opcode_7 != 4'h0 ? _GEN_7203 : _GEN_6935; // @[executor.scala 470:55]
  wire [7:0] _GEN_7704 = opcode_7 != 4'h0 ? _GEN_7204 : _GEN_6936; // @[executor.scala 470:55]
  wire [7:0] _GEN_7705 = opcode_7 != 4'h0 ? _GEN_7205 : _GEN_6937; // @[executor.scala 470:55]
  wire [7:0] _GEN_7706 = opcode_7 != 4'h0 ? _GEN_7210 : _GEN_6938; // @[executor.scala 470:55]
  wire [7:0] _GEN_7707 = opcode_7 != 4'h0 ? _GEN_7211 : _GEN_6939; // @[executor.scala 470:55]
  wire [7:0] _GEN_7708 = opcode_7 != 4'h0 ? _GEN_7212 : _GEN_6940; // @[executor.scala 470:55]
  wire [7:0] _GEN_7709 = opcode_7 != 4'h0 ? _GEN_7213 : _GEN_6941; // @[executor.scala 470:55]
  wire [7:0] _GEN_7710 = opcode_7 != 4'h0 ? _GEN_7218 : _GEN_6942; // @[executor.scala 470:55]
  wire [7:0] _GEN_7711 = opcode_7 != 4'h0 ? _GEN_7219 : _GEN_6943; // @[executor.scala 470:55]
  wire [7:0] _GEN_7712 = opcode_7 != 4'h0 ? _GEN_7220 : _GEN_6944; // @[executor.scala 470:55]
  wire [7:0] _GEN_7713 = opcode_7 != 4'h0 ? _GEN_7221 : _GEN_6945; // @[executor.scala 470:55]
  wire [7:0] _GEN_7714 = opcode_7 != 4'h0 ? _GEN_7226 : _GEN_6946; // @[executor.scala 470:55]
  wire [7:0] _GEN_7715 = opcode_7 != 4'h0 ? _GEN_7227 : _GEN_6947; // @[executor.scala 470:55]
  wire [7:0] _GEN_7716 = opcode_7 != 4'h0 ? _GEN_7228 : _GEN_6948; // @[executor.scala 470:55]
  wire [7:0] _GEN_7717 = opcode_7 != 4'h0 ? _GEN_7229 : _GEN_6949; // @[executor.scala 470:55]
  wire [7:0] _GEN_7718 = opcode_7 != 4'h0 ? _GEN_7234 : _GEN_6950; // @[executor.scala 470:55]
  wire [7:0] _GEN_7719 = opcode_7 != 4'h0 ? _GEN_7235 : _GEN_6951; // @[executor.scala 470:55]
  wire [7:0] _GEN_7720 = opcode_7 != 4'h0 ? _GEN_7236 : _GEN_6952; // @[executor.scala 470:55]
  wire [7:0] _GEN_7721 = opcode_7 != 4'h0 ? _GEN_7237 : _GEN_6953; // @[executor.scala 470:55]
  wire [7:0] _GEN_7722 = opcode_7 != 4'h0 ? _GEN_7242 : _GEN_6954; // @[executor.scala 470:55]
  wire [7:0] _GEN_7723 = opcode_7 != 4'h0 ? _GEN_7243 : _GEN_6955; // @[executor.scala 470:55]
  wire [7:0] _GEN_7724 = opcode_7 != 4'h0 ? _GEN_7244 : _GEN_6956; // @[executor.scala 470:55]
  wire [7:0] _GEN_7725 = opcode_7 != 4'h0 ? _GEN_7245 : _GEN_6957; // @[executor.scala 470:55]
  wire [7:0] _GEN_7726 = opcode_7 != 4'h0 ? _GEN_7250 : _GEN_6958; // @[executor.scala 470:55]
  wire [7:0] _GEN_7727 = opcode_7 != 4'h0 ? _GEN_7251 : _GEN_6959; // @[executor.scala 470:55]
  wire [7:0] _GEN_7728 = opcode_7 != 4'h0 ? _GEN_7252 : _GEN_6960; // @[executor.scala 470:55]
  wire [7:0] _GEN_7729 = opcode_7 != 4'h0 ? _GEN_7253 : _GEN_6961; // @[executor.scala 470:55]
  wire [7:0] _GEN_7730 = opcode_7 != 4'h0 ? _GEN_7258 : _GEN_6962; // @[executor.scala 470:55]
  wire [7:0] _GEN_7731 = opcode_7 != 4'h0 ? _GEN_7259 : _GEN_6963; // @[executor.scala 470:55]
  wire [7:0] _GEN_7732 = opcode_7 != 4'h0 ? _GEN_7260 : _GEN_6964; // @[executor.scala 470:55]
  wire [7:0] _GEN_7733 = opcode_7 != 4'h0 ? _GEN_7261 : _GEN_6965; // @[executor.scala 470:55]
  wire [7:0] _GEN_7734 = opcode_7 != 4'h0 ? _GEN_7266 : _GEN_6966; // @[executor.scala 470:55]
  wire [7:0] _GEN_7735 = opcode_7 != 4'h0 ? _GEN_7267 : _GEN_6967; // @[executor.scala 470:55]
  wire [7:0] _GEN_7736 = opcode_7 != 4'h0 ? _GEN_7268 : _GEN_6968; // @[executor.scala 470:55]
  wire [7:0] _GEN_7737 = opcode_7 != 4'h0 ? _GEN_7269 : _GEN_6969; // @[executor.scala 470:55]
  wire [7:0] _GEN_7738 = opcode_7 != 4'h0 ? _GEN_7274 : _GEN_6970; // @[executor.scala 470:55]
  wire [7:0] _GEN_7739 = opcode_7 != 4'h0 ? _GEN_7275 : _GEN_6971; // @[executor.scala 470:55]
  wire [7:0] _GEN_7740 = opcode_7 != 4'h0 ? _GEN_7276 : _GEN_6972; // @[executor.scala 470:55]
  wire [7:0] _GEN_7741 = opcode_7 != 4'h0 ? _GEN_7277 : _GEN_6973; // @[executor.scala 470:55]
  wire [7:0] _GEN_7742 = opcode_7 != 4'h0 ? _GEN_7282 : _GEN_6974; // @[executor.scala 470:55]
  wire [7:0] _GEN_7743 = opcode_7 != 4'h0 ? _GEN_7283 : _GEN_6975; // @[executor.scala 470:55]
  wire [7:0] _GEN_7744 = opcode_7 != 4'h0 ? _GEN_7284 : _GEN_6976; // @[executor.scala 470:55]
  wire [7:0] _GEN_7745 = opcode_7 != 4'h0 ? _GEN_7285 : _GEN_6977; // @[executor.scala 470:55]
  wire [7:0] _GEN_7746 = opcode_7 != 4'h0 ? _GEN_7290 : _GEN_6978; // @[executor.scala 470:55]
  wire [7:0] _GEN_7747 = opcode_7 != 4'h0 ? _GEN_7291 : _GEN_6979; // @[executor.scala 470:55]
  wire [7:0] _GEN_7748 = opcode_7 != 4'h0 ? _GEN_7292 : _GEN_6980; // @[executor.scala 470:55]
  wire [7:0] _GEN_7749 = opcode_7 != 4'h0 ? _GEN_7293 : _GEN_6981; // @[executor.scala 470:55]
  wire [7:0] _GEN_7750 = opcode_7 != 4'h0 ? _GEN_7298 : _GEN_6982; // @[executor.scala 470:55]
  wire [7:0] _GEN_7751 = opcode_7 != 4'h0 ? _GEN_7299 : _GEN_6983; // @[executor.scala 470:55]
  wire [7:0] _GEN_7752 = opcode_7 != 4'h0 ? _GEN_7300 : _GEN_6984; // @[executor.scala 470:55]
  wire [7:0] _GEN_7753 = opcode_7 != 4'h0 ? _GEN_7301 : _GEN_6985; // @[executor.scala 470:55]
  wire [7:0] _GEN_7754 = opcode_7 != 4'h0 ? _GEN_7306 : _GEN_6986; // @[executor.scala 470:55]
  wire [7:0] _GEN_7755 = opcode_7 != 4'h0 ? _GEN_7307 : _GEN_6987; // @[executor.scala 470:55]
  wire [7:0] _GEN_7756 = opcode_7 != 4'h0 ? _GEN_7308 : _GEN_6988; // @[executor.scala 470:55]
  wire [7:0] _GEN_7757 = opcode_7 != 4'h0 ? _GEN_7309 : _GEN_6989; // @[executor.scala 470:55]
  wire [7:0] _GEN_7758 = opcode_7 != 4'h0 ? _GEN_7314 : _GEN_6990; // @[executor.scala 470:55]
  wire [7:0] _GEN_7759 = opcode_7 != 4'h0 ? _GEN_7315 : _GEN_6991; // @[executor.scala 470:55]
  wire [7:0] _GEN_7760 = opcode_7 != 4'h0 ? _GEN_7316 : _GEN_6992; // @[executor.scala 470:55]
  wire [7:0] _GEN_7761 = opcode_7 != 4'h0 ? _GEN_7317 : _GEN_6993; // @[executor.scala 470:55]
  wire [7:0] _GEN_7762 = opcode_7 != 4'h0 ? _GEN_7322 : _GEN_6994; // @[executor.scala 470:55]
  wire [7:0] _GEN_7763 = opcode_7 != 4'h0 ? _GEN_7323 : _GEN_6995; // @[executor.scala 470:55]
  wire [7:0] _GEN_7764 = opcode_7 != 4'h0 ? _GEN_7324 : _GEN_6996; // @[executor.scala 470:55]
  wire [7:0] _GEN_7765 = opcode_7 != 4'h0 ? _GEN_7325 : _GEN_6997; // @[executor.scala 470:55]
  wire [7:0] _GEN_7766 = opcode_7 != 4'h0 ? _GEN_7330 : _GEN_6998; // @[executor.scala 470:55]
  wire [7:0] _GEN_7767 = opcode_7 != 4'h0 ? _GEN_7331 : _GEN_6999; // @[executor.scala 470:55]
  wire [7:0] _GEN_7768 = opcode_7 != 4'h0 ? _GEN_7332 : _GEN_7000; // @[executor.scala 470:55]
  wire [7:0] _GEN_7769 = opcode_7 != 4'h0 ? _GEN_7333 : _GEN_7001; // @[executor.scala 470:55]
  wire [7:0] _GEN_7770 = opcode_7 != 4'h0 ? _GEN_7338 : _GEN_7002; // @[executor.scala 470:55]
  wire [7:0] _GEN_7771 = opcode_7 != 4'h0 ? _GEN_7339 : _GEN_7003; // @[executor.scala 470:55]
  wire [7:0] _GEN_7772 = opcode_7 != 4'h0 ? _GEN_7340 : _GEN_7004; // @[executor.scala 470:55]
  wire [7:0] _GEN_7773 = opcode_7 != 4'h0 ? _GEN_7341 : _GEN_7005; // @[executor.scala 470:55]
  wire [7:0] _GEN_7774 = opcode_7 != 4'h0 ? _GEN_7346 : _GEN_7006; // @[executor.scala 470:55]
  wire [7:0] _GEN_7775 = opcode_7 != 4'h0 ? _GEN_7347 : _GEN_7007; // @[executor.scala 470:55]
  wire [7:0] _GEN_7776 = opcode_7 != 4'h0 ? _GEN_7348 : _GEN_7008; // @[executor.scala 470:55]
  wire [7:0] _GEN_7777 = opcode_7 != 4'h0 ? _GEN_7349 : _GEN_7009; // @[executor.scala 470:55]
  wire [7:0] _GEN_7778 = opcode_7 != 4'h0 ? _GEN_7354 : _GEN_7010; // @[executor.scala 470:55]
  wire [7:0] _GEN_7779 = opcode_7 != 4'h0 ? _GEN_7355 : _GEN_7011; // @[executor.scala 470:55]
  wire [7:0] _GEN_7780 = opcode_7 != 4'h0 ? _GEN_7356 : _GEN_7012; // @[executor.scala 470:55]
  wire [7:0] _GEN_7781 = opcode_7 != 4'h0 ? _GEN_7357 : _GEN_7013; // @[executor.scala 470:55]
  wire [7:0] _GEN_7782 = opcode_7 != 4'h0 ? _GEN_7362 : _GEN_7014; // @[executor.scala 470:55]
  wire [7:0] _GEN_7783 = opcode_7 != 4'h0 ? _GEN_7363 : _GEN_7015; // @[executor.scala 470:55]
  wire [7:0] _GEN_7784 = opcode_7 != 4'h0 ? _GEN_7364 : _GEN_7016; // @[executor.scala 470:55]
  wire [7:0] _GEN_7785 = opcode_7 != 4'h0 ? _GEN_7365 : _GEN_7017; // @[executor.scala 470:55]
  wire [7:0] _GEN_7786 = opcode_7 != 4'h0 ? _GEN_7370 : _GEN_7018; // @[executor.scala 470:55]
  wire [7:0] _GEN_7787 = opcode_7 != 4'h0 ? _GEN_7371 : _GEN_7019; // @[executor.scala 470:55]
  wire [7:0] _GEN_7788 = opcode_7 != 4'h0 ? _GEN_7372 : _GEN_7020; // @[executor.scala 470:55]
  wire [7:0] _GEN_7789 = opcode_7 != 4'h0 ? _GEN_7373 : _GEN_7021; // @[executor.scala 470:55]
  wire [7:0] _GEN_7790 = opcode_7 != 4'h0 ? _GEN_7378 : _GEN_7022; // @[executor.scala 470:55]
  wire [7:0] _GEN_7791 = opcode_7 != 4'h0 ? _GEN_7379 : _GEN_7023; // @[executor.scala 470:55]
  wire [7:0] _GEN_7792 = opcode_7 != 4'h0 ? _GEN_7380 : _GEN_7024; // @[executor.scala 470:55]
  wire [7:0] _GEN_7793 = opcode_7 != 4'h0 ? _GEN_7381 : _GEN_7025; // @[executor.scala 470:55]
  wire [7:0] _GEN_7794 = opcode_7 != 4'h0 ? _GEN_7386 : _GEN_7026; // @[executor.scala 470:55]
  wire [7:0] _GEN_7795 = opcode_7 != 4'h0 ? _GEN_7387 : _GEN_7027; // @[executor.scala 470:55]
  wire [7:0] _GEN_7796 = opcode_7 != 4'h0 ? _GEN_7388 : _GEN_7028; // @[executor.scala 470:55]
  wire [7:0] _GEN_7797 = opcode_7 != 4'h0 ? _GEN_7389 : _GEN_7029; // @[executor.scala 470:55]
  wire [7:0] _GEN_7798 = opcode_7 != 4'h0 ? _GEN_7394 : _GEN_7030; // @[executor.scala 470:55]
  wire [7:0] _GEN_7799 = opcode_7 != 4'h0 ? _GEN_7395 : _GEN_7031; // @[executor.scala 470:55]
  wire [7:0] _GEN_7800 = opcode_7 != 4'h0 ? _GEN_7396 : _GEN_7032; // @[executor.scala 470:55]
  wire [7:0] _GEN_7801 = opcode_7 != 4'h0 ? _GEN_7397 : _GEN_7033; // @[executor.scala 470:55]
  wire [7:0] _GEN_7802 = opcode_7 != 4'h0 ? _GEN_7402 : _GEN_7034; // @[executor.scala 470:55]
  wire [7:0] _GEN_7803 = opcode_7 != 4'h0 ? _GEN_7403 : _GEN_7035; // @[executor.scala 470:55]
  wire [7:0] _GEN_7804 = opcode_7 != 4'h0 ? _GEN_7404 : _GEN_7036; // @[executor.scala 470:55]
  wire [7:0] _GEN_7805 = opcode_7 != 4'h0 ? _GEN_7405 : _GEN_7037; // @[executor.scala 470:55]
  wire [7:0] _GEN_7806 = opcode_7 != 4'h0 ? _GEN_7410 : _GEN_7038; // @[executor.scala 470:55]
  wire [7:0] _GEN_7807 = opcode_7 != 4'h0 ? _GEN_7411 : _GEN_7039; // @[executor.scala 470:55]
  wire [7:0] _GEN_7808 = opcode_7 != 4'h0 ? _GEN_7412 : _GEN_7040; // @[executor.scala 470:55]
  wire [7:0] _GEN_7809 = opcode_7 != 4'h0 ? _GEN_7413 : _GEN_7041; // @[executor.scala 470:55]
  wire [7:0] _GEN_7810 = opcode_7 != 4'h0 ? _GEN_7418 : _GEN_7042; // @[executor.scala 470:55]
  wire [7:0] _GEN_7811 = opcode_7 != 4'h0 ? _GEN_7419 : _GEN_7043; // @[executor.scala 470:55]
  wire [7:0] _GEN_7812 = opcode_7 != 4'h0 ? _GEN_7420 : _GEN_7044; // @[executor.scala 470:55]
  wire [7:0] _GEN_7813 = opcode_7 != 4'h0 ? _GEN_7421 : _GEN_7045; // @[executor.scala 470:55]
  wire [7:0] _GEN_7814 = opcode_7 != 4'h0 ? _GEN_7426 : _GEN_7046; // @[executor.scala 470:55]
  wire [7:0] _GEN_7815 = opcode_7 != 4'h0 ? _GEN_7427 : _GEN_7047; // @[executor.scala 470:55]
  wire [7:0] _GEN_7816 = opcode_7 != 4'h0 ? _GEN_7428 : _GEN_7048; // @[executor.scala 470:55]
  wire [7:0] _GEN_7817 = opcode_7 != 4'h0 ? _GEN_7429 : _GEN_7049; // @[executor.scala 470:55]
  wire [7:0] _GEN_7818 = opcode_7 != 4'h0 ? _GEN_7434 : _GEN_7050; // @[executor.scala 470:55]
  wire [7:0] _GEN_7819 = opcode_7 != 4'h0 ? _GEN_7435 : _GEN_7051; // @[executor.scala 470:55]
  wire [7:0] _GEN_7820 = opcode_7 != 4'h0 ? _GEN_7436 : _GEN_7052; // @[executor.scala 470:55]
  wire [7:0] _GEN_7821 = opcode_7 != 4'h0 ? _GEN_7437 : _GEN_7053; // @[executor.scala 470:55]
  wire [7:0] _GEN_7822 = opcode_7 != 4'h0 ? _GEN_7442 : _GEN_7054; // @[executor.scala 470:55]
  wire [7:0] _GEN_7823 = opcode_7 != 4'h0 ? _GEN_7443 : _GEN_7055; // @[executor.scala 470:55]
  wire [7:0] _GEN_7824 = opcode_7 != 4'h0 ? _GEN_7444 : _GEN_7056; // @[executor.scala 470:55]
  wire [7:0] _GEN_7825 = opcode_7 != 4'h0 ? _GEN_7445 : _GEN_7057; // @[executor.scala 470:55]
  wire [7:0] _GEN_7826 = opcode_7 != 4'h0 ? _GEN_7450 : _GEN_7058; // @[executor.scala 470:55]
  wire [7:0] _GEN_7827 = opcode_7 != 4'h0 ? _GEN_7451 : _GEN_7059; // @[executor.scala 470:55]
  wire [7:0] _GEN_7828 = opcode_7 != 4'h0 ? _GEN_7452 : _GEN_7060; // @[executor.scala 470:55]
  wire [7:0] _GEN_7829 = opcode_7 != 4'h0 ? _GEN_7453 : _GEN_7061; // @[executor.scala 470:55]
  wire [7:0] _GEN_7830 = opcode_7 != 4'h0 ? _GEN_7458 : _GEN_7062; // @[executor.scala 470:55]
  wire [7:0] _GEN_7831 = opcode_7 != 4'h0 ? _GEN_7459 : _GEN_7063; // @[executor.scala 470:55]
  wire [7:0] _GEN_7832 = opcode_7 != 4'h0 ? _GEN_7460 : _GEN_7064; // @[executor.scala 470:55]
  wire [7:0] _GEN_7833 = opcode_7 != 4'h0 ? _GEN_7461 : _GEN_7065; // @[executor.scala 470:55]
  wire [7:0] _GEN_7834 = opcode_7 != 4'h0 ? _GEN_7466 : _GEN_7066; // @[executor.scala 470:55]
  wire [7:0] _GEN_7835 = opcode_7 != 4'h0 ? _GEN_7467 : _GEN_7067; // @[executor.scala 470:55]
  wire [7:0] _GEN_7836 = opcode_7 != 4'h0 ? _GEN_7468 : _GEN_7068; // @[executor.scala 470:55]
  wire [7:0] _GEN_7837 = opcode_7 != 4'h0 ? _GEN_7469 : _GEN_7069; // @[executor.scala 470:55]
  wire [7:0] _GEN_7838 = opcode_7 != 4'h0 ? _GEN_7474 : _GEN_7070; // @[executor.scala 470:55]
  wire [7:0] _GEN_7839 = opcode_7 != 4'h0 ? _GEN_7475 : _GEN_7071; // @[executor.scala 470:55]
  wire [7:0] _GEN_7840 = opcode_7 != 4'h0 ? _GEN_7476 : _GEN_7072; // @[executor.scala 470:55]
  wire [7:0] _GEN_7841 = opcode_7 != 4'h0 ? _GEN_7477 : _GEN_7073; // @[executor.scala 470:55]
  wire [7:0] _GEN_7842 = opcode_7 != 4'h0 ? _GEN_7482 : _GEN_7074; // @[executor.scala 470:55]
  wire [7:0] _GEN_7843 = opcode_7 != 4'h0 ? _GEN_7483 : _GEN_7075; // @[executor.scala 470:55]
  wire [7:0] _GEN_7844 = opcode_7 != 4'h0 ? _GEN_7484 : _GEN_7076; // @[executor.scala 470:55]
  wire [7:0] _GEN_7845 = opcode_7 != 4'h0 ? _GEN_7485 : _GEN_7077; // @[executor.scala 470:55]
  wire [7:0] _GEN_7846 = opcode_7 != 4'h0 ? _GEN_7490 : _GEN_7078; // @[executor.scala 470:55]
  wire [7:0] _GEN_7847 = opcode_7 != 4'h0 ? _GEN_7491 : _GEN_7079; // @[executor.scala 470:55]
  wire [7:0] _GEN_7848 = opcode_7 != 4'h0 ? _GEN_7492 : _GEN_7080; // @[executor.scala 470:55]
  wire [7:0] _GEN_7849 = opcode_7 != 4'h0 ? _GEN_7493 : _GEN_7081; // @[executor.scala 470:55]
  wire [7:0] _GEN_7850 = opcode_7 != 4'h0 ? _GEN_7498 : _GEN_7082; // @[executor.scala 470:55]
  wire [7:0] _GEN_7851 = opcode_7 != 4'h0 ? _GEN_7499 : _GEN_7083; // @[executor.scala 470:55]
  wire [7:0] _GEN_7852 = opcode_7 != 4'h0 ? _GEN_7500 : _GEN_7084; // @[executor.scala 470:55]
  wire [7:0] _GEN_7853 = opcode_7 != 4'h0 ? _GEN_7501 : _GEN_7085; // @[executor.scala 470:55]
  wire [7:0] _GEN_7854 = opcode_7 != 4'h0 ? _GEN_7506 : _GEN_7086; // @[executor.scala 470:55]
  wire [7:0] _GEN_7855 = opcode_7 != 4'h0 ? _GEN_7507 : _GEN_7087; // @[executor.scala 470:55]
  wire [7:0] _GEN_7856 = opcode_7 != 4'h0 ? _GEN_7508 : _GEN_7088; // @[executor.scala 470:55]
  wire [7:0] _GEN_7857 = opcode_7 != 4'h0 ? _GEN_7509 : _GEN_7089; // @[executor.scala 470:55]
  wire [7:0] _GEN_7858 = opcode_7 != 4'h0 ? _GEN_7514 : _GEN_7090; // @[executor.scala 470:55]
  wire [7:0] _GEN_7859 = opcode_7 != 4'h0 ? _GEN_7515 : _GEN_7091; // @[executor.scala 470:55]
  wire [7:0] _GEN_7860 = opcode_7 != 4'h0 ? _GEN_7516 : _GEN_7092; // @[executor.scala 470:55]
  wire [7:0] _GEN_7861 = opcode_7 != 4'h0 ? _GEN_7517 : _GEN_7093; // @[executor.scala 470:55]
  wire [7:0] _GEN_7862 = opcode_7 != 4'h0 ? _GEN_7522 : _GEN_7094; // @[executor.scala 470:55]
  wire [7:0] _GEN_7863 = opcode_7 != 4'h0 ? _GEN_7523 : _GEN_7095; // @[executor.scala 470:55]
  wire [7:0] _GEN_7864 = opcode_7 != 4'h0 ? _GEN_7524 : _GEN_7096; // @[executor.scala 470:55]
  wire [7:0] _GEN_7865 = opcode_7 != 4'h0 ? _GEN_7525 : _GEN_7097; // @[executor.scala 470:55]
  wire [7:0] _GEN_7866 = opcode_7 != 4'h0 ? _GEN_7530 : _GEN_7098; // @[executor.scala 470:55]
  wire [7:0] _GEN_7867 = opcode_7 != 4'h0 ? _GEN_7531 : _GEN_7099; // @[executor.scala 470:55]
  wire [7:0] _GEN_7868 = opcode_7 != 4'h0 ? _GEN_7532 : _GEN_7100; // @[executor.scala 470:55]
  wire [7:0] _GEN_7869 = opcode_7 != 4'h0 ? _GEN_7533 : _GEN_7101; // @[executor.scala 470:55]
  wire [7:0] _GEN_7870 = opcode_7 != 4'h0 ? _GEN_7538 : _GEN_7102; // @[executor.scala 470:55]
  wire [7:0] _GEN_7871 = opcode_7 != 4'h0 ? _GEN_7539 : _GEN_7103; // @[executor.scala 470:55]
  wire [7:0] _GEN_7872 = opcode_7 != 4'h0 ? _GEN_7540 : _GEN_7104; // @[executor.scala 470:55]
  wire [7:0] _GEN_7873 = opcode_7 != 4'h0 ? _GEN_7541 : _GEN_7105; // @[executor.scala 470:55]
  wire [7:0] _GEN_7874 = opcode_7 != 4'h0 ? _GEN_7546 : _GEN_7106; // @[executor.scala 470:55]
  wire [7:0] _GEN_7875 = opcode_7 != 4'h0 ? _GEN_7547 : _GEN_7107; // @[executor.scala 470:55]
  wire [7:0] _GEN_7876 = opcode_7 != 4'h0 ? _GEN_7548 : _GEN_7108; // @[executor.scala 470:55]
  wire [7:0] _GEN_7877 = opcode_7 != 4'h0 ? _GEN_7549 : _GEN_7109; // @[executor.scala 470:55]
  wire [7:0] _GEN_7878 = opcode_7 != 4'h0 ? _GEN_7554 : _GEN_7110; // @[executor.scala 470:55]
  wire [7:0] _GEN_7879 = opcode_7 != 4'h0 ? _GEN_7555 : _GEN_7111; // @[executor.scala 470:55]
  wire [7:0] _GEN_7880 = opcode_7 != 4'h0 ? _GEN_7556 : _GEN_7112; // @[executor.scala 470:55]
  wire [7:0] _GEN_7881 = opcode_7 != 4'h0 ? _GEN_7557 : _GEN_7113; // @[executor.scala 470:55]
  wire [7:0] _GEN_7882 = opcode_7 != 4'h0 ? _GEN_7562 : _GEN_7114; // @[executor.scala 470:55]
  wire [7:0] _GEN_7883 = opcode_7 != 4'h0 ? _GEN_7563 : _GEN_7115; // @[executor.scala 470:55]
  wire [7:0] _GEN_7884 = opcode_7 != 4'h0 ? _GEN_7564 : _GEN_7116; // @[executor.scala 470:55]
  wire [7:0] _GEN_7885 = opcode_7 != 4'h0 ? _GEN_7565 : _GEN_7117; // @[executor.scala 470:55]
  wire [7:0] _GEN_7886 = opcode_7 != 4'h0 ? _GEN_7570 : _GEN_7118; // @[executor.scala 470:55]
  wire [7:0] _GEN_7887 = opcode_7 != 4'h0 ? _GEN_7571 : _GEN_7119; // @[executor.scala 470:55]
  wire [7:0] _GEN_7888 = opcode_7 != 4'h0 ? _GEN_7572 : _GEN_7120; // @[executor.scala 470:55]
  wire [7:0] _GEN_7889 = opcode_7 != 4'h0 ? _GEN_7573 : _GEN_7121; // @[executor.scala 470:55]
  wire [7:0] _GEN_7890 = opcode_7 != 4'h0 ? _GEN_7578 : _GEN_7122; // @[executor.scala 470:55]
  wire [7:0] _GEN_7891 = opcode_7 != 4'h0 ? _GEN_7579 : _GEN_7123; // @[executor.scala 470:55]
  wire [7:0] _GEN_7892 = opcode_7 != 4'h0 ? _GEN_7580 : _GEN_7124; // @[executor.scala 470:55]
  wire [7:0] _GEN_7893 = opcode_7 != 4'h0 ? _GEN_7581 : _GEN_7125; // @[executor.scala 470:55]
  wire [7:0] _GEN_7894 = opcode_7 != 4'h0 ? _GEN_7586 : _GEN_7126; // @[executor.scala 470:55]
  wire [7:0] _GEN_7895 = opcode_7 != 4'h0 ? _GEN_7587 : _GEN_7127; // @[executor.scala 470:55]
  wire [7:0] _GEN_7896 = opcode_7 != 4'h0 ? _GEN_7588 : _GEN_7128; // @[executor.scala 470:55]
  wire [7:0] _GEN_7897 = opcode_7 != 4'h0 ? _GEN_7589 : _GEN_7129; // @[executor.scala 470:55]
  wire [7:0] _GEN_7898 = opcode_7 != 4'h0 ? _GEN_7594 : _GEN_7130; // @[executor.scala 470:55]
  wire [7:0] _GEN_7899 = opcode_7 != 4'h0 ? _GEN_7595 : _GEN_7131; // @[executor.scala 470:55]
  wire [7:0] _GEN_7900 = opcode_7 != 4'h0 ? _GEN_7596 : _GEN_7132; // @[executor.scala 470:55]
  wire [7:0] _GEN_7901 = opcode_7 != 4'h0 ? _GEN_7597 : _GEN_7133; // @[executor.scala 470:55]
  wire [7:0] _GEN_7902 = opcode_7 != 4'h0 ? _GEN_7602 : _GEN_7134; // @[executor.scala 470:55]
  wire [7:0] _GEN_7903 = opcode_7 != 4'h0 ? _GEN_7603 : _GEN_7135; // @[executor.scala 470:55]
  wire [7:0] _GEN_7904 = opcode_7 != 4'h0 ? _GEN_7604 : _GEN_7136; // @[executor.scala 470:55]
  wire [7:0] _GEN_7905 = opcode_7 != 4'h0 ? _GEN_7605 : _GEN_7137; // @[executor.scala 470:55]
  wire [7:0] _GEN_7906 = opcode_7 != 4'h0 ? _GEN_7610 : _GEN_7138; // @[executor.scala 470:55]
  wire [7:0] _GEN_7907 = opcode_7 != 4'h0 ? _GEN_7611 : _GEN_7139; // @[executor.scala 470:55]
  wire [7:0] _GEN_7908 = opcode_7 != 4'h0 ? _GEN_7612 : _GEN_7140; // @[executor.scala 470:55]
  wire [7:0] _GEN_7909 = opcode_7 != 4'h0 ? _GEN_7613 : _GEN_7141; // @[executor.scala 470:55]
  wire [7:0] _GEN_7910 = opcode_7 != 4'h0 ? _GEN_7618 : _GEN_7142; // @[executor.scala 470:55]
  wire [7:0] _GEN_7911 = opcode_7 != 4'h0 ? _GEN_7619 : _GEN_7143; // @[executor.scala 470:55]
  wire [7:0] _GEN_7912 = opcode_7 != 4'h0 ? _GEN_7620 : _GEN_7144; // @[executor.scala 470:55]
  wire [7:0] _GEN_7913 = opcode_7 != 4'h0 ? _GEN_7621 : _GEN_7145; // @[executor.scala 470:55]
  wire [7:0] _GEN_7914 = opcode_7 != 4'h0 ? _GEN_7626 : _GEN_7146; // @[executor.scala 470:55]
  wire [7:0] _GEN_7915 = opcode_7 != 4'h0 ? _GEN_7627 : _GEN_7147; // @[executor.scala 470:55]
  wire [7:0] _GEN_7916 = opcode_7 != 4'h0 ? _GEN_7628 : _GEN_7148; // @[executor.scala 470:55]
  wire [7:0] _GEN_7917 = opcode_7 != 4'h0 ? _GEN_7629 : _GEN_7149; // @[executor.scala 470:55]
  wire [7:0] _GEN_7918 = opcode_7 != 4'h0 ? _GEN_7634 : _GEN_7150; // @[executor.scala 470:55]
  wire [7:0] _GEN_7919 = opcode_7 != 4'h0 ? _GEN_7635 : _GEN_7151; // @[executor.scala 470:55]
  wire [7:0] _GEN_7920 = opcode_7 != 4'h0 ? _GEN_7636 : _GEN_7152; // @[executor.scala 470:55]
  wire [7:0] _GEN_7921 = opcode_7 != 4'h0 ? _GEN_7637 : _GEN_7153; // @[executor.scala 470:55]
  wire [7:0] _GEN_7922 = opcode_7 != 4'h0 ? _GEN_7642 : _GEN_7154; // @[executor.scala 470:55]
  wire [7:0] _GEN_7923 = opcode_7 != 4'h0 ? _GEN_7643 : _GEN_7155; // @[executor.scala 470:55]
  wire [7:0] _GEN_7924 = opcode_7 != 4'h0 ? _GEN_7644 : _GEN_7156; // @[executor.scala 470:55]
  wire [7:0] _GEN_7925 = opcode_7 != 4'h0 ? _GEN_7645 : _GEN_7157; // @[executor.scala 470:55]
  wire [7:0] _GEN_7926 = opcode_7 != 4'h0 ? _GEN_7650 : _GEN_7158; // @[executor.scala 470:55]
  wire [7:0] _GEN_7927 = opcode_7 != 4'h0 ? _GEN_7651 : _GEN_7159; // @[executor.scala 470:55]
  wire [7:0] _GEN_7928 = opcode_7 != 4'h0 ? _GEN_7652 : _GEN_7160; // @[executor.scala 470:55]
  wire [7:0] _GEN_7929 = opcode_7 != 4'h0 ? _GEN_7653 : _GEN_7161; // @[executor.scala 470:55]
  wire [7:0] _GEN_7930 = opcode_7 != 4'h0 ? _GEN_7658 : _GEN_7162; // @[executor.scala 470:55]
  wire [7:0] _GEN_7931 = opcode_7 != 4'h0 ? _GEN_7659 : _GEN_7163; // @[executor.scala 470:55]
  wire [7:0] _GEN_7932 = opcode_7 != 4'h0 ? _GEN_7660 : _GEN_7164; // @[executor.scala 470:55]
  wire [7:0] _GEN_7933 = opcode_7 != 4'h0 ? _GEN_7661 : _GEN_7165; // @[executor.scala 470:55]
  wire [7:0] _GEN_7934 = opcode_7 != 4'h0 ? _GEN_7666 : _GEN_7166; // @[executor.scala 470:55]
  wire [7:0] _GEN_7935 = opcode_7 != 4'h0 ? _GEN_7667 : _GEN_7167; // @[executor.scala 470:55]
  wire [7:0] _GEN_7936 = opcode_7 != 4'h0 ? _GEN_7668 : _GEN_7168; // @[executor.scala 470:55]
  wire [7:0] _GEN_7937 = opcode_7 != 4'h0 ? _GEN_7669 : _GEN_7169; // @[executor.scala 470:55]
  wire [7:0] _GEN_7938 = opcode_7 != 4'h0 ? _GEN_7674 : _GEN_7170; // @[executor.scala 470:55]
  wire [7:0] _GEN_7939 = opcode_7 != 4'h0 ? _GEN_7675 : _GEN_7171; // @[executor.scala 470:55]
  wire [7:0] _GEN_7940 = opcode_7 != 4'h0 ? _GEN_7676 : _GEN_7172; // @[executor.scala 470:55]
  wire [7:0] _GEN_7941 = opcode_7 != 4'h0 ? _GEN_7677 : _GEN_7173; // @[executor.scala 470:55]
  wire [7:0] _GEN_7942 = opcode_7 != 4'h0 ? _GEN_7682 : _GEN_7174; // @[executor.scala 470:55]
  wire [7:0] _GEN_7943 = opcode_7 != 4'h0 ? _GEN_7683 : _GEN_7175; // @[executor.scala 470:55]
  wire [7:0] _GEN_7944 = opcode_7 != 4'h0 ? _GEN_7684 : _GEN_7176; // @[executor.scala 470:55]
  wire [7:0] _GEN_7945 = opcode_7 != 4'h0 ? _GEN_7685 : _GEN_7177; // @[executor.scala 470:55]
  wire [7:0] _GEN_7946 = opcode_7 != 4'h0 ? _GEN_7690 : _GEN_7178; // @[executor.scala 470:55]
  wire [7:0] _GEN_7947 = opcode_7 != 4'h0 ? _GEN_7691 : _GEN_7179; // @[executor.scala 470:55]
  wire [7:0] _GEN_7948 = opcode_7 != 4'h0 ? _GEN_7692 : _GEN_7180; // @[executor.scala 470:55]
  wire [7:0] _GEN_7949 = opcode_7 != 4'h0 ? _GEN_7693 : _GEN_7181; // @[executor.scala 470:55]
  wire [3:0] _GEN_7950 = opcode_7 == 4'hf ? parameter_2_7[13:10] : _GEN_6924; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_7951 = opcode_7 == 4'hf ? parameter_2_7[0] : _GEN_6925; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_7952 = opcode_7 == 4'hf ? _GEN_6926 : _GEN_7694; // @[executor.scala 466:52]
  wire [7:0] _GEN_7953 = opcode_7 == 4'hf ? _GEN_6927 : _GEN_7695; // @[executor.scala 466:52]
  wire [7:0] _GEN_7954 = opcode_7 == 4'hf ? _GEN_6928 : _GEN_7696; // @[executor.scala 466:52]
  wire [7:0] _GEN_7955 = opcode_7 == 4'hf ? _GEN_6929 : _GEN_7697; // @[executor.scala 466:52]
  wire [7:0] _GEN_7956 = opcode_7 == 4'hf ? _GEN_6930 : _GEN_7698; // @[executor.scala 466:52]
  wire [7:0] _GEN_7957 = opcode_7 == 4'hf ? _GEN_6931 : _GEN_7699; // @[executor.scala 466:52]
  wire [7:0] _GEN_7958 = opcode_7 == 4'hf ? _GEN_6932 : _GEN_7700; // @[executor.scala 466:52]
  wire [7:0] _GEN_7959 = opcode_7 == 4'hf ? _GEN_6933 : _GEN_7701; // @[executor.scala 466:52]
  wire [7:0] _GEN_7960 = opcode_7 == 4'hf ? _GEN_6934 : _GEN_7702; // @[executor.scala 466:52]
  wire [7:0] _GEN_7961 = opcode_7 == 4'hf ? _GEN_6935 : _GEN_7703; // @[executor.scala 466:52]
  wire [7:0] _GEN_7962 = opcode_7 == 4'hf ? _GEN_6936 : _GEN_7704; // @[executor.scala 466:52]
  wire [7:0] _GEN_7963 = opcode_7 == 4'hf ? _GEN_6937 : _GEN_7705; // @[executor.scala 466:52]
  wire [7:0] _GEN_7964 = opcode_7 == 4'hf ? _GEN_6938 : _GEN_7706; // @[executor.scala 466:52]
  wire [7:0] _GEN_7965 = opcode_7 == 4'hf ? _GEN_6939 : _GEN_7707; // @[executor.scala 466:52]
  wire [7:0] _GEN_7966 = opcode_7 == 4'hf ? _GEN_6940 : _GEN_7708; // @[executor.scala 466:52]
  wire [7:0] _GEN_7967 = opcode_7 == 4'hf ? _GEN_6941 : _GEN_7709; // @[executor.scala 466:52]
  wire [7:0] _GEN_7968 = opcode_7 == 4'hf ? _GEN_6942 : _GEN_7710; // @[executor.scala 466:52]
  wire [7:0] _GEN_7969 = opcode_7 == 4'hf ? _GEN_6943 : _GEN_7711; // @[executor.scala 466:52]
  wire [7:0] _GEN_7970 = opcode_7 == 4'hf ? _GEN_6944 : _GEN_7712; // @[executor.scala 466:52]
  wire [7:0] _GEN_7971 = opcode_7 == 4'hf ? _GEN_6945 : _GEN_7713; // @[executor.scala 466:52]
  wire [7:0] _GEN_7972 = opcode_7 == 4'hf ? _GEN_6946 : _GEN_7714; // @[executor.scala 466:52]
  wire [7:0] _GEN_7973 = opcode_7 == 4'hf ? _GEN_6947 : _GEN_7715; // @[executor.scala 466:52]
  wire [7:0] _GEN_7974 = opcode_7 == 4'hf ? _GEN_6948 : _GEN_7716; // @[executor.scala 466:52]
  wire [7:0] _GEN_7975 = opcode_7 == 4'hf ? _GEN_6949 : _GEN_7717; // @[executor.scala 466:52]
  wire [7:0] _GEN_7976 = opcode_7 == 4'hf ? _GEN_6950 : _GEN_7718; // @[executor.scala 466:52]
  wire [7:0] _GEN_7977 = opcode_7 == 4'hf ? _GEN_6951 : _GEN_7719; // @[executor.scala 466:52]
  wire [7:0] _GEN_7978 = opcode_7 == 4'hf ? _GEN_6952 : _GEN_7720; // @[executor.scala 466:52]
  wire [7:0] _GEN_7979 = opcode_7 == 4'hf ? _GEN_6953 : _GEN_7721; // @[executor.scala 466:52]
  wire [7:0] _GEN_7980 = opcode_7 == 4'hf ? _GEN_6954 : _GEN_7722; // @[executor.scala 466:52]
  wire [7:0] _GEN_7981 = opcode_7 == 4'hf ? _GEN_6955 : _GEN_7723; // @[executor.scala 466:52]
  wire [7:0] _GEN_7982 = opcode_7 == 4'hf ? _GEN_6956 : _GEN_7724; // @[executor.scala 466:52]
  wire [7:0] _GEN_7983 = opcode_7 == 4'hf ? _GEN_6957 : _GEN_7725; // @[executor.scala 466:52]
  wire [7:0] _GEN_7984 = opcode_7 == 4'hf ? _GEN_6958 : _GEN_7726; // @[executor.scala 466:52]
  wire [7:0] _GEN_7985 = opcode_7 == 4'hf ? _GEN_6959 : _GEN_7727; // @[executor.scala 466:52]
  wire [7:0] _GEN_7986 = opcode_7 == 4'hf ? _GEN_6960 : _GEN_7728; // @[executor.scala 466:52]
  wire [7:0] _GEN_7987 = opcode_7 == 4'hf ? _GEN_6961 : _GEN_7729; // @[executor.scala 466:52]
  wire [7:0] _GEN_7988 = opcode_7 == 4'hf ? _GEN_6962 : _GEN_7730; // @[executor.scala 466:52]
  wire [7:0] _GEN_7989 = opcode_7 == 4'hf ? _GEN_6963 : _GEN_7731; // @[executor.scala 466:52]
  wire [7:0] _GEN_7990 = opcode_7 == 4'hf ? _GEN_6964 : _GEN_7732; // @[executor.scala 466:52]
  wire [7:0] _GEN_7991 = opcode_7 == 4'hf ? _GEN_6965 : _GEN_7733; // @[executor.scala 466:52]
  wire [7:0] _GEN_7992 = opcode_7 == 4'hf ? _GEN_6966 : _GEN_7734; // @[executor.scala 466:52]
  wire [7:0] _GEN_7993 = opcode_7 == 4'hf ? _GEN_6967 : _GEN_7735; // @[executor.scala 466:52]
  wire [7:0] _GEN_7994 = opcode_7 == 4'hf ? _GEN_6968 : _GEN_7736; // @[executor.scala 466:52]
  wire [7:0] _GEN_7995 = opcode_7 == 4'hf ? _GEN_6969 : _GEN_7737; // @[executor.scala 466:52]
  wire [7:0] _GEN_7996 = opcode_7 == 4'hf ? _GEN_6970 : _GEN_7738; // @[executor.scala 466:52]
  wire [7:0] _GEN_7997 = opcode_7 == 4'hf ? _GEN_6971 : _GEN_7739; // @[executor.scala 466:52]
  wire [7:0] _GEN_7998 = opcode_7 == 4'hf ? _GEN_6972 : _GEN_7740; // @[executor.scala 466:52]
  wire [7:0] _GEN_7999 = opcode_7 == 4'hf ? _GEN_6973 : _GEN_7741; // @[executor.scala 466:52]
  wire [7:0] _GEN_8000 = opcode_7 == 4'hf ? _GEN_6974 : _GEN_7742; // @[executor.scala 466:52]
  wire [7:0] _GEN_8001 = opcode_7 == 4'hf ? _GEN_6975 : _GEN_7743; // @[executor.scala 466:52]
  wire [7:0] _GEN_8002 = opcode_7 == 4'hf ? _GEN_6976 : _GEN_7744; // @[executor.scala 466:52]
  wire [7:0] _GEN_8003 = opcode_7 == 4'hf ? _GEN_6977 : _GEN_7745; // @[executor.scala 466:52]
  wire [7:0] _GEN_8004 = opcode_7 == 4'hf ? _GEN_6978 : _GEN_7746; // @[executor.scala 466:52]
  wire [7:0] _GEN_8005 = opcode_7 == 4'hf ? _GEN_6979 : _GEN_7747; // @[executor.scala 466:52]
  wire [7:0] _GEN_8006 = opcode_7 == 4'hf ? _GEN_6980 : _GEN_7748; // @[executor.scala 466:52]
  wire [7:0] _GEN_8007 = opcode_7 == 4'hf ? _GEN_6981 : _GEN_7749; // @[executor.scala 466:52]
  wire [7:0] _GEN_8008 = opcode_7 == 4'hf ? _GEN_6982 : _GEN_7750; // @[executor.scala 466:52]
  wire [7:0] _GEN_8009 = opcode_7 == 4'hf ? _GEN_6983 : _GEN_7751; // @[executor.scala 466:52]
  wire [7:0] _GEN_8010 = opcode_7 == 4'hf ? _GEN_6984 : _GEN_7752; // @[executor.scala 466:52]
  wire [7:0] _GEN_8011 = opcode_7 == 4'hf ? _GEN_6985 : _GEN_7753; // @[executor.scala 466:52]
  wire [7:0] _GEN_8012 = opcode_7 == 4'hf ? _GEN_6986 : _GEN_7754; // @[executor.scala 466:52]
  wire [7:0] _GEN_8013 = opcode_7 == 4'hf ? _GEN_6987 : _GEN_7755; // @[executor.scala 466:52]
  wire [7:0] _GEN_8014 = opcode_7 == 4'hf ? _GEN_6988 : _GEN_7756; // @[executor.scala 466:52]
  wire [7:0] _GEN_8015 = opcode_7 == 4'hf ? _GEN_6989 : _GEN_7757; // @[executor.scala 466:52]
  wire [7:0] _GEN_8016 = opcode_7 == 4'hf ? _GEN_6990 : _GEN_7758; // @[executor.scala 466:52]
  wire [7:0] _GEN_8017 = opcode_7 == 4'hf ? _GEN_6991 : _GEN_7759; // @[executor.scala 466:52]
  wire [7:0] _GEN_8018 = opcode_7 == 4'hf ? _GEN_6992 : _GEN_7760; // @[executor.scala 466:52]
  wire [7:0] _GEN_8019 = opcode_7 == 4'hf ? _GEN_6993 : _GEN_7761; // @[executor.scala 466:52]
  wire [7:0] _GEN_8020 = opcode_7 == 4'hf ? _GEN_6994 : _GEN_7762; // @[executor.scala 466:52]
  wire [7:0] _GEN_8021 = opcode_7 == 4'hf ? _GEN_6995 : _GEN_7763; // @[executor.scala 466:52]
  wire [7:0] _GEN_8022 = opcode_7 == 4'hf ? _GEN_6996 : _GEN_7764; // @[executor.scala 466:52]
  wire [7:0] _GEN_8023 = opcode_7 == 4'hf ? _GEN_6997 : _GEN_7765; // @[executor.scala 466:52]
  wire [7:0] _GEN_8024 = opcode_7 == 4'hf ? _GEN_6998 : _GEN_7766; // @[executor.scala 466:52]
  wire [7:0] _GEN_8025 = opcode_7 == 4'hf ? _GEN_6999 : _GEN_7767; // @[executor.scala 466:52]
  wire [7:0] _GEN_8026 = opcode_7 == 4'hf ? _GEN_7000 : _GEN_7768; // @[executor.scala 466:52]
  wire [7:0] _GEN_8027 = opcode_7 == 4'hf ? _GEN_7001 : _GEN_7769; // @[executor.scala 466:52]
  wire [7:0] _GEN_8028 = opcode_7 == 4'hf ? _GEN_7002 : _GEN_7770; // @[executor.scala 466:52]
  wire [7:0] _GEN_8029 = opcode_7 == 4'hf ? _GEN_7003 : _GEN_7771; // @[executor.scala 466:52]
  wire [7:0] _GEN_8030 = opcode_7 == 4'hf ? _GEN_7004 : _GEN_7772; // @[executor.scala 466:52]
  wire [7:0] _GEN_8031 = opcode_7 == 4'hf ? _GEN_7005 : _GEN_7773; // @[executor.scala 466:52]
  wire [7:0] _GEN_8032 = opcode_7 == 4'hf ? _GEN_7006 : _GEN_7774; // @[executor.scala 466:52]
  wire [7:0] _GEN_8033 = opcode_7 == 4'hf ? _GEN_7007 : _GEN_7775; // @[executor.scala 466:52]
  wire [7:0] _GEN_8034 = opcode_7 == 4'hf ? _GEN_7008 : _GEN_7776; // @[executor.scala 466:52]
  wire [7:0] _GEN_8035 = opcode_7 == 4'hf ? _GEN_7009 : _GEN_7777; // @[executor.scala 466:52]
  wire [7:0] _GEN_8036 = opcode_7 == 4'hf ? _GEN_7010 : _GEN_7778; // @[executor.scala 466:52]
  wire [7:0] _GEN_8037 = opcode_7 == 4'hf ? _GEN_7011 : _GEN_7779; // @[executor.scala 466:52]
  wire [7:0] _GEN_8038 = opcode_7 == 4'hf ? _GEN_7012 : _GEN_7780; // @[executor.scala 466:52]
  wire [7:0] _GEN_8039 = opcode_7 == 4'hf ? _GEN_7013 : _GEN_7781; // @[executor.scala 466:52]
  wire [7:0] _GEN_8040 = opcode_7 == 4'hf ? _GEN_7014 : _GEN_7782; // @[executor.scala 466:52]
  wire [7:0] _GEN_8041 = opcode_7 == 4'hf ? _GEN_7015 : _GEN_7783; // @[executor.scala 466:52]
  wire [7:0] _GEN_8042 = opcode_7 == 4'hf ? _GEN_7016 : _GEN_7784; // @[executor.scala 466:52]
  wire [7:0] _GEN_8043 = opcode_7 == 4'hf ? _GEN_7017 : _GEN_7785; // @[executor.scala 466:52]
  wire [7:0] _GEN_8044 = opcode_7 == 4'hf ? _GEN_7018 : _GEN_7786; // @[executor.scala 466:52]
  wire [7:0] _GEN_8045 = opcode_7 == 4'hf ? _GEN_7019 : _GEN_7787; // @[executor.scala 466:52]
  wire [7:0] _GEN_8046 = opcode_7 == 4'hf ? _GEN_7020 : _GEN_7788; // @[executor.scala 466:52]
  wire [7:0] _GEN_8047 = opcode_7 == 4'hf ? _GEN_7021 : _GEN_7789; // @[executor.scala 466:52]
  wire [7:0] _GEN_8048 = opcode_7 == 4'hf ? _GEN_7022 : _GEN_7790; // @[executor.scala 466:52]
  wire [7:0] _GEN_8049 = opcode_7 == 4'hf ? _GEN_7023 : _GEN_7791; // @[executor.scala 466:52]
  wire [7:0] _GEN_8050 = opcode_7 == 4'hf ? _GEN_7024 : _GEN_7792; // @[executor.scala 466:52]
  wire [7:0] _GEN_8051 = opcode_7 == 4'hf ? _GEN_7025 : _GEN_7793; // @[executor.scala 466:52]
  wire [7:0] _GEN_8052 = opcode_7 == 4'hf ? _GEN_7026 : _GEN_7794; // @[executor.scala 466:52]
  wire [7:0] _GEN_8053 = opcode_7 == 4'hf ? _GEN_7027 : _GEN_7795; // @[executor.scala 466:52]
  wire [7:0] _GEN_8054 = opcode_7 == 4'hf ? _GEN_7028 : _GEN_7796; // @[executor.scala 466:52]
  wire [7:0] _GEN_8055 = opcode_7 == 4'hf ? _GEN_7029 : _GEN_7797; // @[executor.scala 466:52]
  wire [7:0] _GEN_8056 = opcode_7 == 4'hf ? _GEN_7030 : _GEN_7798; // @[executor.scala 466:52]
  wire [7:0] _GEN_8057 = opcode_7 == 4'hf ? _GEN_7031 : _GEN_7799; // @[executor.scala 466:52]
  wire [7:0] _GEN_8058 = opcode_7 == 4'hf ? _GEN_7032 : _GEN_7800; // @[executor.scala 466:52]
  wire [7:0] _GEN_8059 = opcode_7 == 4'hf ? _GEN_7033 : _GEN_7801; // @[executor.scala 466:52]
  wire [7:0] _GEN_8060 = opcode_7 == 4'hf ? _GEN_7034 : _GEN_7802; // @[executor.scala 466:52]
  wire [7:0] _GEN_8061 = opcode_7 == 4'hf ? _GEN_7035 : _GEN_7803; // @[executor.scala 466:52]
  wire [7:0] _GEN_8062 = opcode_7 == 4'hf ? _GEN_7036 : _GEN_7804; // @[executor.scala 466:52]
  wire [7:0] _GEN_8063 = opcode_7 == 4'hf ? _GEN_7037 : _GEN_7805; // @[executor.scala 466:52]
  wire [7:0] _GEN_8064 = opcode_7 == 4'hf ? _GEN_7038 : _GEN_7806; // @[executor.scala 466:52]
  wire [7:0] _GEN_8065 = opcode_7 == 4'hf ? _GEN_7039 : _GEN_7807; // @[executor.scala 466:52]
  wire [7:0] _GEN_8066 = opcode_7 == 4'hf ? _GEN_7040 : _GEN_7808; // @[executor.scala 466:52]
  wire [7:0] _GEN_8067 = opcode_7 == 4'hf ? _GEN_7041 : _GEN_7809; // @[executor.scala 466:52]
  wire [7:0] _GEN_8068 = opcode_7 == 4'hf ? _GEN_7042 : _GEN_7810; // @[executor.scala 466:52]
  wire [7:0] _GEN_8069 = opcode_7 == 4'hf ? _GEN_7043 : _GEN_7811; // @[executor.scala 466:52]
  wire [7:0] _GEN_8070 = opcode_7 == 4'hf ? _GEN_7044 : _GEN_7812; // @[executor.scala 466:52]
  wire [7:0] _GEN_8071 = opcode_7 == 4'hf ? _GEN_7045 : _GEN_7813; // @[executor.scala 466:52]
  wire [7:0] _GEN_8072 = opcode_7 == 4'hf ? _GEN_7046 : _GEN_7814; // @[executor.scala 466:52]
  wire [7:0] _GEN_8073 = opcode_7 == 4'hf ? _GEN_7047 : _GEN_7815; // @[executor.scala 466:52]
  wire [7:0] _GEN_8074 = opcode_7 == 4'hf ? _GEN_7048 : _GEN_7816; // @[executor.scala 466:52]
  wire [7:0] _GEN_8075 = opcode_7 == 4'hf ? _GEN_7049 : _GEN_7817; // @[executor.scala 466:52]
  wire [7:0] _GEN_8076 = opcode_7 == 4'hf ? _GEN_7050 : _GEN_7818; // @[executor.scala 466:52]
  wire [7:0] _GEN_8077 = opcode_7 == 4'hf ? _GEN_7051 : _GEN_7819; // @[executor.scala 466:52]
  wire [7:0] _GEN_8078 = opcode_7 == 4'hf ? _GEN_7052 : _GEN_7820; // @[executor.scala 466:52]
  wire [7:0] _GEN_8079 = opcode_7 == 4'hf ? _GEN_7053 : _GEN_7821; // @[executor.scala 466:52]
  wire [7:0] _GEN_8080 = opcode_7 == 4'hf ? _GEN_7054 : _GEN_7822; // @[executor.scala 466:52]
  wire [7:0] _GEN_8081 = opcode_7 == 4'hf ? _GEN_7055 : _GEN_7823; // @[executor.scala 466:52]
  wire [7:0] _GEN_8082 = opcode_7 == 4'hf ? _GEN_7056 : _GEN_7824; // @[executor.scala 466:52]
  wire [7:0] _GEN_8083 = opcode_7 == 4'hf ? _GEN_7057 : _GEN_7825; // @[executor.scala 466:52]
  wire [7:0] _GEN_8084 = opcode_7 == 4'hf ? _GEN_7058 : _GEN_7826; // @[executor.scala 466:52]
  wire [7:0] _GEN_8085 = opcode_7 == 4'hf ? _GEN_7059 : _GEN_7827; // @[executor.scala 466:52]
  wire [7:0] _GEN_8086 = opcode_7 == 4'hf ? _GEN_7060 : _GEN_7828; // @[executor.scala 466:52]
  wire [7:0] _GEN_8087 = opcode_7 == 4'hf ? _GEN_7061 : _GEN_7829; // @[executor.scala 466:52]
  wire [7:0] _GEN_8088 = opcode_7 == 4'hf ? _GEN_7062 : _GEN_7830; // @[executor.scala 466:52]
  wire [7:0] _GEN_8089 = opcode_7 == 4'hf ? _GEN_7063 : _GEN_7831; // @[executor.scala 466:52]
  wire [7:0] _GEN_8090 = opcode_7 == 4'hf ? _GEN_7064 : _GEN_7832; // @[executor.scala 466:52]
  wire [7:0] _GEN_8091 = opcode_7 == 4'hf ? _GEN_7065 : _GEN_7833; // @[executor.scala 466:52]
  wire [7:0] _GEN_8092 = opcode_7 == 4'hf ? _GEN_7066 : _GEN_7834; // @[executor.scala 466:52]
  wire [7:0] _GEN_8093 = opcode_7 == 4'hf ? _GEN_7067 : _GEN_7835; // @[executor.scala 466:52]
  wire [7:0] _GEN_8094 = opcode_7 == 4'hf ? _GEN_7068 : _GEN_7836; // @[executor.scala 466:52]
  wire [7:0] _GEN_8095 = opcode_7 == 4'hf ? _GEN_7069 : _GEN_7837; // @[executor.scala 466:52]
  wire [7:0] _GEN_8096 = opcode_7 == 4'hf ? _GEN_7070 : _GEN_7838; // @[executor.scala 466:52]
  wire [7:0] _GEN_8097 = opcode_7 == 4'hf ? _GEN_7071 : _GEN_7839; // @[executor.scala 466:52]
  wire [7:0] _GEN_8098 = opcode_7 == 4'hf ? _GEN_7072 : _GEN_7840; // @[executor.scala 466:52]
  wire [7:0] _GEN_8099 = opcode_7 == 4'hf ? _GEN_7073 : _GEN_7841; // @[executor.scala 466:52]
  wire [7:0] _GEN_8100 = opcode_7 == 4'hf ? _GEN_7074 : _GEN_7842; // @[executor.scala 466:52]
  wire [7:0] _GEN_8101 = opcode_7 == 4'hf ? _GEN_7075 : _GEN_7843; // @[executor.scala 466:52]
  wire [7:0] _GEN_8102 = opcode_7 == 4'hf ? _GEN_7076 : _GEN_7844; // @[executor.scala 466:52]
  wire [7:0] _GEN_8103 = opcode_7 == 4'hf ? _GEN_7077 : _GEN_7845; // @[executor.scala 466:52]
  wire [7:0] _GEN_8104 = opcode_7 == 4'hf ? _GEN_7078 : _GEN_7846; // @[executor.scala 466:52]
  wire [7:0] _GEN_8105 = opcode_7 == 4'hf ? _GEN_7079 : _GEN_7847; // @[executor.scala 466:52]
  wire [7:0] _GEN_8106 = opcode_7 == 4'hf ? _GEN_7080 : _GEN_7848; // @[executor.scala 466:52]
  wire [7:0] _GEN_8107 = opcode_7 == 4'hf ? _GEN_7081 : _GEN_7849; // @[executor.scala 466:52]
  wire [7:0] _GEN_8108 = opcode_7 == 4'hf ? _GEN_7082 : _GEN_7850; // @[executor.scala 466:52]
  wire [7:0] _GEN_8109 = opcode_7 == 4'hf ? _GEN_7083 : _GEN_7851; // @[executor.scala 466:52]
  wire [7:0] _GEN_8110 = opcode_7 == 4'hf ? _GEN_7084 : _GEN_7852; // @[executor.scala 466:52]
  wire [7:0] _GEN_8111 = opcode_7 == 4'hf ? _GEN_7085 : _GEN_7853; // @[executor.scala 466:52]
  wire [7:0] _GEN_8112 = opcode_7 == 4'hf ? _GEN_7086 : _GEN_7854; // @[executor.scala 466:52]
  wire [7:0] _GEN_8113 = opcode_7 == 4'hf ? _GEN_7087 : _GEN_7855; // @[executor.scala 466:52]
  wire [7:0] _GEN_8114 = opcode_7 == 4'hf ? _GEN_7088 : _GEN_7856; // @[executor.scala 466:52]
  wire [7:0] _GEN_8115 = opcode_7 == 4'hf ? _GEN_7089 : _GEN_7857; // @[executor.scala 466:52]
  wire [7:0] _GEN_8116 = opcode_7 == 4'hf ? _GEN_7090 : _GEN_7858; // @[executor.scala 466:52]
  wire [7:0] _GEN_8117 = opcode_7 == 4'hf ? _GEN_7091 : _GEN_7859; // @[executor.scala 466:52]
  wire [7:0] _GEN_8118 = opcode_7 == 4'hf ? _GEN_7092 : _GEN_7860; // @[executor.scala 466:52]
  wire [7:0] _GEN_8119 = opcode_7 == 4'hf ? _GEN_7093 : _GEN_7861; // @[executor.scala 466:52]
  wire [7:0] _GEN_8120 = opcode_7 == 4'hf ? _GEN_7094 : _GEN_7862; // @[executor.scala 466:52]
  wire [7:0] _GEN_8121 = opcode_7 == 4'hf ? _GEN_7095 : _GEN_7863; // @[executor.scala 466:52]
  wire [7:0] _GEN_8122 = opcode_7 == 4'hf ? _GEN_7096 : _GEN_7864; // @[executor.scala 466:52]
  wire [7:0] _GEN_8123 = opcode_7 == 4'hf ? _GEN_7097 : _GEN_7865; // @[executor.scala 466:52]
  wire [7:0] _GEN_8124 = opcode_7 == 4'hf ? _GEN_7098 : _GEN_7866; // @[executor.scala 466:52]
  wire [7:0] _GEN_8125 = opcode_7 == 4'hf ? _GEN_7099 : _GEN_7867; // @[executor.scala 466:52]
  wire [7:0] _GEN_8126 = opcode_7 == 4'hf ? _GEN_7100 : _GEN_7868; // @[executor.scala 466:52]
  wire [7:0] _GEN_8127 = opcode_7 == 4'hf ? _GEN_7101 : _GEN_7869; // @[executor.scala 466:52]
  wire [7:0] _GEN_8128 = opcode_7 == 4'hf ? _GEN_7102 : _GEN_7870; // @[executor.scala 466:52]
  wire [7:0] _GEN_8129 = opcode_7 == 4'hf ? _GEN_7103 : _GEN_7871; // @[executor.scala 466:52]
  wire [7:0] _GEN_8130 = opcode_7 == 4'hf ? _GEN_7104 : _GEN_7872; // @[executor.scala 466:52]
  wire [7:0] _GEN_8131 = opcode_7 == 4'hf ? _GEN_7105 : _GEN_7873; // @[executor.scala 466:52]
  wire [7:0] _GEN_8132 = opcode_7 == 4'hf ? _GEN_7106 : _GEN_7874; // @[executor.scala 466:52]
  wire [7:0] _GEN_8133 = opcode_7 == 4'hf ? _GEN_7107 : _GEN_7875; // @[executor.scala 466:52]
  wire [7:0] _GEN_8134 = opcode_7 == 4'hf ? _GEN_7108 : _GEN_7876; // @[executor.scala 466:52]
  wire [7:0] _GEN_8135 = opcode_7 == 4'hf ? _GEN_7109 : _GEN_7877; // @[executor.scala 466:52]
  wire [7:0] _GEN_8136 = opcode_7 == 4'hf ? _GEN_7110 : _GEN_7878; // @[executor.scala 466:52]
  wire [7:0] _GEN_8137 = opcode_7 == 4'hf ? _GEN_7111 : _GEN_7879; // @[executor.scala 466:52]
  wire [7:0] _GEN_8138 = opcode_7 == 4'hf ? _GEN_7112 : _GEN_7880; // @[executor.scala 466:52]
  wire [7:0] _GEN_8139 = opcode_7 == 4'hf ? _GEN_7113 : _GEN_7881; // @[executor.scala 466:52]
  wire [7:0] _GEN_8140 = opcode_7 == 4'hf ? _GEN_7114 : _GEN_7882; // @[executor.scala 466:52]
  wire [7:0] _GEN_8141 = opcode_7 == 4'hf ? _GEN_7115 : _GEN_7883; // @[executor.scala 466:52]
  wire [7:0] _GEN_8142 = opcode_7 == 4'hf ? _GEN_7116 : _GEN_7884; // @[executor.scala 466:52]
  wire [7:0] _GEN_8143 = opcode_7 == 4'hf ? _GEN_7117 : _GEN_7885; // @[executor.scala 466:52]
  wire [7:0] _GEN_8144 = opcode_7 == 4'hf ? _GEN_7118 : _GEN_7886; // @[executor.scala 466:52]
  wire [7:0] _GEN_8145 = opcode_7 == 4'hf ? _GEN_7119 : _GEN_7887; // @[executor.scala 466:52]
  wire [7:0] _GEN_8146 = opcode_7 == 4'hf ? _GEN_7120 : _GEN_7888; // @[executor.scala 466:52]
  wire [7:0] _GEN_8147 = opcode_7 == 4'hf ? _GEN_7121 : _GEN_7889; // @[executor.scala 466:52]
  wire [7:0] _GEN_8148 = opcode_7 == 4'hf ? _GEN_7122 : _GEN_7890; // @[executor.scala 466:52]
  wire [7:0] _GEN_8149 = opcode_7 == 4'hf ? _GEN_7123 : _GEN_7891; // @[executor.scala 466:52]
  wire [7:0] _GEN_8150 = opcode_7 == 4'hf ? _GEN_7124 : _GEN_7892; // @[executor.scala 466:52]
  wire [7:0] _GEN_8151 = opcode_7 == 4'hf ? _GEN_7125 : _GEN_7893; // @[executor.scala 466:52]
  wire [7:0] _GEN_8152 = opcode_7 == 4'hf ? _GEN_7126 : _GEN_7894; // @[executor.scala 466:52]
  wire [7:0] _GEN_8153 = opcode_7 == 4'hf ? _GEN_7127 : _GEN_7895; // @[executor.scala 466:52]
  wire [7:0] _GEN_8154 = opcode_7 == 4'hf ? _GEN_7128 : _GEN_7896; // @[executor.scala 466:52]
  wire [7:0] _GEN_8155 = opcode_7 == 4'hf ? _GEN_7129 : _GEN_7897; // @[executor.scala 466:52]
  wire [7:0] _GEN_8156 = opcode_7 == 4'hf ? _GEN_7130 : _GEN_7898; // @[executor.scala 466:52]
  wire [7:0] _GEN_8157 = opcode_7 == 4'hf ? _GEN_7131 : _GEN_7899; // @[executor.scala 466:52]
  wire [7:0] _GEN_8158 = opcode_7 == 4'hf ? _GEN_7132 : _GEN_7900; // @[executor.scala 466:52]
  wire [7:0] _GEN_8159 = opcode_7 == 4'hf ? _GEN_7133 : _GEN_7901; // @[executor.scala 466:52]
  wire [7:0] _GEN_8160 = opcode_7 == 4'hf ? _GEN_7134 : _GEN_7902; // @[executor.scala 466:52]
  wire [7:0] _GEN_8161 = opcode_7 == 4'hf ? _GEN_7135 : _GEN_7903; // @[executor.scala 466:52]
  wire [7:0] _GEN_8162 = opcode_7 == 4'hf ? _GEN_7136 : _GEN_7904; // @[executor.scala 466:52]
  wire [7:0] _GEN_8163 = opcode_7 == 4'hf ? _GEN_7137 : _GEN_7905; // @[executor.scala 466:52]
  wire [7:0] _GEN_8164 = opcode_7 == 4'hf ? _GEN_7138 : _GEN_7906; // @[executor.scala 466:52]
  wire [7:0] _GEN_8165 = opcode_7 == 4'hf ? _GEN_7139 : _GEN_7907; // @[executor.scala 466:52]
  wire [7:0] _GEN_8166 = opcode_7 == 4'hf ? _GEN_7140 : _GEN_7908; // @[executor.scala 466:52]
  wire [7:0] _GEN_8167 = opcode_7 == 4'hf ? _GEN_7141 : _GEN_7909; // @[executor.scala 466:52]
  wire [7:0] _GEN_8168 = opcode_7 == 4'hf ? _GEN_7142 : _GEN_7910; // @[executor.scala 466:52]
  wire [7:0] _GEN_8169 = opcode_7 == 4'hf ? _GEN_7143 : _GEN_7911; // @[executor.scala 466:52]
  wire [7:0] _GEN_8170 = opcode_7 == 4'hf ? _GEN_7144 : _GEN_7912; // @[executor.scala 466:52]
  wire [7:0] _GEN_8171 = opcode_7 == 4'hf ? _GEN_7145 : _GEN_7913; // @[executor.scala 466:52]
  wire [7:0] _GEN_8172 = opcode_7 == 4'hf ? _GEN_7146 : _GEN_7914; // @[executor.scala 466:52]
  wire [7:0] _GEN_8173 = opcode_7 == 4'hf ? _GEN_7147 : _GEN_7915; // @[executor.scala 466:52]
  wire [7:0] _GEN_8174 = opcode_7 == 4'hf ? _GEN_7148 : _GEN_7916; // @[executor.scala 466:52]
  wire [7:0] _GEN_8175 = opcode_7 == 4'hf ? _GEN_7149 : _GEN_7917; // @[executor.scala 466:52]
  wire [7:0] _GEN_8176 = opcode_7 == 4'hf ? _GEN_7150 : _GEN_7918; // @[executor.scala 466:52]
  wire [7:0] _GEN_8177 = opcode_7 == 4'hf ? _GEN_7151 : _GEN_7919; // @[executor.scala 466:52]
  wire [7:0] _GEN_8178 = opcode_7 == 4'hf ? _GEN_7152 : _GEN_7920; // @[executor.scala 466:52]
  wire [7:0] _GEN_8179 = opcode_7 == 4'hf ? _GEN_7153 : _GEN_7921; // @[executor.scala 466:52]
  wire [7:0] _GEN_8180 = opcode_7 == 4'hf ? _GEN_7154 : _GEN_7922; // @[executor.scala 466:52]
  wire [7:0] _GEN_8181 = opcode_7 == 4'hf ? _GEN_7155 : _GEN_7923; // @[executor.scala 466:52]
  wire [7:0] _GEN_8182 = opcode_7 == 4'hf ? _GEN_7156 : _GEN_7924; // @[executor.scala 466:52]
  wire [7:0] _GEN_8183 = opcode_7 == 4'hf ? _GEN_7157 : _GEN_7925; // @[executor.scala 466:52]
  wire [7:0] _GEN_8184 = opcode_7 == 4'hf ? _GEN_7158 : _GEN_7926; // @[executor.scala 466:52]
  wire [7:0] _GEN_8185 = opcode_7 == 4'hf ? _GEN_7159 : _GEN_7927; // @[executor.scala 466:52]
  wire [7:0] _GEN_8186 = opcode_7 == 4'hf ? _GEN_7160 : _GEN_7928; // @[executor.scala 466:52]
  wire [7:0] _GEN_8187 = opcode_7 == 4'hf ? _GEN_7161 : _GEN_7929; // @[executor.scala 466:52]
  wire [7:0] _GEN_8188 = opcode_7 == 4'hf ? _GEN_7162 : _GEN_7930; // @[executor.scala 466:52]
  wire [7:0] _GEN_8189 = opcode_7 == 4'hf ? _GEN_7163 : _GEN_7931; // @[executor.scala 466:52]
  wire [7:0] _GEN_8190 = opcode_7 == 4'hf ? _GEN_7164 : _GEN_7932; // @[executor.scala 466:52]
  wire [7:0] _GEN_8191 = opcode_7 == 4'hf ? _GEN_7165 : _GEN_7933; // @[executor.scala 466:52]
  wire [7:0] _GEN_8192 = opcode_7 == 4'hf ? _GEN_7166 : _GEN_7934; // @[executor.scala 466:52]
  wire [7:0] _GEN_8193 = opcode_7 == 4'hf ? _GEN_7167 : _GEN_7935; // @[executor.scala 466:52]
  wire [7:0] _GEN_8194 = opcode_7 == 4'hf ? _GEN_7168 : _GEN_7936; // @[executor.scala 466:52]
  wire [7:0] _GEN_8195 = opcode_7 == 4'hf ? _GEN_7169 : _GEN_7937; // @[executor.scala 466:52]
  wire [7:0] _GEN_8196 = opcode_7 == 4'hf ? _GEN_7170 : _GEN_7938; // @[executor.scala 466:52]
  wire [7:0] _GEN_8197 = opcode_7 == 4'hf ? _GEN_7171 : _GEN_7939; // @[executor.scala 466:52]
  wire [7:0] _GEN_8198 = opcode_7 == 4'hf ? _GEN_7172 : _GEN_7940; // @[executor.scala 466:52]
  wire [7:0] _GEN_8199 = opcode_7 == 4'hf ? _GEN_7173 : _GEN_7941; // @[executor.scala 466:52]
  wire [7:0] _GEN_8200 = opcode_7 == 4'hf ? _GEN_7174 : _GEN_7942; // @[executor.scala 466:52]
  wire [7:0] _GEN_8201 = opcode_7 == 4'hf ? _GEN_7175 : _GEN_7943; // @[executor.scala 466:52]
  wire [7:0] _GEN_8202 = opcode_7 == 4'hf ? _GEN_7176 : _GEN_7944; // @[executor.scala 466:52]
  wire [7:0] _GEN_8203 = opcode_7 == 4'hf ? _GEN_7177 : _GEN_7945; // @[executor.scala 466:52]
  wire [7:0] _GEN_8204 = opcode_7 == 4'hf ? _GEN_7178 : _GEN_7946; // @[executor.scala 466:52]
  wire [7:0] _GEN_8205 = opcode_7 == 4'hf ? _GEN_7179 : _GEN_7947; // @[executor.scala 466:52]
  wire [7:0] _GEN_8206 = opcode_7 == 4'hf ? _GEN_7180 : _GEN_7948; // @[executor.scala 466:52]
  wire [7:0] _GEN_8207 = opcode_7 == 4'hf ? _GEN_7181 : _GEN_7949; // @[executor.scala 466:52]
  assign io_pipe_phv_out_data_0 = phv_is_valid_processor ? _GEN_7955 : phv_data_0; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_1 = phv_is_valid_processor ? _GEN_7954 : phv_data_1; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_2 = phv_is_valid_processor ? _GEN_7953 : phv_data_2; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_3 = phv_is_valid_processor ? _GEN_7952 : phv_data_3; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_4 = phv_is_valid_processor ? _GEN_7959 : phv_data_4; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_5 = phv_is_valid_processor ? _GEN_7958 : phv_data_5; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_6 = phv_is_valid_processor ? _GEN_7957 : phv_data_6; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_7 = phv_is_valid_processor ? _GEN_7956 : phv_data_7; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_8 = phv_is_valid_processor ? _GEN_7963 : phv_data_8; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_9 = phv_is_valid_processor ? _GEN_7962 : phv_data_9; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_10 = phv_is_valid_processor ? _GEN_7961 : phv_data_10; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_11 = phv_is_valid_processor ? _GEN_7960 : phv_data_11; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_12 = phv_is_valid_processor ? _GEN_7967 : phv_data_12; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_13 = phv_is_valid_processor ? _GEN_7966 : phv_data_13; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_14 = phv_is_valid_processor ? _GEN_7965 : phv_data_14; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_15 = phv_is_valid_processor ? _GEN_7964 : phv_data_15; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_16 = phv_is_valid_processor ? _GEN_7971 : phv_data_16; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_17 = phv_is_valid_processor ? _GEN_7970 : phv_data_17; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_18 = phv_is_valid_processor ? _GEN_7969 : phv_data_18; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_19 = phv_is_valid_processor ? _GEN_7968 : phv_data_19; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_20 = phv_is_valid_processor ? _GEN_7975 : phv_data_20; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_21 = phv_is_valid_processor ? _GEN_7974 : phv_data_21; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_22 = phv_is_valid_processor ? _GEN_7973 : phv_data_22; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_23 = phv_is_valid_processor ? _GEN_7972 : phv_data_23; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_24 = phv_is_valid_processor ? _GEN_7979 : phv_data_24; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_25 = phv_is_valid_processor ? _GEN_7978 : phv_data_25; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_26 = phv_is_valid_processor ? _GEN_7977 : phv_data_26; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_27 = phv_is_valid_processor ? _GEN_7976 : phv_data_27; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_28 = phv_is_valid_processor ? _GEN_7983 : phv_data_28; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_29 = phv_is_valid_processor ? _GEN_7982 : phv_data_29; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_30 = phv_is_valid_processor ? _GEN_7981 : phv_data_30; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_31 = phv_is_valid_processor ? _GEN_7980 : phv_data_31; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_32 = phv_is_valid_processor ? _GEN_7987 : phv_data_32; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_33 = phv_is_valid_processor ? _GEN_7986 : phv_data_33; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_34 = phv_is_valid_processor ? _GEN_7985 : phv_data_34; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_35 = phv_is_valid_processor ? _GEN_7984 : phv_data_35; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_36 = phv_is_valid_processor ? _GEN_7991 : phv_data_36; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_37 = phv_is_valid_processor ? _GEN_7990 : phv_data_37; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_38 = phv_is_valid_processor ? _GEN_7989 : phv_data_38; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_39 = phv_is_valid_processor ? _GEN_7988 : phv_data_39; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_40 = phv_is_valid_processor ? _GEN_7995 : phv_data_40; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_41 = phv_is_valid_processor ? _GEN_7994 : phv_data_41; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_42 = phv_is_valid_processor ? _GEN_7993 : phv_data_42; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_43 = phv_is_valid_processor ? _GEN_7992 : phv_data_43; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_44 = phv_is_valid_processor ? _GEN_7999 : phv_data_44; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_45 = phv_is_valid_processor ? _GEN_7998 : phv_data_45; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_46 = phv_is_valid_processor ? _GEN_7997 : phv_data_46; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_47 = phv_is_valid_processor ? _GEN_7996 : phv_data_47; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_48 = phv_is_valid_processor ? _GEN_8003 : phv_data_48; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_49 = phv_is_valid_processor ? _GEN_8002 : phv_data_49; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_50 = phv_is_valid_processor ? _GEN_8001 : phv_data_50; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_51 = phv_is_valid_processor ? _GEN_8000 : phv_data_51; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_52 = phv_is_valid_processor ? _GEN_8007 : phv_data_52; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_53 = phv_is_valid_processor ? _GEN_8006 : phv_data_53; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_54 = phv_is_valid_processor ? _GEN_8005 : phv_data_54; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_55 = phv_is_valid_processor ? _GEN_8004 : phv_data_55; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_56 = phv_is_valid_processor ? _GEN_8011 : phv_data_56; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_57 = phv_is_valid_processor ? _GEN_8010 : phv_data_57; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_58 = phv_is_valid_processor ? _GEN_8009 : phv_data_58; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_59 = phv_is_valid_processor ? _GEN_8008 : phv_data_59; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_60 = phv_is_valid_processor ? _GEN_8015 : phv_data_60; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_61 = phv_is_valid_processor ? _GEN_8014 : phv_data_61; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_62 = phv_is_valid_processor ? _GEN_8013 : phv_data_62; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_63 = phv_is_valid_processor ? _GEN_8012 : phv_data_63; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_64 = phv_is_valid_processor ? _GEN_8019 : phv_data_64; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_65 = phv_is_valid_processor ? _GEN_8018 : phv_data_65; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_66 = phv_is_valid_processor ? _GEN_8017 : phv_data_66; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_67 = phv_is_valid_processor ? _GEN_8016 : phv_data_67; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_68 = phv_is_valid_processor ? _GEN_8023 : phv_data_68; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_69 = phv_is_valid_processor ? _GEN_8022 : phv_data_69; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_70 = phv_is_valid_processor ? _GEN_8021 : phv_data_70; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_71 = phv_is_valid_processor ? _GEN_8020 : phv_data_71; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_72 = phv_is_valid_processor ? _GEN_8027 : phv_data_72; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_73 = phv_is_valid_processor ? _GEN_8026 : phv_data_73; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_74 = phv_is_valid_processor ? _GEN_8025 : phv_data_74; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_75 = phv_is_valid_processor ? _GEN_8024 : phv_data_75; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_76 = phv_is_valid_processor ? _GEN_8031 : phv_data_76; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_77 = phv_is_valid_processor ? _GEN_8030 : phv_data_77; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_78 = phv_is_valid_processor ? _GEN_8029 : phv_data_78; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_79 = phv_is_valid_processor ? _GEN_8028 : phv_data_79; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_80 = phv_is_valid_processor ? _GEN_8035 : phv_data_80; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_81 = phv_is_valid_processor ? _GEN_8034 : phv_data_81; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_82 = phv_is_valid_processor ? _GEN_8033 : phv_data_82; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_83 = phv_is_valid_processor ? _GEN_8032 : phv_data_83; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_84 = phv_is_valid_processor ? _GEN_8039 : phv_data_84; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_85 = phv_is_valid_processor ? _GEN_8038 : phv_data_85; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_86 = phv_is_valid_processor ? _GEN_8037 : phv_data_86; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_87 = phv_is_valid_processor ? _GEN_8036 : phv_data_87; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_88 = phv_is_valid_processor ? _GEN_8043 : phv_data_88; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_89 = phv_is_valid_processor ? _GEN_8042 : phv_data_89; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_90 = phv_is_valid_processor ? _GEN_8041 : phv_data_90; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_91 = phv_is_valid_processor ? _GEN_8040 : phv_data_91; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_92 = phv_is_valid_processor ? _GEN_8047 : phv_data_92; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_93 = phv_is_valid_processor ? _GEN_8046 : phv_data_93; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_94 = phv_is_valid_processor ? _GEN_8045 : phv_data_94; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_95 = phv_is_valid_processor ? _GEN_8044 : phv_data_95; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_96 = phv_is_valid_processor ? _GEN_8051 : phv_data_96; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_97 = phv_is_valid_processor ? _GEN_8050 : phv_data_97; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_98 = phv_is_valid_processor ? _GEN_8049 : phv_data_98; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_99 = phv_is_valid_processor ? _GEN_8048 : phv_data_99; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_100 = phv_is_valid_processor ? _GEN_8055 : phv_data_100; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_101 = phv_is_valid_processor ? _GEN_8054 : phv_data_101; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_102 = phv_is_valid_processor ? _GEN_8053 : phv_data_102; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_103 = phv_is_valid_processor ? _GEN_8052 : phv_data_103; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_104 = phv_is_valid_processor ? _GEN_8059 : phv_data_104; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_105 = phv_is_valid_processor ? _GEN_8058 : phv_data_105; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_106 = phv_is_valid_processor ? _GEN_8057 : phv_data_106; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_107 = phv_is_valid_processor ? _GEN_8056 : phv_data_107; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_108 = phv_is_valid_processor ? _GEN_8063 : phv_data_108; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_109 = phv_is_valid_processor ? _GEN_8062 : phv_data_109; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_110 = phv_is_valid_processor ? _GEN_8061 : phv_data_110; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_111 = phv_is_valid_processor ? _GEN_8060 : phv_data_111; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_112 = phv_is_valid_processor ? _GEN_8067 : phv_data_112; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_113 = phv_is_valid_processor ? _GEN_8066 : phv_data_113; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_114 = phv_is_valid_processor ? _GEN_8065 : phv_data_114; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_115 = phv_is_valid_processor ? _GEN_8064 : phv_data_115; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_116 = phv_is_valid_processor ? _GEN_8071 : phv_data_116; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_117 = phv_is_valid_processor ? _GEN_8070 : phv_data_117; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_118 = phv_is_valid_processor ? _GEN_8069 : phv_data_118; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_119 = phv_is_valid_processor ? _GEN_8068 : phv_data_119; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_120 = phv_is_valid_processor ? _GEN_8075 : phv_data_120; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_121 = phv_is_valid_processor ? _GEN_8074 : phv_data_121; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_122 = phv_is_valid_processor ? _GEN_8073 : phv_data_122; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_123 = phv_is_valid_processor ? _GEN_8072 : phv_data_123; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_124 = phv_is_valid_processor ? _GEN_8079 : phv_data_124; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_125 = phv_is_valid_processor ? _GEN_8078 : phv_data_125; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_126 = phv_is_valid_processor ? _GEN_8077 : phv_data_126; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_127 = phv_is_valid_processor ? _GEN_8076 : phv_data_127; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_128 = phv_is_valid_processor ? _GEN_8083 : phv_data_128; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_129 = phv_is_valid_processor ? _GEN_8082 : phv_data_129; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_130 = phv_is_valid_processor ? _GEN_8081 : phv_data_130; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_131 = phv_is_valid_processor ? _GEN_8080 : phv_data_131; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_132 = phv_is_valid_processor ? _GEN_8087 : phv_data_132; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_133 = phv_is_valid_processor ? _GEN_8086 : phv_data_133; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_134 = phv_is_valid_processor ? _GEN_8085 : phv_data_134; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_135 = phv_is_valid_processor ? _GEN_8084 : phv_data_135; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_136 = phv_is_valid_processor ? _GEN_8091 : phv_data_136; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_137 = phv_is_valid_processor ? _GEN_8090 : phv_data_137; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_138 = phv_is_valid_processor ? _GEN_8089 : phv_data_138; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_139 = phv_is_valid_processor ? _GEN_8088 : phv_data_139; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_140 = phv_is_valid_processor ? _GEN_8095 : phv_data_140; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_141 = phv_is_valid_processor ? _GEN_8094 : phv_data_141; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_142 = phv_is_valid_processor ? _GEN_8093 : phv_data_142; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_143 = phv_is_valid_processor ? _GEN_8092 : phv_data_143; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_144 = phv_is_valid_processor ? _GEN_8099 : phv_data_144; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_145 = phv_is_valid_processor ? _GEN_8098 : phv_data_145; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_146 = phv_is_valid_processor ? _GEN_8097 : phv_data_146; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_147 = phv_is_valid_processor ? _GEN_8096 : phv_data_147; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_148 = phv_is_valid_processor ? _GEN_8103 : phv_data_148; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_149 = phv_is_valid_processor ? _GEN_8102 : phv_data_149; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_150 = phv_is_valid_processor ? _GEN_8101 : phv_data_150; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_151 = phv_is_valid_processor ? _GEN_8100 : phv_data_151; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_152 = phv_is_valid_processor ? _GEN_8107 : phv_data_152; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_153 = phv_is_valid_processor ? _GEN_8106 : phv_data_153; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_154 = phv_is_valid_processor ? _GEN_8105 : phv_data_154; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_155 = phv_is_valid_processor ? _GEN_8104 : phv_data_155; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_156 = phv_is_valid_processor ? _GEN_8111 : phv_data_156; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_157 = phv_is_valid_processor ? _GEN_8110 : phv_data_157; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_158 = phv_is_valid_processor ? _GEN_8109 : phv_data_158; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_159 = phv_is_valid_processor ? _GEN_8108 : phv_data_159; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_160 = phv_is_valid_processor ? _GEN_8115 : phv_data_160; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_161 = phv_is_valid_processor ? _GEN_8114 : phv_data_161; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_162 = phv_is_valid_processor ? _GEN_8113 : phv_data_162; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_163 = phv_is_valid_processor ? _GEN_8112 : phv_data_163; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_164 = phv_is_valid_processor ? _GEN_8119 : phv_data_164; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_165 = phv_is_valid_processor ? _GEN_8118 : phv_data_165; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_166 = phv_is_valid_processor ? _GEN_8117 : phv_data_166; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_167 = phv_is_valid_processor ? _GEN_8116 : phv_data_167; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_168 = phv_is_valid_processor ? _GEN_8123 : phv_data_168; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_169 = phv_is_valid_processor ? _GEN_8122 : phv_data_169; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_170 = phv_is_valid_processor ? _GEN_8121 : phv_data_170; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_171 = phv_is_valid_processor ? _GEN_8120 : phv_data_171; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_172 = phv_is_valid_processor ? _GEN_8127 : phv_data_172; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_173 = phv_is_valid_processor ? _GEN_8126 : phv_data_173; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_174 = phv_is_valid_processor ? _GEN_8125 : phv_data_174; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_175 = phv_is_valid_processor ? _GEN_8124 : phv_data_175; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_176 = phv_is_valid_processor ? _GEN_8131 : phv_data_176; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_177 = phv_is_valid_processor ? _GEN_8130 : phv_data_177; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_178 = phv_is_valid_processor ? _GEN_8129 : phv_data_178; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_179 = phv_is_valid_processor ? _GEN_8128 : phv_data_179; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_180 = phv_is_valid_processor ? _GEN_8135 : phv_data_180; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_181 = phv_is_valid_processor ? _GEN_8134 : phv_data_181; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_182 = phv_is_valid_processor ? _GEN_8133 : phv_data_182; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_183 = phv_is_valid_processor ? _GEN_8132 : phv_data_183; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_184 = phv_is_valid_processor ? _GEN_8139 : phv_data_184; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_185 = phv_is_valid_processor ? _GEN_8138 : phv_data_185; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_186 = phv_is_valid_processor ? _GEN_8137 : phv_data_186; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_187 = phv_is_valid_processor ? _GEN_8136 : phv_data_187; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_188 = phv_is_valid_processor ? _GEN_8143 : phv_data_188; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_189 = phv_is_valid_processor ? _GEN_8142 : phv_data_189; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_190 = phv_is_valid_processor ? _GEN_8141 : phv_data_190; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_191 = phv_is_valid_processor ? _GEN_8140 : phv_data_191; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_192 = phv_is_valid_processor ? _GEN_8147 : phv_data_192; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_193 = phv_is_valid_processor ? _GEN_8146 : phv_data_193; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_194 = phv_is_valid_processor ? _GEN_8145 : phv_data_194; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_195 = phv_is_valid_processor ? _GEN_8144 : phv_data_195; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_196 = phv_is_valid_processor ? _GEN_8151 : phv_data_196; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_197 = phv_is_valid_processor ? _GEN_8150 : phv_data_197; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_198 = phv_is_valid_processor ? _GEN_8149 : phv_data_198; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_199 = phv_is_valid_processor ? _GEN_8148 : phv_data_199; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_200 = phv_is_valid_processor ? _GEN_8155 : phv_data_200; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_201 = phv_is_valid_processor ? _GEN_8154 : phv_data_201; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_202 = phv_is_valid_processor ? _GEN_8153 : phv_data_202; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_203 = phv_is_valid_processor ? _GEN_8152 : phv_data_203; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_204 = phv_is_valid_processor ? _GEN_8159 : phv_data_204; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_205 = phv_is_valid_processor ? _GEN_8158 : phv_data_205; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_206 = phv_is_valid_processor ? _GEN_8157 : phv_data_206; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_207 = phv_is_valid_processor ? _GEN_8156 : phv_data_207; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_208 = phv_is_valid_processor ? _GEN_8163 : phv_data_208; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_209 = phv_is_valid_processor ? _GEN_8162 : phv_data_209; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_210 = phv_is_valid_processor ? _GEN_8161 : phv_data_210; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_211 = phv_is_valid_processor ? _GEN_8160 : phv_data_211; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_212 = phv_is_valid_processor ? _GEN_8167 : phv_data_212; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_213 = phv_is_valid_processor ? _GEN_8166 : phv_data_213; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_214 = phv_is_valid_processor ? _GEN_8165 : phv_data_214; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_215 = phv_is_valid_processor ? _GEN_8164 : phv_data_215; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_216 = phv_is_valid_processor ? _GEN_8171 : phv_data_216; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_217 = phv_is_valid_processor ? _GEN_8170 : phv_data_217; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_218 = phv_is_valid_processor ? _GEN_8169 : phv_data_218; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_219 = phv_is_valid_processor ? _GEN_8168 : phv_data_219; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_220 = phv_is_valid_processor ? _GEN_8175 : phv_data_220; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_221 = phv_is_valid_processor ? _GEN_8174 : phv_data_221; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_222 = phv_is_valid_processor ? _GEN_8173 : phv_data_222; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_223 = phv_is_valid_processor ? _GEN_8172 : phv_data_223; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_224 = phv_is_valid_processor ? _GEN_8179 : phv_data_224; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_225 = phv_is_valid_processor ? _GEN_8178 : phv_data_225; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_226 = phv_is_valid_processor ? _GEN_8177 : phv_data_226; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_227 = phv_is_valid_processor ? _GEN_8176 : phv_data_227; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_228 = phv_is_valid_processor ? _GEN_8183 : phv_data_228; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_229 = phv_is_valid_processor ? _GEN_8182 : phv_data_229; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_230 = phv_is_valid_processor ? _GEN_8181 : phv_data_230; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_231 = phv_is_valid_processor ? _GEN_8180 : phv_data_231; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_232 = phv_is_valid_processor ? _GEN_8187 : phv_data_232; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_233 = phv_is_valid_processor ? _GEN_8186 : phv_data_233; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_234 = phv_is_valid_processor ? _GEN_8185 : phv_data_234; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_235 = phv_is_valid_processor ? _GEN_8184 : phv_data_235; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_236 = phv_is_valid_processor ? _GEN_8191 : phv_data_236; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_237 = phv_is_valid_processor ? _GEN_8190 : phv_data_237; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_238 = phv_is_valid_processor ? _GEN_8189 : phv_data_238; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_239 = phv_is_valid_processor ? _GEN_8188 : phv_data_239; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_240 = phv_is_valid_processor ? _GEN_8195 : phv_data_240; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_241 = phv_is_valid_processor ? _GEN_8194 : phv_data_241; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_242 = phv_is_valid_processor ? _GEN_8193 : phv_data_242; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_243 = phv_is_valid_processor ? _GEN_8192 : phv_data_243; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_244 = phv_is_valid_processor ? _GEN_8199 : phv_data_244; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_245 = phv_is_valid_processor ? _GEN_8198 : phv_data_245; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_246 = phv_is_valid_processor ? _GEN_8197 : phv_data_246; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_247 = phv_is_valid_processor ? _GEN_8196 : phv_data_247; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_248 = phv_is_valid_processor ? _GEN_8203 : phv_data_248; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_249 = phv_is_valid_processor ? _GEN_8202 : phv_data_249; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_250 = phv_is_valid_processor ? _GEN_8201 : phv_data_250; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_251 = phv_is_valid_processor ? _GEN_8200 : phv_data_251; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_252 = phv_is_valid_processor ? _GEN_8207 : phv_data_252; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_253 = phv_is_valid_processor ? _GEN_8206 : phv_data_253; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_254 = phv_is_valid_processor ? _GEN_8205 : phv_data_254; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_255 = phv_is_valid_processor ? _GEN_8204 : phv_data_255; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 450:25]
  assign io_pipe_phv_out_next_processor_id = phv_is_valid_processor ? _GEN_7950 : phv_next_processor_id; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_next_config_id = phv_is_valid_processor ? _GEN_7951 : phv_next_config_id; // @[executor.scala 461:39 executor.scala 450:25]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 449:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 449:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 449:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 449:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 449:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 449:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 449:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 449:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 449:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 449:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 449:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 449:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 449:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 449:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 449:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 449:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 449:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 449:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 449:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 449:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 449:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 449:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 449:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 449:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 449:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 449:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 449:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 449:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 449:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 449:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 449:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 449:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 449:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 449:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 449:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 449:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 449:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 449:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 449:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 449:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 449:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 449:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 449:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 449:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 449:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 449:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 449:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 449:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 449:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 449:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 449:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 449:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 449:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 449:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 449:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 449:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 449:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 449:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 449:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 449:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 449:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 449:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 449:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 449:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 449:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 449:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 449:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 449:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 449:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 449:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 449:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 449:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 449:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 449:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 449:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 449:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 449:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 449:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 449:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 449:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 449:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 449:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 449:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 449:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 449:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 449:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 449:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 449:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 449:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 449:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 449:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 449:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 449:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 449:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 449:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 449:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor.scala 449:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor.scala 449:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor.scala 449:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor.scala 449:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor.scala 449:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor.scala 449:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor.scala 449:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor.scala 449:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor.scala 449:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor.scala 449:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor.scala 449:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor.scala 449:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor.scala 449:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor.scala 449:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor.scala 449:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor.scala 449:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor.scala 449:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor.scala 449:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor.scala 449:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor.scala 449:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor.scala 449:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor.scala 449:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor.scala 449:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor.scala 449:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor.scala 449:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor.scala 449:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor.scala 449:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor.scala 449:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor.scala 449:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor.scala 449:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor.scala 449:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor.scala 449:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor.scala 449:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor.scala 449:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor.scala 449:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor.scala 449:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor.scala 449:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor.scala 449:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor.scala 449:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor.scala 449:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor.scala 449:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor.scala 449:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor.scala 449:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor.scala 449:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor.scala 449:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor.scala 449:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor.scala 449:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor.scala 449:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor.scala 449:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor.scala 449:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor.scala 449:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor.scala 449:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor.scala 449:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor.scala 449:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor.scala 449:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor.scala 449:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor.scala 449:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor.scala 449:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor.scala 449:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor.scala 449:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor.scala 449:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor.scala 449:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor.scala 449:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor.scala 449:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor.scala 449:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor.scala 449:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor.scala 449:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor.scala 449:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor.scala 449:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor.scala 449:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor.scala 449:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor.scala 449:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor.scala 449:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor.scala 449:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor.scala 449:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor.scala 449:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor.scala 449:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor.scala 449:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor.scala 449:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor.scala 449:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor.scala 449:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor.scala 449:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor.scala 449:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor.scala 449:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor.scala 449:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor.scala 449:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor.scala 449:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor.scala 449:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor.scala 449:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor.scala 449:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor.scala 449:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor.scala 449:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor.scala 449:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor.scala 449:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor.scala 449:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor.scala 449:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor.scala 449:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor.scala 449:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor.scala 449:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor.scala 449:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor.scala 449:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor.scala 449:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor.scala 449:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor.scala 449:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor.scala 449:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor.scala 449:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor.scala 449:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor.scala 449:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor.scala 449:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor.scala 449:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor.scala 449:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor.scala 449:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor.scala 449:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor.scala 449:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor.scala 449:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor.scala 449:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor.scala 449:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor.scala 449:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor.scala 449:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor.scala 449:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor.scala 449:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor.scala 449:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor.scala 449:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor.scala 449:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor.scala 449:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor.scala 449:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor.scala 449:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor.scala 449:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor.scala 449:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor.scala 449:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor.scala 449:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor.scala 449:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor.scala 449:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor.scala 449:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor.scala 449:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor.scala 449:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor.scala 449:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor.scala 449:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor.scala 449:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor.scala 449:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor.scala 449:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor.scala 449:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor.scala 449:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor.scala 449:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor.scala 449:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor.scala 449:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor.scala 449:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor.scala 449:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor.scala 449:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor.scala 449:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor.scala 449:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor.scala 449:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor.scala 449:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor.scala 449:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor.scala 449:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor.scala 449:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor.scala 449:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor.scala 449:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor.scala 449:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor.scala 449:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 449:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 449:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 449:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 449:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 449:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 449:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 449:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 449:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 449:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 449:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 449:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 449:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 449:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 449:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 449:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 449:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 449:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 449:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 449:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 449:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor.scala 449:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 449:13]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 453:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 453:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 453:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 453:14]
    vliw_4 <= io_vliw_in_4; // @[executor.scala 453:14]
    vliw_5 <= io_vliw_in_5; // @[executor.scala 453:14]
    vliw_6 <= io_vliw_in_6; // @[executor.scala 453:14]
    vliw_7 <= io_vliw_in_7; // @[executor.scala 453:14]
    field_0 <= io_field_in_0; // @[executor.scala 455:15]
    field_1 <= io_field_in_1; // @[executor.scala 455:15]
    field_2 <= io_field_in_2; // @[executor.scala 455:15]
    field_3 <= io_field_in_3; // @[executor.scala 455:15]
    field_4 <= io_field_in_4; // @[executor.scala 455:15]
    field_5 <= io_field_in_5; // @[executor.scala 455:15]
    field_6 <= io_field_in_6; // @[executor.scala 455:15]
    field_7 <= io_field_in_7; // @[executor.scala 455:15]
    mask_0 <= io_mask_in_0; // @[executor.scala 457:14]
    mask_1 <= io_mask_in_1; // @[executor.scala 457:14]
    mask_2 <= io_mask_in_2; // @[executor.scala 457:14]
    mask_3 <= io_mask_in_3; // @[executor.scala 457:14]
    mask_4 <= io_mask_in_4; // @[executor.scala 457:14]
    mask_5 <= io_mask_in_5; // @[executor.scala 457:14]
    mask_6 <= io_mask_in_6; // @[executor.scala 457:14]
    mask_7 <= io_mask_in_7; // @[executor.scala 457:14]
    dst_offset_0 <= io_dst_offset_in_0; // @[executor.scala 459:20]
    dst_offset_1 <= io_dst_offset_in_1; // @[executor.scala 459:20]
    dst_offset_2 <= io_dst_offset_in_2; // @[executor.scala 459:20]
    dst_offset_3 <= io_dst_offset_in_3; // @[executor.scala 459:20]
    dst_offset_4 <= io_dst_offset_in_4; // @[executor.scala 459:20]
    dst_offset_5 <= io_dst_offset_in_5; // @[executor.scala 459:20]
    dst_offset_6 <= io_dst_offset_in_6; // @[executor.scala 459:20]
    dst_offset_7 <= io_dst_offset_in_7; // @[executor.scala 459:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_header_0 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  phv_header_1 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  phv_header_2 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  phv_header_3 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  phv_header_4 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  phv_header_5 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  phv_header_6 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  phv_header_7 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  phv_header_8 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  phv_header_9 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  phv_header_10 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  phv_header_11 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  phv_header_12 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  phv_header_13 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  phv_header_14 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  phv_header_15 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  phv_next_config_id = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  vliw_0 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  vliw_1 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  vliw_2 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  vliw_3 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  vliw_4 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  vliw_5 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  vliw_6 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  vliw_7 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  field_0 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  field_1 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  field_2 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  field_3 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  field_4 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  field_5 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  field_6 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  field_7 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  mask_0 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  mask_1 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  mask_2 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  mask_3 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  mask_4 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  mask_5 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  mask_6 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  mask_7 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  dst_offset_0 = _RAND_302[5:0];
  _RAND_303 = {1{`RANDOM}};
  dst_offset_1 = _RAND_303[5:0];
  _RAND_304 = {1{`RANDOM}};
  dst_offset_2 = _RAND_304[5:0];
  _RAND_305 = {1{`RANDOM}};
  dst_offset_3 = _RAND_305[5:0];
  _RAND_306 = {1{`RANDOM}};
  dst_offset_4 = _RAND_306[5:0];
  _RAND_307 = {1{`RANDOM}};
  dst_offset_5 = _RAND_307[5:0];
  _RAND_308 = {1{`RANDOM}};
  dst_offset_6 = _RAND_308[5:0];
  _RAND_309 = {1{`RANDOM}};
  dst_offset_7 = _RAND_309[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
