module PrimitiveGetSourcePISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [17:0] io_vliw_in_0,
  input  [17:0] io_vliw_in_1,
  input  [17:0] io_vliw_in_2,
  input  [17:0] io_vliw_in_3,
  input  [17:0] io_vliw_in_4,
  input  [17:0] io_vliw_in_5,
  input  [17:0] io_vliw_in_6,
  input  [17:0] io_vliw_in_7,
  input  [17:0] io_vliw_in_8,
  input  [17:0] io_vliw_in_9,
  input  [17:0] io_vliw_in_10,
  input  [17:0] io_vliw_in_11,
  input  [17:0] io_vliw_in_12,
  input  [17:0] io_vliw_in_13,
  input  [17:0] io_vliw_in_14,
  input  [17:0] io_vliw_in_15,
  input  [17:0] io_vliw_in_16,
  input  [17:0] io_vliw_in_17,
  input  [17:0] io_vliw_in_18,
  input  [17:0] io_vliw_in_19,
  input  [17:0] io_vliw_in_20,
  input  [17:0] io_vliw_in_21,
  input  [17:0] io_vliw_in_22,
  input  [17:0] io_vliw_in_23,
  input  [17:0] io_vliw_in_24,
  input  [17:0] io_vliw_in_25,
  input  [17:0] io_vliw_in_26,
  input  [17:0] io_vliw_in_27,
  input  [17:0] io_vliw_in_28,
  input  [17:0] io_vliw_in_29,
  input  [17:0] io_vliw_in_30,
  input  [17:0] io_vliw_in_31,
  input  [17:0] io_vliw_in_32,
  input  [17:0] io_vliw_in_33,
  input  [17:0] io_vliw_in_34,
  input  [17:0] io_vliw_in_35,
  input  [17:0] io_vliw_in_36,
  input  [17:0] io_vliw_in_37,
  input  [17:0] io_vliw_in_38,
  input  [17:0] io_vliw_in_39,
  input  [17:0] io_vliw_in_40,
  input  [17:0] io_vliw_in_41,
  input  [17:0] io_vliw_in_42,
  input  [17:0] io_vliw_in_43,
  input  [17:0] io_vliw_in_44,
  input  [17:0] io_vliw_in_45,
  input  [17:0] io_vliw_in_46,
  input  [17:0] io_vliw_in_47,
  input  [17:0] io_vliw_in_48,
  input  [17:0] io_vliw_in_49,
  input  [17:0] io_vliw_in_50,
  input  [17:0] io_vliw_in_51,
  input  [17:0] io_vliw_in_52,
  input  [17:0] io_vliw_in_53,
  input  [17:0] io_vliw_in_54,
  input  [17:0] io_vliw_in_55,
  input  [17:0] io_vliw_in_56,
  input  [17:0] io_vliw_in_57,
  input  [17:0] io_vliw_in_58,
  input  [17:0] io_vliw_in_59,
  input  [17:0] io_vliw_in_60,
  input  [17:0] io_vliw_in_61,
  input  [17:0] io_vliw_in_62,
  input  [17:0] io_vliw_in_63,
  input  [17:0] io_vliw_in_64,
  input  [17:0] io_vliw_in_65,
  input  [17:0] io_vliw_in_66,
  input  [17:0] io_vliw_in_67,
  input  [17:0] io_vliw_in_68,
  input  [17:0] io_vliw_in_69,
  input  [14:0] io_nid_in,
  output [14:0] io_nid_out,
  output [1:0]  io_tag_out_0,
  output [1:0]  io_tag_out_1,
  output [1:0]  io_tag_out_2,
  output [1:0]  io_tag_out_3,
  output [1:0]  io_tag_out_4,
  output [1:0]  io_tag_out_5,
  output [1:0]  io_tag_out_6,
  output [1:0]  io_tag_out_7,
  output [1:0]  io_tag_out_8,
  output [1:0]  io_tag_out_9,
  output [1:0]  io_tag_out_10,
  output [1:0]  io_tag_out_11,
  output [1:0]  io_tag_out_12,
  output [1:0]  io_tag_out_13,
  output [1:0]  io_tag_out_14,
  output [1:0]  io_tag_out_15,
  output [1:0]  io_tag_out_16,
  output [1:0]  io_tag_out_17,
  output [1:0]  io_tag_out_18,
  output [1:0]  io_tag_out_19,
  output [1:0]  io_tag_out_20,
  output [1:0]  io_tag_out_21,
  output [1:0]  io_tag_out_22,
  output [1:0]  io_tag_out_23,
  output [1:0]  io_tag_out_24,
  output [1:0]  io_tag_out_25,
  output [1:0]  io_tag_out_26,
  output [1:0]  io_tag_out_27,
  output [1:0]  io_tag_out_28,
  output [1:0]  io_tag_out_29,
  output [1:0]  io_tag_out_30,
  output [1:0]  io_tag_out_31,
  output [1:0]  io_tag_out_32,
  output [1:0]  io_tag_out_33,
  output [1:0]  io_tag_out_34,
  output [1:0]  io_tag_out_35,
  output [1:0]  io_tag_out_36,
  output [1:0]  io_tag_out_37,
  output [1:0]  io_tag_out_38,
  output [1:0]  io_tag_out_39,
  output [1:0]  io_tag_out_40,
  output [1:0]  io_tag_out_41,
  output [1:0]  io_tag_out_42,
  output [1:0]  io_tag_out_43,
  output [1:0]  io_tag_out_44,
  output [1:0]  io_tag_out_45,
  output [1:0]  io_tag_out_46,
  output [1:0]  io_tag_out_47,
  output [1:0]  io_tag_out_48,
  output [1:0]  io_tag_out_49,
  output [1:0]  io_tag_out_50,
  output [1:0]  io_tag_out_51,
  output [1:0]  io_tag_out_52,
  output [1:0]  io_tag_out_53,
  output [1:0]  io_tag_out_54,
  output [1:0]  io_tag_out_55,
  output [1:0]  io_tag_out_56,
  output [1:0]  io_tag_out_57,
  output [1:0]  io_tag_out_58,
  output [1:0]  io_tag_out_59,
  output [1:0]  io_tag_out_60,
  output [1:0]  io_tag_out_61,
  output [1:0]  io_tag_out_62,
  output [1:0]  io_tag_out_63,
  output [1:0]  io_tag_out_64,
  output [1:0]  io_tag_out_65,
  output [1:0]  io_tag_out_66,
  output [1:0]  io_tag_out_67,
  output [1:0]  io_tag_out_68,
  output [1:0]  io_tag_out_69,
  output [7:0]  io_field_set_field8_0,
  output [7:0]  io_field_set_field8_1,
  output [7:0]  io_field_set_field8_2,
  output [7:0]  io_field_set_field8_3,
  output [7:0]  io_field_set_field8_4,
  output [7:0]  io_field_set_field8_5,
  output [7:0]  io_field_set_field8_6,
  output [7:0]  io_field_set_field8_7,
  output [7:0]  io_field_set_field8_8,
  output [7:0]  io_field_set_field8_9,
  output [7:0]  io_field_set_field8_10,
  output [7:0]  io_field_set_field8_11,
  output [7:0]  io_field_set_field8_12,
  output [7:0]  io_field_set_field8_13,
  output [7:0]  io_field_set_field8_14,
  output [7:0]  io_field_set_field8_15,
  output [7:0]  io_field_set_field8_16,
  output [7:0]  io_field_set_field8_17,
  output [7:0]  io_field_set_field8_18,
  output [7:0]  io_field_set_field8_19,
  output [15:0] io_field_set_field16_0,
  output [15:0] io_field_set_field16_1,
  output [15:0] io_field_set_field16_2,
  output [15:0] io_field_set_field16_3,
  output [15:0] io_field_set_field16_4,
  output [15:0] io_field_set_field16_5,
  output [15:0] io_field_set_field16_6,
  output [15:0] io_field_set_field16_7,
  output [15:0] io_field_set_field16_8,
  output [15:0] io_field_set_field16_9,
  output [15:0] io_field_set_field16_10,
  output [15:0] io_field_set_field16_11,
  output [15:0] io_field_set_field16_12,
  output [15:0] io_field_set_field16_13,
  output [15:0] io_field_set_field16_14,
  output [15:0] io_field_set_field16_15,
  output [15:0] io_field_set_field16_16,
  output [15:0] io_field_set_field16_17,
  output [15:0] io_field_set_field16_18,
  output [15:0] io_field_set_field16_19,
  output [15:0] io_field_set_field16_20,
  output [15:0] io_field_set_field16_21,
  output [15:0] io_field_set_field16_22,
  output [15:0] io_field_set_field16_23,
  output [15:0] io_field_set_field16_24,
  output [15:0] io_field_set_field16_25,
  output [15:0] io_field_set_field16_26,
  output [15:0] io_field_set_field16_27,
  output [15:0] io_field_set_field16_28,
  output [15:0] io_field_set_field16_29,
  output [31:0] io_field_set_field32_0,
  output [31:0] io_field_set_field32_1,
  output [31:0] io_field_set_field32_2,
  output [31:0] io_field_set_field32_3,
  output [31:0] io_field_set_field32_4,
  output [31:0] io_field_set_field32_5,
  output [31:0] io_field_set_field32_6,
  output [31:0] io_field_set_field32_7,
  output [31:0] io_field_set_field32_8,
  output [31:0] io_field_set_field32_9,
  output [31:0] io_field_set_field32_10,
  output [31:0] io_field_set_field32_11,
  output [31:0] io_field_set_field32_12,
  output [31:0] io_field_set_field32_13,
  output [31:0] io_field_set_field32_14,
  output [31:0] io_field_set_field32_15,
  output [31:0] io_field_set_field32_16,
  output [31:0] io_field_set_field32_17,
  output [31:0] io_field_set_field32_18,
  output [31:0] io_field_set_field32_19
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_1; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_2; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_3; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_4; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_5; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_6; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_7; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_8; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_9; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_10; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_11; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_12; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_13; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_14; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_15; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_16; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_17; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_18; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_19; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_20; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_21; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_22; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_23; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_24; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_25; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_26; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_27; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_28; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_29; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_30; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_31; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_32; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_33; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_34; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_35; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_36; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_37; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_38; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_39; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_40; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_41; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_42; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_43; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_44; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_45; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_46; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_47; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_48; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_49; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_50; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_51; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_52; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_53; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_54; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_55; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_56; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_57; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_58; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_59; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_60; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_61; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_62; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_63; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_64; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_65; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_66; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_67; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_68; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_69; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_70; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_71; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_72; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_73; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_74; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_75; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_76; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_77; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_78; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_79; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_80; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_81; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_82; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_83; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_84; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_85; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_86; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_87; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_88; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_89; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_90; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_91; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_92; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_93; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_94; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_95; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_96; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_97; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_98; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_99; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_100; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_101; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_102; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_103; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_104; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_105; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_106; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_107; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_108; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_109; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_110; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_111; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_112; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_113; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_114; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_115; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_116; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_117; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_118; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_119; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_120; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_121; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_122; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_123; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_124; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_125; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_126; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_127; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_128; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_129; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_130; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_131; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_132; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_133; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_134; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_135; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_136; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_137; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_138; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_139; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_140; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_141; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_142; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_143; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_144; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_145; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_146; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_147; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_148; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_149; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_150; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_151; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_152; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_153; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_154; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_155; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_156; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_157; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_158; // @[executor_pisa.scala 161:22]
  reg [7:0] phv_data_159; // @[executor_pisa.scala 161:22]
  reg [3:0] phv_next_processor_id; // @[executor_pisa.scala 161:22]
  reg  phv_next_config_id; // @[executor_pisa.scala 161:22]
  reg [7:0] args_0; // @[executor_pisa.scala 165:23]
  reg [7:0] args_1; // @[executor_pisa.scala 165:23]
  reg [7:0] args_2; // @[executor_pisa.scala 165:23]
  reg [7:0] args_3; // @[executor_pisa.scala 165:23]
  reg [7:0] args_4; // @[executor_pisa.scala 165:23]
  reg [7:0] args_5; // @[executor_pisa.scala 165:23]
  reg [7:0] args_6; // @[executor_pisa.scala 165:23]
  reg [17:0] vliw_0; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_1; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_2; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_3; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_4; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_5; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_6; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_7; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_8; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_9; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_10; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_11; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_12; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_13; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_14; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_15; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_16; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_17; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_18; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_19; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_20; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_21; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_22; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_23; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_24; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_25; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_26; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_27; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_28; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_29; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_30; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_31; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_32; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_33; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_34; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_35; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_36; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_37; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_38; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_39; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_40; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_41; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_42; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_43; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_44; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_45; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_46; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_47; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_48; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_49; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_50; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_51; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_52; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_53; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_54; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_55; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_56; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_57; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_58; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_59; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_60; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_61; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_62; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_63; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_64; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_65; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_66; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_67; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_68; // @[executor_pisa.scala 168:23]
  reg [17:0] vliw_69; // @[executor_pisa.scala 168:23]
  reg [14:0] nid; // @[executor_pisa.scala 171:23]
  wire [3:0] opcode = vliw_0[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2 = vliw_0[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset = parameter_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length = parameter_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T = {{1'd0}, args_offset}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset = _total_offset_T[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1 = 3'h1 == total_offset ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2 = 3'h2 == total_offset ? args_2 : _GEN_1; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3 = 3'h3 == total_offset ? args_3 : _GEN_2; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_4 = 3'h4 == total_offset ? args_4 : _GEN_3; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_5 = 3'h5 == total_offset ? args_5 : _GEN_4; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_6 = 3'h6 == total_offset ? args_6 : _GEN_5; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_7 = total_offset < 3'h7 ? _GEN_6 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_0 = 3'h0 < args_length ? _GEN_7 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_9 = opcode == 4'ha ? field_bytes_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_10 = opcode == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_3 = opcode == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_1 = _T_3 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_11 = opcode == 4'h8 | opcode == 4'hb ? parameter_2[7:0] : _GEN_9; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_12 = opcode == 4'h8 | opcode == 4'hb ? _field_tag_T_1 : _GEN_10; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_13 = 14'h0 == parameter_2 ? phv_data_0 : _GEN_11; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_14 = 14'h1 == parameter_2 ? phv_data_1 : _GEN_13; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_15 = 14'h2 == parameter_2 ? phv_data_2 : _GEN_14; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_16 = 14'h3 == parameter_2 ? phv_data_3 : _GEN_15; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_17 = 14'h4 == parameter_2 ? phv_data_4 : _GEN_16; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_18 = 14'h5 == parameter_2 ? phv_data_5 : _GEN_17; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_19 = 14'h6 == parameter_2 ? phv_data_6 : _GEN_18; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_20 = 14'h7 == parameter_2 ? phv_data_7 : _GEN_19; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_21 = 14'h8 == parameter_2 ? phv_data_8 : _GEN_20; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_22 = 14'h9 == parameter_2 ? phv_data_9 : _GEN_21; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_23 = 14'ha == parameter_2 ? phv_data_10 : _GEN_22; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_24 = 14'hb == parameter_2 ? phv_data_11 : _GEN_23; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_25 = 14'hc == parameter_2 ? phv_data_12 : _GEN_24; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_26 = 14'hd == parameter_2 ? phv_data_13 : _GEN_25; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_27 = 14'he == parameter_2 ? phv_data_14 : _GEN_26; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_28 = 14'hf == parameter_2 ? phv_data_15 : _GEN_27; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_29 = 14'h10 == parameter_2 ? phv_data_16 : _GEN_28; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_30 = 14'h11 == parameter_2 ? phv_data_17 : _GEN_29; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_31 = 14'h12 == parameter_2 ? phv_data_18 : _GEN_30; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_32 = 14'h13 == parameter_2 ? phv_data_19 : _GEN_31; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_1 = vliw_1[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_1 = vliw_1[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_1 = parameter_2_1[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_1 = parameter_2_1[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_1 = {{1'd0}, args_offset_1}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_1 = _total_offset_T_1[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_36 = 3'h1 == total_offset_1 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_37 = 3'h2 == total_offset_1 ? args_2 : _GEN_36; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_38 = 3'h3 == total_offset_1 ? args_3 : _GEN_37; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_39 = 3'h4 == total_offset_1 ? args_4 : _GEN_38; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_40 = 3'h5 == total_offset_1 ? args_5 : _GEN_39; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_41 = 3'h6 == total_offset_1 ? args_6 : _GEN_40; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_42 = total_offset_1 < 3'h7 ? _GEN_41 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_1_0 = 3'h0 < args_length_1 ? _GEN_42 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_44 = opcode_1 == 4'ha ? field_bytes_1_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_45 = opcode_1 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_30 = opcode_1 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_3 = _T_30 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_46 = opcode_1 == 4'h8 | opcode_1 == 4'hb ? parameter_2_1[7:0] : _GEN_44; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_47 = opcode_1 == 4'h8 | opcode_1 == 4'hb ? _field_tag_T_3 : _GEN_45; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_48 = 14'h0 == parameter_2_1 ? phv_data_0 : _GEN_46; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_49 = 14'h1 == parameter_2_1 ? phv_data_1 : _GEN_48; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_50 = 14'h2 == parameter_2_1 ? phv_data_2 : _GEN_49; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_51 = 14'h3 == parameter_2_1 ? phv_data_3 : _GEN_50; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_52 = 14'h4 == parameter_2_1 ? phv_data_4 : _GEN_51; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_53 = 14'h5 == parameter_2_1 ? phv_data_5 : _GEN_52; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_54 = 14'h6 == parameter_2_1 ? phv_data_6 : _GEN_53; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_55 = 14'h7 == parameter_2_1 ? phv_data_7 : _GEN_54; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_56 = 14'h8 == parameter_2_1 ? phv_data_8 : _GEN_55; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_57 = 14'h9 == parameter_2_1 ? phv_data_9 : _GEN_56; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_58 = 14'ha == parameter_2_1 ? phv_data_10 : _GEN_57; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_59 = 14'hb == parameter_2_1 ? phv_data_11 : _GEN_58; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_60 = 14'hc == parameter_2_1 ? phv_data_12 : _GEN_59; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_61 = 14'hd == parameter_2_1 ? phv_data_13 : _GEN_60; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_62 = 14'he == parameter_2_1 ? phv_data_14 : _GEN_61; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_63 = 14'hf == parameter_2_1 ? phv_data_15 : _GEN_62; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_64 = 14'h10 == parameter_2_1 ? phv_data_16 : _GEN_63; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_65 = 14'h11 == parameter_2_1 ? phv_data_17 : _GEN_64; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_66 = 14'h12 == parameter_2_1 ? phv_data_18 : _GEN_65; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_67 = 14'h13 == parameter_2_1 ? phv_data_19 : _GEN_66; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_2 = vliw_2[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_2 = vliw_2[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_2 = parameter_2_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_2 = parameter_2_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_2 = {{1'd0}, args_offset_2}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_2 = _total_offset_T_2[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_71 = 3'h1 == total_offset_2 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_72 = 3'h2 == total_offset_2 ? args_2 : _GEN_71; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_73 = 3'h3 == total_offset_2 ? args_3 : _GEN_72; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_74 = 3'h4 == total_offset_2 ? args_4 : _GEN_73; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_75 = 3'h5 == total_offset_2 ? args_5 : _GEN_74; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_76 = 3'h6 == total_offset_2 ? args_6 : _GEN_75; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_77 = total_offset_2 < 3'h7 ? _GEN_76 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_2_0 = 3'h0 < args_length_2 ? _GEN_77 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_79 = opcode_2 == 4'ha ? field_bytes_2_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_80 = opcode_2 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_57 = opcode_2 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_5 = _T_57 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_81 = opcode_2 == 4'h8 | opcode_2 == 4'hb ? parameter_2_2[7:0] : _GEN_79; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_82 = opcode_2 == 4'h8 | opcode_2 == 4'hb ? _field_tag_T_5 : _GEN_80; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_83 = 14'h0 == parameter_2_2 ? phv_data_0 : _GEN_81; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_84 = 14'h1 == parameter_2_2 ? phv_data_1 : _GEN_83; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_85 = 14'h2 == parameter_2_2 ? phv_data_2 : _GEN_84; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_86 = 14'h3 == parameter_2_2 ? phv_data_3 : _GEN_85; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_87 = 14'h4 == parameter_2_2 ? phv_data_4 : _GEN_86; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_88 = 14'h5 == parameter_2_2 ? phv_data_5 : _GEN_87; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_89 = 14'h6 == parameter_2_2 ? phv_data_6 : _GEN_88; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_90 = 14'h7 == parameter_2_2 ? phv_data_7 : _GEN_89; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_91 = 14'h8 == parameter_2_2 ? phv_data_8 : _GEN_90; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_92 = 14'h9 == parameter_2_2 ? phv_data_9 : _GEN_91; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_93 = 14'ha == parameter_2_2 ? phv_data_10 : _GEN_92; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_94 = 14'hb == parameter_2_2 ? phv_data_11 : _GEN_93; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_95 = 14'hc == parameter_2_2 ? phv_data_12 : _GEN_94; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_96 = 14'hd == parameter_2_2 ? phv_data_13 : _GEN_95; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_97 = 14'he == parameter_2_2 ? phv_data_14 : _GEN_96; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_98 = 14'hf == parameter_2_2 ? phv_data_15 : _GEN_97; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_99 = 14'h10 == parameter_2_2 ? phv_data_16 : _GEN_98; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_100 = 14'h11 == parameter_2_2 ? phv_data_17 : _GEN_99; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_101 = 14'h12 == parameter_2_2 ? phv_data_18 : _GEN_100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_102 = 14'h13 == parameter_2_2 ? phv_data_19 : _GEN_101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_3 = vliw_3[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_3 = vliw_3[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_3 = parameter_2_3[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_3 = parameter_2_3[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_3 = {{1'd0}, args_offset_3}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_3 = _total_offset_T_3[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_106 = 3'h1 == total_offset_3 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_107 = 3'h2 == total_offset_3 ? args_2 : _GEN_106; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_108 = 3'h3 == total_offset_3 ? args_3 : _GEN_107; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_109 = 3'h4 == total_offset_3 ? args_4 : _GEN_108; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_110 = 3'h5 == total_offset_3 ? args_5 : _GEN_109; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_111 = 3'h6 == total_offset_3 ? args_6 : _GEN_110; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_112 = total_offset_3 < 3'h7 ? _GEN_111 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_3_0 = 3'h0 < args_length_3 ? _GEN_112 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_114 = opcode_3 == 4'ha ? field_bytes_3_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_115 = opcode_3 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_84 = opcode_3 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_7 = _T_84 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_116 = opcode_3 == 4'h8 | opcode_3 == 4'hb ? parameter_2_3[7:0] : _GEN_114; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_117 = opcode_3 == 4'h8 | opcode_3 == 4'hb ? _field_tag_T_7 : _GEN_115; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_118 = 14'h0 == parameter_2_3 ? phv_data_0 : _GEN_116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_119 = 14'h1 == parameter_2_3 ? phv_data_1 : _GEN_118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_120 = 14'h2 == parameter_2_3 ? phv_data_2 : _GEN_119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_121 = 14'h3 == parameter_2_3 ? phv_data_3 : _GEN_120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_122 = 14'h4 == parameter_2_3 ? phv_data_4 : _GEN_121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_123 = 14'h5 == parameter_2_3 ? phv_data_5 : _GEN_122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_124 = 14'h6 == parameter_2_3 ? phv_data_6 : _GEN_123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_125 = 14'h7 == parameter_2_3 ? phv_data_7 : _GEN_124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_126 = 14'h8 == parameter_2_3 ? phv_data_8 : _GEN_125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_127 = 14'h9 == parameter_2_3 ? phv_data_9 : _GEN_126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_128 = 14'ha == parameter_2_3 ? phv_data_10 : _GEN_127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_129 = 14'hb == parameter_2_3 ? phv_data_11 : _GEN_128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_130 = 14'hc == parameter_2_3 ? phv_data_12 : _GEN_129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_131 = 14'hd == parameter_2_3 ? phv_data_13 : _GEN_130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_132 = 14'he == parameter_2_3 ? phv_data_14 : _GEN_131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_133 = 14'hf == parameter_2_3 ? phv_data_15 : _GEN_132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_134 = 14'h10 == parameter_2_3 ? phv_data_16 : _GEN_133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_135 = 14'h11 == parameter_2_3 ? phv_data_17 : _GEN_134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_136 = 14'h12 == parameter_2_3 ? phv_data_18 : _GEN_135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_137 = 14'h13 == parameter_2_3 ? phv_data_19 : _GEN_136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_4 = vliw_4[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_4 = vliw_4[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_4 = parameter_2_4[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_4 = parameter_2_4[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_4 = {{1'd0}, args_offset_4}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_4 = _total_offset_T_4[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_141 = 3'h1 == total_offset_4 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_142 = 3'h2 == total_offset_4 ? args_2 : _GEN_141; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_143 = 3'h3 == total_offset_4 ? args_3 : _GEN_142; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_144 = 3'h4 == total_offset_4 ? args_4 : _GEN_143; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_145 = 3'h5 == total_offset_4 ? args_5 : _GEN_144; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_146 = 3'h6 == total_offset_4 ? args_6 : _GEN_145; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_147 = total_offset_4 < 3'h7 ? _GEN_146 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_4_0 = 3'h0 < args_length_4 ? _GEN_147 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_149 = opcode_4 == 4'ha ? field_bytes_4_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_150 = opcode_4 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_111 = opcode_4 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_9 = _T_111 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_151 = opcode_4 == 4'h8 | opcode_4 == 4'hb ? parameter_2_4[7:0] : _GEN_149; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_152 = opcode_4 == 4'h8 | opcode_4 == 4'hb ? _field_tag_T_9 : _GEN_150; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_153 = 14'h0 == parameter_2_4 ? phv_data_0 : _GEN_151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_154 = 14'h1 == parameter_2_4 ? phv_data_1 : _GEN_153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_155 = 14'h2 == parameter_2_4 ? phv_data_2 : _GEN_154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_156 = 14'h3 == parameter_2_4 ? phv_data_3 : _GEN_155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_157 = 14'h4 == parameter_2_4 ? phv_data_4 : _GEN_156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_158 = 14'h5 == parameter_2_4 ? phv_data_5 : _GEN_157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_159 = 14'h6 == parameter_2_4 ? phv_data_6 : _GEN_158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_160 = 14'h7 == parameter_2_4 ? phv_data_7 : _GEN_159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_161 = 14'h8 == parameter_2_4 ? phv_data_8 : _GEN_160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_162 = 14'h9 == parameter_2_4 ? phv_data_9 : _GEN_161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_163 = 14'ha == parameter_2_4 ? phv_data_10 : _GEN_162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_164 = 14'hb == parameter_2_4 ? phv_data_11 : _GEN_163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_165 = 14'hc == parameter_2_4 ? phv_data_12 : _GEN_164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_166 = 14'hd == parameter_2_4 ? phv_data_13 : _GEN_165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_167 = 14'he == parameter_2_4 ? phv_data_14 : _GEN_166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_168 = 14'hf == parameter_2_4 ? phv_data_15 : _GEN_167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_169 = 14'h10 == parameter_2_4 ? phv_data_16 : _GEN_168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_170 = 14'h11 == parameter_2_4 ? phv_data_17 : _GEN_169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_171 = 14'h12 == parameter_2_4 ? phv_data_18 : _GEN_170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_172 = 14'h13 == parameter_2_4 ? phv_data_19 : _GEN_171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_5 = vliw_5[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_5 = vliw_5[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_5 = parameter_2_5[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_5 = parameter_2_5[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_5 = {{1'd0}, args_offset_5}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_5 = _total_offset_T_5[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_176 = 3'h1 == total_offset_5 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_177 = 3'h2 == total_offset_5 ? args_2 : _GEN_176; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_178 = 3'h3 == total_offset_5 ? args_3 : _GEN_177; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_179 = 3'h4 == total_offset_5 ? args_4 : _GEN_178; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_180 = 3'h5 == total_offset_5 ? args_5 : _GEN_179; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_181 = 3'h6 == total_offset_5 ? args_6 : _GEN_180; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_182 = total_offset_5 < 3'h7 ? _GEN_181 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_5_0 = 3'h0 < args_length_5 ? _GEN_182 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_184 = opcode_5 == 4'ha ? field_bytes_5_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_185 = opcode_5 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_138 = opcode_5 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_11 = _T_138 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_186 = opcode_5 == 4'h8 | opcode_5 == 4'hb ? parameter_2_5[7:0] : _GEN_184; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_187 = opcode_5 == 4'h8 | opcode_5 == 4'hb ? _field_tag_T_11 : _GEN_185; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_188 = 14'h0 == parameter_2_5 ? phv_data_0 : _GEN_186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_189 = 14'h1 == parameter_2_5 ? phv_data_1 : _GEN_188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_190 = 14'h2 == parameter_2_5 ? phv_data_2 : _GEN_189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_191 = 14'h3 == parameter_2_5 ? phv_data_3 : _GEN_190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_192 = 14'h4 == parameter_2_5 ? phv_data_4 : _GEN_191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_193 = 14'h5 == parameter_2_5 ? phv_data_5 : _GEN_192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_194 = 14'h6 == parameter_2_5 ? phv_data_6 : _GEN_193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_195 = 14'h7 == parameter_2_5 ? phv_data_7 : _GEN_194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_196 = 14'h8 == parameter_2_5 ? phv_data_8 : _GEN_195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_197 = 14'h9 == parameter_2_5 ? phv_data_9 : _GEN_196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_198 = 14'ha == parameter_2_5 ? phv_data_10 : _GEN_197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_199 = 14'hb == parameter_2_5 ? phv_data_11 : _GEN_198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_200 = 14'hc == parameter_2_5 ? phv_data_12 : _GEN_199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_201 = 14'hd == parameter_2_5 ? phv_data_13 : _GEN_200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_202 = 14'he == parameter_2_5 ? phv_data_14 : _GEN_201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_203 = 14'hf == parameter_2_5 ? phv_data_15 : _GEN_202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_204 = 14'h10 == parameter_2_5 ? phv_data_16 : _GEN_203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_205 = 14'h11 == parameter_2_5 ? phv_data_17 : _GEN_204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_206 = 14'h12 == parameter_2_5 ? phv_data_18 : _GEN_205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_207 = 14'h13 == parameter_2_5 ? phv_data_19 : _GEN_206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_6 = vliw_6[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_6 = vliw_6[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_6 = parameter_2_6[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_6 = parameter_2_6[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_6 = {{1'd0}, args_offset_6}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_6 = _total_offset_T_6[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_211 = 3'h1 == total_offset_6 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_212 = 3'h2 == total_offset_6 ? args_2 : _GEN_211; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_213 = 3'h3 == total_offset_6 ? args_3 : _GEN_212; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_214 = 3'h4 == total_offset_6 ? args_4 : _GEN_213; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_215 = 3'h5 == total_offset_6 ? args_5 : _GEN_214; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_216 = 3'h6 == total_offset_6 ? args_6 : _GEN_215; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_217 = total_offset_6 < 3'h7 ? _GEN_216 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_6_0 = 3'h0 < args_length_6 ? _GEN_217 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_219 = opcode_6 == 4'ha ? field_bytes_6_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_220 = opcode_6 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_165 = opcode_6 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_13 = _T_165 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_221 = opcode_6 == 4'h8 | opcode_6 == 4'hb ? parameter_2_6[7:0] : _GEN_219; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_222 = opcode_6 == 4'h8 | opcode_6 == 4'hb ? _field_tag_T_13 : _GEN_220; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_223 = 14'h0 == parameter_2_6 ? phv_data_0 : _GEN_221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_224 = 14'h1 == parameter_2_6 ? phv_data_1 : _GEN_223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_225 = 14'h2 == parameter_2_6 ? phv_data_2 : _GEN_224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_226 = 14'h3 == parameter_2_6 ? phv_data_3 : _GEN_225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_227 = 14'h4 == parameter_2_6 ? phv_data_4 : _GEN_226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_228 = 14'h5 == parameter_2_6 ? phv_data_5 : _GEN_227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_229 = 14'h6 == parameter_2_6 ? phv_data_6 : _GEN_228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_230 = 14'h7 == parameter_2_6 ? phv_data_7 : _GEN_229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_231 = 14'h8 == parameter_2_6 ? phv_data_8 : _GEN_230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_232 = 14'h9 == parameter_2_6 ? phv_data_9 : _GEN_231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_233 = 14'ha == parameter_2_6 ? phv_data_10 : _GEN_232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_234 = 14'hb == parameter_2_6 ? phv_data_11 : _GEN_233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_235 = 14'hc == parameter_2_6 ? phv_data_12 : _GEN_234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_236 = 14'hd == parameter_2_6 ? phv_data_13 : _GEN_235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_237 = 14'he == parameter_2_6 ? phv_data_14 : _GEN_236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_238 = 14'hf == parameter_2_6 ? phv_data_15 : _GEN_237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_239 = 14'h10 == parameter_2_6 ? phv_data_16 : _GEN_238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_240 = 14'h11 == parameter_2_6 ? phv_data_17 : _GEN_239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_241 = 14'h12 == parameter_2_6 ? phv_data_18 : _GEN_240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_242 = 14'h13 == parameter_2_6 ? phv_data_19 : _GEN_241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_7 = vliw_7[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_7 = vliw_7[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_7 = parameter_2_7[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_7 = parameter_2_7[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_7 = {{1'd0}, args_offset_7}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_7 = _total_offset_T_7[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_246 = 3'h1 == total_offset_7 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_247 = 3'h2 == total_offset_7 ? args_2 : _GEN_246; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_248 = 3'h3 == total_offset_7 ? args_3 : _GEN_247; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_249 = 3'h4 == total_offset_7 ? args_4 : _GEN_248; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_250 = 3'h5 == total_offset_7 ? args_5 : _GEN_249; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_251 = 3'h6 == total_offset_7 ? args_6 : _GEN_250; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_252 = total_offset_7 < 3'h7 ? _GEN_251 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_7_0 = 3'h0 < args_length_7 ? _GEN_252 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_254 = opcode_7 == 4'ha ? field_bytes_7_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_255 = opcode_7 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_192 = opcode_7 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_15 = _T_192 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_256 = opcode_7 == 4'h8 | opcode_7 == 4'hb ? parameter_2_7[7:0] : _GEN_254; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_257 = opcode_7 == 4'h8 | opcode_7 == 4'hb ? _field_tag_T_15 : _GEN_255; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_258 = 14'h0 == parameter_2_7 ? phv_data_0 : _GEN_256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_259 = 14'h1 == parameter_2_7 ? phv_data_1 : _GEN_258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_260 = 14'h2 == parameter_2_7 ? phv_data_2 : _GEN_259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_261 = 14'h3 == parameter_2_7 ? phv_data_3 : _GEN_260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_262 = 14'h4 == parameter_2_7 ? phv_data_4 : _GEN_261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_263 = 14'h5 == parameter_2_7 ? phv_data_5 : _GEN_262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_264 = 14'h6 == parameter_2_7 ? phv_data_6 : _GEN_263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_265 = 14'h7 == parameter_2_7 ? phv_data_7 : _GEN_264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_266 = 14'h8 == parameter_2_7 ? phv_data_8 : _GEN_265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_267 = 14'h9 == parameter_2_7 ? phv_data_9 : _GEN_266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_268 = 14'ha == parameter_2_7 ? phv_data_10 : _GEN_267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_269 = 14'hb == parameter_2_7 ? phv_data_11 : _GEN_268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_270 = 14'hc == parameter_2_7 ? phv_data_12 : _GEN_269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_271 = 14'hd == parameter_2_7 ? phv_data_13 : _GEN_270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_272 = 14'he == parameter_2_7 ? phv_data_14 : _GEN_271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_273 = 14'hf == parameter_2_7 ? phv_data_15 : _GEN_272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_274 = 14'h10 == parameter_2_7 ? phv_data_16 : _GEN_273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_275 = 14'h11 == parameter_2_7 ? phv_data_17 : _GEN_274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_276 = 14'h12 == parameter_2_7 ? phv_data_18 : _GEN_275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_277 = 14'h13 == parameter_2_7 ? phv_data_19 : _GEN_276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_8 = vliw_8[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_8 = vliw_8[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_8 = parameter_2_8[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_8 = parameter_2_8[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_8 = {{1'd0}, args_offset_8}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_8 = _total_offset_T_8[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_281 = 3'h1 == total_offset_8 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_282 = 3'h2 == total_offset_8 ? args_2 : _GEN_281; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_283 = 3'h3 == total_offset_8 ? args_3 : _GEN_282; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_284 = 3'h4 == total_offset_8 ? args_4 : _GEN_283; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_285 = 3'h5 == total_offset_8 ? args_5 : _GEN_284; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_286 = 3'h6 == total_offset_8 ? args_6 : _GEN_285; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_287 = total_offset_8 < 3'h7 ? _GEN_286 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_8_0 = 3'h0 < args_length_8 ? _GEN_287 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_289 = opcode_8 == 4'ha ? field_bytes_8_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_290 = opcode_8 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_219 = opcode_8 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_17 = _T_219 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_291 = opcode_8 == 4'h8 | opcode_8 == 4'hb ? parameter_2_8[7:0] : _GEN_289; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_292 = opcode_8 == 4'h8 | opcode_8 == 4'hb ? _field_tag_T_17 : _GEN_290; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_293 = 14'h0 == parameter_2_8 ? phv_data_0 : _GEN_291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_294 = 14'h1 == parameter_2_8 ? phv_data_1 : _GEN_293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_295 = 14'h2 == parameter_2_8 ? phv_data_2 : _GEN_294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_296 = 14'h3 == parameter_2_8 ? phv_data_3 : _GEN_295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_297 = 14'h4 == parameter_2_8 ? phv_data_4 : _GEN_296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_298 = 14'h5 == parameter_2_8 ? phv_data_5 : _GEN_297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_299 = 14'h6 == parameter_2_8 ? phv_data_6 : _GEN_298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_300 = 14'h7 == parameter_2_8 ? phv_data_7 : _GEN_299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_301 = 14'h8 == parameter_2_8 ? phv_data_8 : _GEN_300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_302 = 14'h9 == parameter_2_8 ? phv_data_9 : _GEN_301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_303 = 14'ha == parameter_2_8 ? phv_data_10 : _GEN_302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_304 = 14'hb == parameter_2_8 ? phv_data_11 : _GEN_303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_305 = 14'hc == parameter_2_8 ? phv_data_12 : _GEN_304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_306 = 14'hd == parameter_2_8 ? phv_data_13 : _GEN_305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_307 = 14'he == parameter_2_8 ? phv_data_14 : _GEN_306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_308 = 14'hf == parameter_2_8 ? phv_data_15 : _GEN_307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_309 = 14'h10 == parameter_2_8 ? phv_data_16 : _GEN_308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_310 = 14'h11 == parameter_2_8 ? phv_data_17 : _GEN_309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_311 = 14'h12 == parameter_2_8 ? phv_data_18 : _GEN_310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_312 = 14'h13 == parameter_2_8 ? phv_data_19 : _GEN_311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_9 = vliw_9[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_9 = vliw_9[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_9 = parameter_2_9[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_9 = parameter_2_9[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_9 = {{1'd0}, args_offset_9}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_9 = _total_offset_T_9[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_316 = 3'h1 == total_offset_9 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_317 = 3'h2 == total_offset_9 ? args_2 : _GEN_316; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_318 = 3'h3 == total_offset_9 ? args_3 : _GEN_317; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_319 = 3'h4 == total_offset_9 ? args_4 : _GEN_318; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_320 = 3'h5 == total_offset_9 ? args_5 : _GEN_319; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_321 = 3'h6 == total_offset_9 ? args_6 : _GEN_320; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_322 = total_offset_9 < 3'h7 ? _GEN_321 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_9_0 = 3'h0 < args_length_9 ? _GEN_322 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_324 = opcode_9 == 4'ha ? field_bytes_9_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_325 = opcode_9 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_246 = opcode_9 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_19 = _T_246 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_326 = opcode_9 == 4'h8 | opcode_9 == 4'hb ? parameter_2_9[7:0] : _GEN_324; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_327 = opcode_9 == 4'h8 | opcode_9 == 4'hb ? _field_tag_T_19 : _GEN_325; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_328 = 14'h0 == parameter_2_9 ? phv_data_0 : _GEN_326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_329 = 14'h1 == parameter_2_9 ? phv_data_1 : _GEN_328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_330 = 14'h2 == parameter_2_9 ? phv_data_2 : _GEN_329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_331 = 14'h3 == parameter_2_9 ? phv_data_3 : _GEN_330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_332 = 14'h4 == parameter_2_9 ? phv_data_4 : _GEN_331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_333 = 14'h5 == parameter_2_9 ? phv_data_5 : _GEN_332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_334 = 14'h6 == parameter_2_9 ? phv_data_6 : _GEN_333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_335 = 14'h7 == parameter_2_9 ? phv_data_7 : _GEN_334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_336 = 14'h8 == parameter_2_9 ? phv_data_8 : _GEN_335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_337 = 14'h9 == parameter_2_9 ? phv_data_9 : _GEN_336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_338 = 14'ha == parameter_2_9 ? phv_data_10 : _GEN_337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_339 = 14'hb == parameter_2_9 ? phv_data_11 : _GEN_338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_340 = 14'hc == parameter_2_9 ? phv_data_12 : _GEN_339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_341 = 14'hd == parameter_2_9 ? phv_data_13 : _GEN_340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_342 = 14'he == parameter_2_9 ? phv_data_14 : _GEN_341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_343 = 14'hf == parameter_2_9 ? phv_data_15 : _GEN_342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_344 = 14'h10 == parameter_2_9 ? phv_data_16 : _GEN_343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_345 = 14'h11 == parameter_2_9 ? phv_data_17 : _GEN_344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_346 = 14'h12 == parameter_2_9 ? phv_data_18 : _GEN_345; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_347 = 14'h13 == parameter_2_9 ? phv_data_19 : _GEN_346; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_10 = vliw_10[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_10 = vliw_10[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_10 = parameter_2_10[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_10 = parameter_2_10[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_10 = {{1'd0}, args_offset_10}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_10 = _total_offset_T_10[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_351 = 3'h1 == total_offset_10 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_352 = 3'h2 == total_offset_10 ? args_2 : _GEN_351; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_353 = 3'h3 == total_offset_10 ? args_3 : _GEN_352; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_354 = 3'h4 == total_offset_10 ? args_4 : _GEN_353; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_355 = 3'h5 == total_offset_10 ? args_5 : _GEN_354; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_356 = 3'h6 == total_offset_10 ? args_6 : _GEN_355; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_357 = total_offset_10 < 3'h7 ? _GEN_356 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_10_0 = 3'h0 < args_length_10 ? _GEN_357 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_359 = opcode_10 == 4'ha ? field_bytes_10_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_360 = opcode_10 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_273 = opcode_10 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_21 = _T_273 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_361 = opcode_10 == 4'h8 | opcode_10 == 4'hb ? parameter_2_10[7:0] : _GEN_359; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_362 = opcode_10 == 4'h8 | opcode_10 == 4'hb ? _field_tag_T_21 : _GEN_360; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_363 = 14'h0 == parameter_2_10 ? phv_data_0 : _GEN_361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_364 = 14'h1 == parameter_2_10 ? phv_data_1 : _GEN_363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_365 = 14'h2 == parameter_2_10 ? phv_data_2 : _GEN_364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_366 = 14'h3 == parameter_2_10 ? phv_data_3 : _GEN_365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_367 = 14'h4 == parameter_2_10 ? phv_data_4 : _GEN_366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_368 = 14'h5 == parameter_2_10 ? phv_data_5 : _GEN_367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_369 = 14'h6 == parameter_2_10 ? phv_data_6 : _GEN_368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_370 = 14'h7 == parameter_2_10 ? phv_data_7 : _GEN_369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_371 = 14'h8 == parameter_2_10 ? phv_data_8 : _GEN_370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_372 = 14'h9 == parameter_2_10 ? phv_data_9 : _GEN_371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_373 = 14'ha == parameter_2_10 ? phv_data_10 : _GEN_372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_374 = 14'hb == parameter_2_10 ? phv_data_11 : _GEN_373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_375 = 14'hc == parameter_2_10 ? phv_data_12 : _GEN_374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_376 = 14'hd == parameter_2_10 ? phv_data_13 : _GEN_375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_377 = 14'he == parameter_2_10 ? phv_data_14 : _GEN_376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_378 = 14'hf == parameter_2_10 ? phv_data_15 : _GEN_377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_379 = 14'h10 == parameter_2_10 ? phv_data_16 : _GEN_378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_380 = 14'h11 == parameter_2_10 ? phv_data_17 : _GEN_379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_381 = 14'h12 == parameter_2_10 ? phv_data_18 : _GEN_380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_382 = 14'h13 == parameter_2_10 ? phv_data_19 : _GEN_381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_11 = vliw_11[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_11 = vliw_11[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_11 = parameter_2_11[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_11 = parameter_2_11[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_11 = {{1'd0}, args_offset_11}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_11 = _total_offset_T_11[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_386 = 3'h1 == total_offset_11 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_387 = 3'h2 == total_offset_11 ? args_2 : _GEN_386; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_388 = 3'h3 == total_offset_11 ? args_3 : _GEN_387; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_389 = 3'h4 == total_offset_11 ? args_4 : _GEN_388; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_390 = 3'h5 == total_offset_11 ? args_5 : _GEN_389; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_391 = 3'h6 == total_offset_11 ? args_6 : _GEN_390; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_392 = total_offset_11 < 3'h7 ? _GEN_391 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_11_0 = 3'h0 < args_length_11 ? _GEN_392 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_394 = opcode_11 == 4'ha ? field_bytes_11_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_395 = opcode_11 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_300 = opcode_11 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_23 = _T_300 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_396 = opcode_11 == 4'h8 | opcode_11 == 4'hb ? parameter_2_11[7:0] : _GEN_394; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_397 = opcode_11 == 4'h8 | opcode_11 == 4'hb ? _field_tag_T_23 : _GEN_395; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_398 = 14'h0 == parameter_2_11 ? phv_data_0 : _GEN_396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_399 = 14'h1 == parameter_2_11 ? phv_data_1 : _GEN_398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_400 = 14'h2 == parameter_2_11 ? phv_data_2 : _GEN_399; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_401 = 14'h3 == parameter_2_11 ? phv_data_3 : _GEN_400; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_402 = 14'h4 == parameter_2_11 ? phv_data_4 : _GEN_401; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_403 = 14'h5 == parameter_2_11 ? phv_data_5 : _GEN_402; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_404 = 14'h6 == parameter_2_11 ? phv_data_6 : _GEN_403; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_405 = 14'h7 == parameter_2_11 ? phv_data_7 : _GEN_404; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_406 = 14'h8 == parameter_2_11 ? phv_data_8 : _GEN_405; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_407 = 14'h9 == parameter_2_11 ? phv_data_9 : _GEN_406; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_408 = 14'ha == parameter_2_11 ? phv_data_10 : _GEN_407; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_409 = 14'hb == parameter_2_11 ? phv_data_11 : _GEN_408; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_410 = 14'hc == parameter_2_11 ? phv_data_12 : _GEN_409; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_411 = 14'hd == parameter_2_11 ? phv_data_13 : _GEN_410; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_412 = 14'he == parameter_2_11 ? phv_data_14 : _GEN_411; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_413 = 14'hf == parameter_2_11 ? phv_data_15 : _GEN_412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_414 = 14'h10 == parameter_2_11 ? phv_data_16 : _GEN_413; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_415 = 14'h11 == parameter_2_11 ? phv_data_17 : _GEN_414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_416 = 14'h12 == parameter_2_11 ? phv_data_18 : _GEN_415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_417 = 14'h13 == parameter_2_11 ? phv_data_19 : _GEN_416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_12 = vliw_12[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_12 = vliw_12[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_12 = parameter_2_12[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_12 = parameter_2_12[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_12 = {{1'd0}, args_offset_12}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_12 = _total_offset_T_12[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_421 = 3'h1 == total_offset_12 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_422 = 3'h2 == total_offset_12 ? args_2 : _GEN_421; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_423 = 3'h3 == total_offset_12 ? args_3 : _GEN_422; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_424 = 3'h4 == total_offset_12 ? args_4 : _GEN_423; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_425 = 3'h5 == total_offset_12 ? args_5 : _GEN_424; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_426 = 3'h6 == total_offset_12 ? args_6 : _GEN_425; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_427 = total_offset_12 < 3'h7 ? _GEN_426 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_12_0 = 3'h0 < args_length_12 ? _GEN_427 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_429 = opcode_12 == 4'ha ? field_bytes_12_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_430 = opcode_12 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_327 = opcode_12 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_25 = _T_327 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_431 = opcode_12 == 4'h8 | opcode_12 == 4'hb ? parameter_2_12[7:0] : _GEN_429; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_432 = opcode_12 == 4'h8 | opcode_12 == 4'hb ? _field_tag_T_25 : _GEN_430; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_433 = 14'h0 == parameter_2_12 ? phv_data_0 : _GEN_431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_434 = 14'h1 == parameter_2_12 ? phv_data_1 : _GEN_433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_435 = 14'h2 == parameter_2_12 ? phv_data_2 : _GEN_434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_436 = 14'h3 == parameter_2_12 ? phv_data_3 : _GEN_435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_437 = 14'h4 == parameter_2_12 ? phv_data_4 : _GEN_436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_438 = 14'h5 == parameter_2_12 ? phv_data_5 : _GEN_437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_439 = 14'h6 == parameter_2_12 ? phv_data_6 : _GEN_438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_440 = 14'h7 == parameter_2_12 ? phv_data_7 : _GEN_439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_441 = 14'h8 == parameter_2_12 ? phv_data_8 : _GEN_440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_442 = 14'h9 == parameter_2_12 ? phv_data_9 : _GEN_441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_443 = 14'ha == parameter_2_12 ? phv_data_10 : _GEN_442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_444 = 14'hb == parameter_2_12 ? phv_data_11 : _GEN_443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_445 = 14'hc == parameter_2_12 ? phv_data_12 : _GEN_444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_446 = 14'hd == parameter_2_12 ? phv_data_13 : _GEN_445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_447 = 14'he == parameter_2_12 ? phv_data_14 : _GEN_446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_448 = 14'hf == parameter_2_12 ? phv_data_15 : _GEN_447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_449 = 14'h10 == parameter_2_12 ? phv_data_16 : _GEN_448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_450 = 14'h11 == parameter_2_12 ? phv_data_17 : _GEN_449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_451 = 14'h12 == parameter_2_12 ? phv_data_18 : _GEN_450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_452 = 14'h13 == parameter_2_12 ? phv_data_19 : _GEN_451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_13 = vliw_13[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_13 = vliw_13[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_13 = parameter_2_13[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_13 = parameter_2_13[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_13 = {{1'd0}, args_offset_13}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_13 = _total_offset_T_13[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_456 = 3'h1 == total_offset_13 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_457 = 3'h2 == total_offset_13 ? args_2 : _GEN_456; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_458 = 3'h3 == total_offset_13 ? args_3 : _GEN_457; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_459 = 3'h4 == total_offset_13 ? args_4 : _GEN_458; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_460 = 3'h5 == total_offset_13 ? args_5 : _GEN_459; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_461 = 3'h6 == total_offset_13 ? args_6 : _GEN_460; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_462 = total_offset_13 < 3'h7 ? _GEN_461 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_13_0 = 3'h0 < args_length_13 ? _GEN_462 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_464 = opcode_13 == 4'ha ? field_bytes_13_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_465 = opcode_13 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_354 = opcode_13 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_27 = _T_354 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_466 = opcode_13 == 4'h8 | opcode_13 == 4'hb ? parameter_2_13[7:0] : _GEN_464; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_467 = opcode_13 == 4'h8 | opcode_13 == 4'hb ? _field_tag_T_27 : _GEN_465; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_468 = 14'h0 == parameter_2_13 ? phv_data_0 : _GEN_466; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_469 = 14'h1 == parameter_2_13 ? phv_data_1 : _GEN_468; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_470 = 14'h2 == parameter_2_13 ? phv_data_2 : _GEN_469; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_471 = 14'h3 == parameter_2_13 ? phv_data_3 : _GEN_470; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_472 = 14'h4 == parameter_2_13 ? phv_data_4 : _GEN_471; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_473 = 14'h5 == parameter_2_13 ? phv_data_5 : _GEN_472; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_474 = 14'h6 == parameter_2_13 ? phv_data_6 : _GEN_473; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_475 = 14'h7 == parameter_2_13 ? phv_data_7 : _GEN_474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_476 = 14'h8 == parameter_2_13 ? phv_data_8 : _GEN_475; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_477 = 14'h9 == parameter_2_13 ? phv_data_9 : _GEN_476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_478 = 14'ha == parameter_2_13 ? phv_data_10 : _GEN_477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_479 = 14'hb == parameter_2_13 ? phv_data_11 : _GEN_478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_480 = 14'hc == parameter_2_13 ? phv_data_12 : _GEN_479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_481 = 14'hd == parameter_2_13 ? phv_data_13 : _GEN_480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_482 = 14'he == parameter_2_13 ? phv_data_14 : _GEN_481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_483 = 14'hf == parameter_2_13 ? phv_data_15 : _GEN_482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_484 = 14'h10 == parameter_2_13 ? phv_data_16 : _GEN_483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_485 = 14'h11 == parameter_2_13 ? phv_data_17 : _GEN_484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_486 = 14'h12 == parameter_2_13 ? phv_data_18 : _GEN_485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_487 = 14'h13 == parameter_2_13 ? phv_data_19 : _GEN_486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_14 = vliw_14[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_14 = vliw_14[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_14 = parameter_2_14[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_14 = parameter_2_14[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_14 = {{1'd0}, args_offset_14}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_14 = _total_offset_T_14[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_491 = 3'h1 == total_offset_14 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_492 = 3'h2 == total_offset_14 ? args_2 : _GEN_491; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_493 = 3'h3 == total_offset_14 ? args_3 : _GEN_492; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_494 = 3'h4 == total_offset_14 ? args_4 : _GEN_493; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_495 = 3'h5 == total_offset_14 ? args_5 : _GEN_494; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_496 = 3'h6 == total_offset_14 ? args_6 : _GEN_495; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_497 = total_offset_14 < 3'h7 ? _GEN_496 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_14_0 = 3'h0 < args_length_14 ? _GEN_497 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_499 = opcode_14 == 4'ha ? field_bytes_14_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_500 = opcode_14 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_381 = opcode_14 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_29 = _T_381 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_501 = opcode_14 == 4'h8 | opcode_14 == 4'hb ? parameter_2_14[7:0] : _GEN_499; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_502 = opcode_14 == 4'h8 | opcode_14 == 4'hb ? _field_tag_T_29 : _GEN_500; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_503 = 14'h0 == parameter_2_14 ? phv_data_0 : _GEN_501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_504 = 14'h1 == parameter_2_14 ? phv_data_1 : _GEN_503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_505 = 14'h2 == parameter_2_14 ? phv_data_2 : _GEN_504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_506 = 14'h3 == parameter_2_14 ? phv_data_3 : _GEN_505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_507 = 14'h4 == parameter_2_14 ? phv_data_4 : _GEN_506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_508 = 14'h5 == parameter_2_14 ? phv_data_5 : _GEN_507; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_509 = 14'h6 == parameter_2_14 ? phv_data_6 : _GEN_508; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_510 = 14'h7 == parameter_2_14 ? phv_data_7 : _GEN_509; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_511 = 14'h8 == parameter_2_14 ? phv_data_8 : _GEN_510; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_512 = 14'h9 == parameter_2_14 ? phv_data_9 : _GEN_511; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_513 = 14'ha == parameter_2_14 ? phv_data_10 : _GEN_512; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_514 = 14'hb == parameter_2_14 ? phv_data_11 : _GEN_513; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_515 = 14'hc == parameter_2_14 ? phv_data_12 : _GEN_514; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_516 = 14'hd == parameter_2_14 ? phv_data_13 : _GEN_515; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_517 = 14'he == parameter_2_14 ? phv_data_14 : _GEN_516; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_518 = 14'hf == parameter_2_14 ? phv_data_15 : _GEN_517; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_519 = 14'h10 == parameter_2_14 ? phv_data_16 : _GEN_518; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_520 = 14'h11 == parameter_2_14 ? phv_data_17 : _GEN_519; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_521 = 14'h12 == parameter_2_14 ? phv_data_18 : _GEN_520; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_522 = 14'h13 == parameter_2_14 ? phv_data_19 : _GEN_521; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_15 = vliw_15[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_15 = vliw_15[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_15 = parameter_2_15[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_15 = parameter_2_15[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_15 = {{1'd0}, args_offset_15}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_15 = _total_offset_T_15[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_526 = 3'h1 == total_offset_15 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_527 = 3'h2 == total_offset_15 ? args_2 : _GEN_526; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_528 = 3'h3 == total_offset_15 ? args_3 : _GEN_527; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_529 = 3'h4 == total_offset_15 ? args_4 : _GEN_528; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_530 = 3'h5 == total_offset_15 ? args_5 : _GEN_529; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_531 = 3'h6 == total_offset_15 ? args_6 : _GEN_530; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_532 = total_offset_15 < 3'h7 ? _GEN_531 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_15_0 = 3'h0 < args_length_15 ? _GEN_532 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_534 = opcode_15 == 4'ha ? field_bytes_15_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_535 = opcode_15 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_408 = opcode_15 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_31 = _T_408 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_536 = opcode_15 == 4'h8 | opcode_15 == 4'hb ? parameter_2_15[7:0] : _GEN_534; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_537 = opcode_15 == 4'h8 | opcode_15 == 4'hb ? _field_tag_T_31 : _GEN_535; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_538 = 14'h0 == parameter_2_15 ? phv_data_0 : _GEN_536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_539 = 14'h1 == parameter_2_15 ? phv_data_1 : _GEN_538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_540 = 14'h2 == parameter_2_15 ? phv_data_2 : _GEN_539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_541 = 14'h3 == parameter_2_15 ? phv_data_3 : _GEN_540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_542 = 14'h4 == parameter_2_15 ? phv_data_4 : _GEN_541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_543 = 14'h5 == parameter_2_15 ? phv_data_5 : _GEN_542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_544 = 14'h6 == parameter_2_15 ? phv_data_6 : _GEN_543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_545 = 14'h7 == parameter_2_15 ? phv_data_7 : _GEN_544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_546 = 14'h8 == parameter_2_15 ? phv_data_8 : _GEN_545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_547 = 14'h9 == parameter_2_15 ? phv_data_9 : _GEN_546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_548 = 14'ha == parameter_2_15 ? phv_data_10 : _GEN_547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_549 = 14'hb == parameter_2_15 ? phv_data_11 : _GEN_548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_550 = 14'hc == parameter_2_15 ? phv_data_12 : _GEN_549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_551 = 14'hd == parameter_2_15 ? phv_data_13 : _GEN_550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_552 = 14'he == parameter_2_15 ? phv_data_14 : _GEN_551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_553 = 14'hf == parameter_2_15 ? phv_data_15 : _GEN_552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_554 = 14'h10 == parameter_2_15 ? phv_data_16 : _GEN_553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_555 = 14'h11 == parameter_2_15 ? phv_data_17 : _GEN_554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_556 = 14'h12 == parameter_2_15 ? phv_data_18 : _GEN_555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_557 = 14'h13 == parameter_2_15 ? phv_data_19 : _GEN_556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_16 = vliw_16[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_16 = vliw_16[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_16 = parameter_2_16[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_16 = parameter_2_16[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_16 = {{1'd0}, args_offset_16}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_16 = _total_offset_T_16[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_561 = 3'h1 == total_offset_16 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_562 = 3'h2 == total_offset_16 ? args_2 : _GEN_561; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_563 = 3'h3 == total_offset_16 ? args_3 : _GEN_562; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_564 = 3'h4 == total_offset_16 ? args_4 : _GEN_563; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_565 = 3'h5 == total_offset_16 ? args_5 : _GEN_564; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_566 = 3'h6 == total_offset_16 ? args_6 : _GEN_565; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_567 = total_offset_16 < 3'h7 ? _GEN_566 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_16_0 = 3'h0 < args_length_16 ? _GEN_567 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_569 = opcode_16 == 4'ha ? field_bytes_16_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_570 = opcode_16 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_435 = opcode_16 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_33 = _T_435 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_571 = opcode_16 == 4'h8 | opcode_16 == 4'hb ? parameter_2_16[7:0] : _GEN_569; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_572 = opcode_16 == 4'h8 | opcode_16 == 4'hb ? _field_tag_T_33 : _GEN_570; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_573 = 14'h0 == parameter_2_16 ? phv_data_0 : _GEN_571; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_574 = 14'h1 == parameter_2_16 ? phv_data_1 : _GEN_573; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_575 = 14'h2 == parameter_2_16 ? phv_data_2 : _GEN_574; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_576 = 14'h3 == parameter_2_16 ? phv_data_3 : _GEN_575; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_577 = 14'h4 == parameter_2_16 ? phv_data_4 : _GEN_576; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_578 = 14'h5 == parameter_2_16 ? phv_data_5 : _GEN_577; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_579 = 14'h6 == parameter_2_16 ? phv_data_6 : _GEN_578; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_580 = 14'h7 == parameter_2_16 ? phv_data_7 : _GEN_579; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_581 = 14'h8 == parameter_2_16 ? phv_data_8 : _GEN_580; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_582 = 14'h9 == parameter_2_16 ? phv_data_9 : _GEN_581; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_583 = 14'ha == parameter_2_16 ? phv_data_10 : _GEN_582; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_584 = 14'hb == parameter_2_16 ? phv_data_11 : _GEN_583; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_585 = 14'hc == parameter_2_16 ? phv_data_12 : _GEN_584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_586 = 14'hd == parameter_2_16 ? phv_data_13 : _GEN_585; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_587 = 14'he == parameter_2_16 ? phv_data_14 : _GEN_586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_588 = 14'hf == parameter_2_16 ? phv_data_15 : _GEN_587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_589 = 14'h10 == parameter_2_16 ? phv_data_16 : _GEN_588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_590 = 14'h11 == parameter_2_16 ? phv_data_17 : _GEN_589; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_591 = 14'h12 == parameter_2_16 ? phv_data_18 : _GEN_590; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_592 = 14'h13 == parameter_2_16 ? phv_data_19 : _GEN_591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_17 = vliw_17[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_17 = vliw_17[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_17 = parameter_2_17[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_17 = parameter_2_17[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_17 = {{1'd0}, args_offset_17}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_17 = _total_offset_T_17[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_596 = 3'h1 == total_offset_17 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_597 = 3'h2 == total_offset_17 ? args_2 : _GEN_596; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_598 = 3'h3 == total_offset_17 ? args_3 : _GEN_597; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_599 = 3'h4 == total_offset_17 ? args_4 : _GEN_598; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_600 = 3'h5 == total_offset_17 ? args_5 : _GEN_599; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_601 = 3'h6 == total_offset_17 ? args_6 : _GEN_600; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_602 = total_offset_17 < 3'h7 ? _GEN_601 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_17_0 = 3'h0 < args_length_17 ? _GEN_602 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_604 = opcode_17 == 4'ha ? field_bytes_17_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_605 = opcode_17 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_462 = opcode_17 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_35 = _T_462 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_606 = opcode_17 == 4'h8 | opcode_17 == 4'hb ? parameter_2_17[7:0] : _GEN_604; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_607 = opcode_17 == 4'h8 | opcode_17 == 4'hb ? _field_tag_T_35 : _GEN_605; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_608 = 14'h0 == parameter_2_17 ? phv_data_0 : _GEN_606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_609 = 14'h1 == parameter_2_17 ? phv_data_1 : _GEN_608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_610 = 14'h2 == parameter_2_17 ? phv_data_2 : _GEN_609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_611 = 14'h3 == parameter_2_17 ? phv_data_3 : _GEN_610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_612 = 14'h4 == parameter_2_17 ? phv_data_4 : _GEN_611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_613 = 14'h5 == parameter_2_17 ? phv_data_5 : _GEN_612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_614 = 14'h6 == parameter_2_17 ? phv_data_6 : _GEN_613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_615 = 14'h7 == parameter_2_17 ? phv_data_7 : _GEN_614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_616 = 14'h8 == parameter_2_17 ? phv_data_8 : _GEN_615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_617 = 14'h9 == parameter_2_17 ? phv_data_9 : _GEN_616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_618 = 14'ha == parameter_2_17 ? phv_data_10 : _GEN_617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_619 = 14'hb == parameter_2_17 ? phv_data_11 : _GEN_618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_620 = 14'hc == parameter_2_17 ? phv_data_12 : _GEN_619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_621 = 14'hd == parameter_2_17 ? phv_data_13 : _GEN_620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_622 = 14'he == parameter_2_17 ? phv_data_14 : _GEN_621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_623 = 14'hf == parameter_2_17 ? phv_data_15 : _GEN_622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_624 = 14'h10 == parameter_2_17 ? phv_data_16 : _GEN_623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_625 = 14'h11 == parameter_2_17 ? phv_data_17 : _GEN_624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_626 = 14'h12 == parameter_2_17 ? phv_data_18 : _GEN_625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_627 = 14'h13 == parameter_2_17 ? phv_data_19 : _GEN_626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_18 = vliw_18[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_18 = vliw_18[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_18 = parameter_2_18[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_18 = parameter_2_18[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_18 = {{1'd0}, args_offset_18}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_18 = _total_offset_T_18[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_631 = 3'h1 == total_offset_18 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_632 = 3'h2 == total_offset_18 ? args_2 : _GEN_631; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_633 = 3'h3 == total_offset_18 ? args_3 : _GEN_632; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_634 = 3'h4 == total_offset_18 ? args_4 : _GEN_633; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_635 = 3'h5 == total_offset_18 ? args_5 : _GEN_634; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_636 = 3'h6 == total_offset_18 ? args_6 : _GEN_635; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_637 = total_offset_18 < 3'h7 ? _GEN_636 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_18_0 = 3'h0 < args_length_18 ? _GEN_637 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_639 = opcode_18 == 4'ha ? field_bytes_18_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_640 = opcode_18 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_489 = opcode_18 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_37 = _T_489 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_641 = opcode_18 == 4'h8 | opcode_18 == 4'hb ? parameter_2_18[7:0] : _GEN_639; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_642 = opcode_18 == 4'h8 | opcode_18 == 4'hb ? _field_tag_T_37 : _GEN_640; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_643 = 14'h0 == parameter_2_18 ? phv_data_0 : _GEN_641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_644 = 14'h1 == parameter_2_18 ? phv_data_1 : _GEN_643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_645 = 14'h2 == parameter_2_18 ? phv_data_2 : _GEN_644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_646 = 14'h3 == parameter_2_18 ? phv_data_3 : _GEN_645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_647 = 14'h4 == parameter_2_18 ? phv_data_4 : _GEN_646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_648 = 14'h5 == parameter_2_18 ? phv_data_5 : _GEN_647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_649 = 14'h6 == parameter_2_18 ? phv_data_6 : _GEN_648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_650 = 14'h7 == parameter_2_18 ? phv_data_7 : _GEN_649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_651 = 14'h8 == parameter_2_18 ? phv_data_8 : _GEN_650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_652 = 14'h9 == parameter_2_18 ? phv_data_9 : _GEN_651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_653 = 14'ha == parameter_2_18 ? phv_data_10 : _GEN_652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_654 = 14'hb == parameter_2_18 ? phv_data_11 : _GEN_653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_655 = 14'hc == parameter_2_18 ? phv_data_12 : _GEN_654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_656 = 14'hd == parameter_2_18 ? phv_data_13 : _GEN_655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_657 = 14'he == parameter_2_18 ? phv_data_14 : _GEN_656; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_658 = 14'hf == parameter_2_18 ? phv_data_15 : _GEN_657; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_659 = 14'h10 == parameter_2_18 ? phv_data_16 : _GEN_658; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_660 = 14'h11 == parameter_2_18 ? phv_data_17 : _GEN_659; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_661 = 14'h12 == parameter_2_18 ? phv_data_18 : _GEN_660; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_662 = 14'h13 == parameter_2_18 ? phv_data_19 : _GEN_661; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_19 = vliw_19[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] parameter_2_19 = vliw_19[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_19 = parameter_2_19[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_19 = parameter_2_19[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_19 = {{1'd0}, args_offset_19}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_19 = _total_offset_T_19[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_666 = 3'h1 == total_offset_19 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_667 = 3'h2 == total_offset_19 ? args_2 : _GEN_666; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_668 = 3'h3 == total_offset_19 ? args_3 : _GEN_667; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_669 = 3'h4 == total_offset_19 ? args_4 : _GEN_668; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_670 = 3'h5 == total_offset_19 ? args_5 : _GEN_669; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_671 = 3'h6 == total_offset_19 ? args_6 : _GEN_670; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_672 = total_offset_19 < 3'h7 ? _GEN_671 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_19_0 = 3'h0 < args_length_19 ? _GEN_672 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [7:0] _GEN_674 = opcode_19 == 4'ha ? field_bytes_19_0 : 8'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_675 = opcode_19 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_516 = opcode_19 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] _field_tag_T_39 = _T_516 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [7:0] _GEN_676 = opcode_19 == 4'h8 | opcode_19 == 4'hb ? parameter_2_19[7:0] : _GEN_674; // @[executor_pisa.scala 203:79 executor_pisa.scala 206:32]
  wire [1:0] _GEN_677 = opcode_19 == 4'h8 | opcode_19 == 4'hb ? _field_tag_T_39 : _GEN_675; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [7:0] _GEN_678 = 14'h0 == parameter_2_19 ? phv_data_0 : _GEN_676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_679 = 14'h1 == parameter_2_19 ? phv_data_1 : _GEN_678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_680 = 14'h2 == parameter_2_19 ? phv_data_2 : _GEN_679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_681 = 14'h3 == parameter_2_19 ? phv_data_3 : _GEN_680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_682 = 14'h4 == parameter_2_19 ? phv_data_4 : _GEN_681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_683 = 14'h5 == parameter_2_19 ? phv_data_5 : _GEN_682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_684 = 14'h6 == parameter_2_19 ? phv_data_6 : _GEN_683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_685 = 14'h7 == parameter_2_19 ? phv_data_7 : _GEN_684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_686 = 14'h8 == parameter_2_19 ? phv_data_8 : _GEN_685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_687 = 14'h9 == parameter_2_19 ? phv_data_9 : _GEN_686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_688 = 14'ha == parameter_2_19 ? phv_data_10 : _GEN_687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_689 = 14'hb == parameter_2_19 ? phv_data_11 : _GEN_688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_690 = 14'hc == parameter_2_19 ? phv_data_12 : _GEN_689; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_691 = 14'hd == parameter_2_19 ? phv_data_13 : _GEN_690; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_692 = 14'he == parameter_2_19 ? phv_data_14 : _GEN_691; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_693 = 14'hf == parameter_2_19 ? phv_data_15 : _GEN_692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_694 = 14'h10 == parameter_2_19 ? phv_data_16 : _GEN_693; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_695 = 14'h11 == parameter_2_19 ? phv_data_17 : _GEN_694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_696 = 14'h12 == parameter_2_19 ? phv_data_18 : _GEN_695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [7:0] _GEN_697 = 14'h13 == parameter_2_19 ? phv_data_19 : _GEN_696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_20 = vliw_20[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo = vliw_20[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_20 = field_data_lo[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_20 = field_data_lo[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_20 = {{1'd0}, args_offset_20}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_20 = _total_offset_T_20[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_701 = 3'h1 == total_offset_20 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_702 = 3'h2 == total_offset_20 ? args_2 : _GEN_701; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_703 = 3'h3 == total_offset_20 ? args_3 : _GEN_702; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_704 = 3'h4 == total_offset_20 ? args_4 : _GEN_703; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_705 = 3'h5 == total_offset_20 ? args_5 : _GEN_704; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_706 = 3'h6 == total_offset_20 ? args_6 : _GEN_705; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_707 = total_offset_20 < 3'h7 ? _GEN_706 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_20_1 = 3'h0 < args_length_20 ? _GEN_707 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_21 = args_offset_20 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_710 = 3'h1 == total_offset_21 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_711 = 3'h2 == total_offset_21 ? args_2 : _GEN_710; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_712 = 3'h3 == total_offset_21 ? args_3 : _GEN_711; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_713 = 3'h4 == total_offset_21 ? args_4 : _GEN_712; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_714 = 3'h5 == total_offset_21 ? args_5 : _GEN_713; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_715 = 3'h6 == total_offset_21 ? args_6 : _GEN_714; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_716 = total_offset_21 < 3'h7 ? _GEN_715 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_20_0 = 3'h1 < args_length_20 ? _GEN_716 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_20 = {field_bytes_20_0,field_bytes_20_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_718 = opcode_20 == 4'ha ? _field_data_T_20 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_719 = opcode_20 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_545 = opcode_20 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi = field_data_lo[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_23 = {field_data_hi,field_data_lo}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_41 = _T_545 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_720 = opcode_20 == 4'h8 | opcode_20 == 4'hb ? _field_data_T_23 : _GEN_718; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_721 = opcode_20 == 4'h8 | opcode_20 == 4'hb ? _field_tag_T_41 : _GEN_719; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _field_data_T_24 = {phv_data_20,phv_data_21}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_722 = 14'h14 == field_data_lo ? _field_data_T_24 : _GEN_720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_25 = {phv_data_22,phv_data_23}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_723 = 14'h15 == field_data_lo ? _field_data_T_25 : _GEN_722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_26 = {phv_data_24,phv_data_25}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_724 = 14'h16 == field_data_lo ? _field_data_T_26 : _GEN_723; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_27 = {phv_data_26,phv_data_27}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_725 = 14'h17 == field_data_lo ? _field_data_T_27 : _GEN_724; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_28 = {phv_data_28,phv_data_29}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_726 = 14'h18 == field_data_lo ? _field_data_T_28 : _GEN_725; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_29 = {phv_data_30,phv_data_31}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_727 = 14'h19 == field_data_lo ? _field_data_T_29 : _GEN_726; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_30 = {phv_data_32,phv_data_33}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_728 = 14'h1a == field_data_lo ? _field_data_T_30 : _GEN_727; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_31 = {phv_data_34,phv_data_35}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_729 = 14'h1b == field_data_lo ? _field_data_T_31 : _GEN_728; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_32 = {phv_data_36,phv_data_37}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_730 = 14'h1c == field_data_lo ? _field_data_T_32 : _GEN_729; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_33 = {phv_data_38,phv_data_39}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_731 = 14'h1d == field_data_lo ? _field_data_T_33 : _GEN_730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_34 = {phv_data_40,phv_data_41}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_732 = 14'h1e == field_data_lo ? _field_data_T_34 : _GEN_731; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_35 = {phv_data_42,phv_data_43}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_733 = 14'h1f == field_data_lo ? _field_data_T_35 : _GEN_732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_36 = {phv_data_44,phv_data_45}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_734 = 14'h20 == field_data_lo ? _field_data_T_36 : _GEN_733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_37 = {phv_data_46,phv_data_47}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_735 = 14'h21 == field_data_lo ? _field_data_T_37 : _GEN_734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_38 = {phv_data_48,phv_data_49}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_736 = 14'h22 == field_data_lo ? _field_data_T_38 : _GEN_735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_39 = {phv_data_50,phv_data_51}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_737 = 14'h23 == field_data_lo ? _field_data_T_39 : _GEN_736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_40 = {phv_data_52,phv_data_53}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_738 = 14'h24 == field_data_lo ? _field_data_T_40 : _GEN_737; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_41 = {phv_data_54,phv_data_55}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_739 = 14'h25 == field_data_lo ? _field_data_T_41 : _GEN_738; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_42 = {phv_data_56,phv_data_57}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_740 = 14'h26 == field_data_lo ? _field_data_T_42 : _GEN_739; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_43 = {phv_data_58,phv_data_59}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_741 = 14'h27 == field_data_lo ? _field_data_T_43 : _GEN_740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_44 = {phv_data_60,phv_data_61}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_742 = 14'h28 == field_data_lo ? _field_data_T_44 : _GEN_741; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_45 = {phv_data_62,phv_data_63}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_743 = 14'h29 == field_data_lo ? _field_data_T_45 : _GEN_742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_46 = {phv_data_64,phv_data_65}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_744 = 14'h2a == field_data_lo ? _field_data_T_46 : _GEN_743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_47 = {phv_data_66,phv_data_67}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_745 = 14'h2b == field_data_lo ? _field_data_T_47 : _GEN_744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_48 = {phv_data_68,phv_data_69}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_746 = 14'h2c == field_data_lo ? _field_data_T_48 : _GEN_745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_49 = {phv_data_70,phv_data_71}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_747 = 14'h2d == field_data_lo ? _field_data_T_49 : _GEN_746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_50 = {phv_data_72,phv_data_73}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_748 = 14'h2e == field_data_lo ? _field_data_T_50 : _GEN_747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_51 = {phv_data_74,phv_data_75}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_749 = 14'h2f == field_data_lo ? _field_data_T_51 : _GEN_748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_52 = {phv_data_76,phv_data_77}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_750 = 14'h30 == field_data_lo ? _field_data_T_52 : _GEN_749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _field_data_T_53 = {phv_data_78,phv_data_79}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_751 = 14'h31 == field_data_lo ? _field_data_T_53 : _GEN_750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_21 = vliw_21[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_1 = vliw_21[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_21 = field_data_lo_1[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_21 = field_data_lo_1[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_22 = {{1'd0}, args_offset_21}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_22 = _total_offset_T_22[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_755 = 3'h1 == total_offset_22 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_756 = 3'h2 == total_offset_22 ? args_2 : _GEN_755; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_757 = 3'h3 == total_offset_22 ? args_3 : _GEN_756; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_758 = 3'h4 == total_offset_22 ? args_4 : _GEN_757; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_759 = 3'h5 == total_offset_22 ? args_5 : _GEN_758; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_760 = 3'h6 == total_offset_22 ? args_6 : _GEN_759; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_761 = total_offset_22 < 3'h7 ? _GEN_760 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_21_1 = 3'h0 < args_length_21 ? _GEN_761 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_23 = args_offset_21 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_764 = 3'h1 == total_offset_23 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_765 = 3'h2 == total_offset_23 ? args_2 : _GEN_764; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_766 = 3'h3 == total_offset_23 ? args_3 : _GEN_765; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_767 = 3'h4 == total_offset_23 ? args_4 : _GEN_766; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_768 = 3'h5 == total_offset_23 ? args_5 : _GEN_767; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_769 = 3'h6 == total_offset_23 ? args_6 : _GEN_768; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_770 = total_offset_23 < 3'h7 ? _GEN_769 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_21_0 = 3'h1 < args_length_21 ? _GEN_770 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_54 = {field_bytes_21_0,field_bytes_21_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_772 = opcode_21 == 4'ha ? _field_data_T_54 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_773 = opcode_21 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_584 = opcode_21 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_1 = field_data_lo_1[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_57 = {field_data_hi_1,field_data_lo_1}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_43 = _T_584 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_774 = opcode_21 == 4'h8 | opcode_21 == 4'hb ? _field_data_T_57 : _GEN_772; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_775 = opcode_21 == 4'h8 | opcode_21 == 4'hb ? _field_tag_T_43 : _GEN_773; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_776 = 14'h14 == field_data_lo_1 ? _field_data_T_24 : _GEN_774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_777 = 14'h15 == field_data_lo_1 ? _field_data_T_25 : _GEN_776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_778 = 14'h16 == field_data_lo_1 ? _field_data_T_26 : _GEN_777; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_779 = 14'h17 == field_data_lo_1 ? _field_data_T_27 : _GEN_778; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_780 = 14'h18 == field_data_lo_1 ? _field_data_T_28 : _GEN_779; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_781 = 14'h19 == field_data_lo_1 ? _field_data_T_29 : _GEN_780; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_782 = 14'h1a == field_data_lo_1 ? _field_data_T_30 : _GEN_781; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_783 = 14'h1b == field_data_lo_1 ? _field_data_T_31 : _GEN_782; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_784 = 14'h1c == field_data_lo_1 ? _field_data_T_32 : _GEN_783; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_785 = 14'h1d == field_data_lo_1 ? _field_data_T_33 : _GEN_784; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_786 = 14'h1e == field_data_lo_1 ? _field_data_T_34 : _GEN_785; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_787 = 14'h1f == field_data_lo_1 ? _field_data_T_35 : _GEN_786; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_788 = 14'h20 == field_data_lo_1 ? _field_data_T_36 : _GEN_787; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_789 = 14'h21 == field_data_lo_1 ? _field_data_T_37 : _GEN_788; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_790 = 14'h22 == field_data_lo_1 ? _field_data_T_38 : _GEN_789; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_791 = 14'h23 == field_data_lo_1 ? _field_data_T_39 : _GEN_790; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_792 = 14'h24 == field_data_lo_1 ? _field_data_T_40 : _GEN_791; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_793 = 14'h25 == field_data_lo_1 ? _field_data_T_41 : _GEN_792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_794 = 14'h26 == field_data_lo_1 ? _field_data_T_42 : _GEN_793; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_795 = 14'h27 == field_data_lo_1 ? _field_data_T_43 : _GEN_794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_796 = 14'h28 == field_data_lo_1 ? _field_data_T_44 : _GEN_795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_797 = 14'h29 == field_data_lo_1 ? _field_data_T_45 : _GEN_796; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_798 = 14'h2a == field_data_lo_1 ? _field_data_T_46 : _GEN_797; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_799 = 14'h2b == field_data_lo_1 ? _field_data_T_47 : _GEN_798; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_800 = 14'h2c == field_data_lo_1 ? _field_data_T_48 : _GEN_799; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_801 = 14'h2d == field_data_lo_1 ? _field_data_T_49 : _GEN_800; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_802 = 14'h2e == field_data_lo_1 ? _field_data_T_50 : _GEN_801; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_803 = 14'h2f == field_data_lo_1 ? _field_data_T_51 : _GEN_802; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_804 = 14'h30 == field_data_lo_1 ? _field_data_T_52 : _GEN_803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_805 = 14'h31 == field_data_lo_1 ? _field_data_T_53 : _GEN_804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_22 = vliw_22[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_2 = vliw_22[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_22 = field_data_lo_2[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_22 = field_data_lo_2[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_24 = {{1'd0}, args_offset_22}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_24 = _total_offset_T_24[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_809 = 3'h1 == total_offset_24 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_810 = 3'h2 == total_offset_24 ? args_2 : _GEN_809; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_811 = 3'h3 == total_offset_24 ? args_3 : _GEN_810; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_812 = 3'h4 == total_offset_24 ? args_4 : _GEN_811; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_813 = 3'h5 == total_offset_24 ? args_5 : _GEN_812; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_814 = 3'h6 == total_offset_24 ? args_6 : _GEN_813; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_815 = total_offset_24 < 3'h7 ? _GEN_814 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_22_1 = 3'h0 < args_length_22 ? _GEN_815 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_25 = args_offset_22 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_818 = 3'h1 == total_offset_25 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_819 = 3'h2 == total_offset_25 ? args_2 : _GEN_818; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_820 = 3'h3 == total_offset_25 ? args_3 : _GEN_819; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_821 = 3'h4 == total_offset_25 ? args_4 : _GEN_820; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_822 = 3'h5 == total_offset_25 ? args_5 : _GEN_821; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_823 = 3'h6 == total_offset_25 ? args_6 : _GEN_822; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_824 = total_offset_25 < 3'h7 ? _GEN_823 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_22_0 = 3'h1 < args_length_22 ? _GEN_824 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_88 = {field_bytes_22_0,field_bytes_22_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_826 = opcode_22 == 4'ha ? _field_data_T_88 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_827 = opcode_22 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_623 = opcode_22 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_2 = field_data_lo_2[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_91 = {field_data_hi_2,field_data_lo_2}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_45 = _T_623 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_828 = opcode_22 == 4'h8 | opcode_22 == 4'hb ? _field_data_T_91 : _GEN_826; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_829 = opcode_22 == 4'h8 | opcode_22 == 4'hb ? _field_tag_T_45 : _GEN_827; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_830 = 14'h14 == field_data_lo_2 ? _field_data_T_24 : _GEN_828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_831 = 14'h15 == field_data_lo_2 ? _field_data_T_25 : _GEN_830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_832 = 14'h16 == field_data_lo_2 ? _field_data_T_26 : _GEN_831; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_833 = 14'h17 == field_data_lo_2 ? _field_data_T_27 : _GEN_832; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_834 = 14'h18 == field_data_lo_2 ? _field_data_T_28 : _GEN_833; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_835 = 14'h19 == field_data_lo_2 ? _field_data_T_29 : _GEN_834; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_836 = 14'h1a == field_data_lo_2 ? _field_data_T_30 : _GEN_835; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_837 = 14'h1b == field_data_lo_2 ? _field_data_T_31 : _GEN_836; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_838 = 14'h1c == field_data_lo_2 ? _field_data_T_32 : _GEN_837; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_839 = 14'h1d == field_data_lo_2 ? _field_data_T_33 : _GEN_838; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_840 = 14'h1e == field_data_lo_2 ? _field_data_T_34 : _GEN_839; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_841 = 14'h1f == field_data_lo_2 ? _field_data_T_35 : _GEN_840; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_842 = 14'h20 == field_data_lo_2 ? _field_data_T_36 : _GEN_841; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_843 = 14'h21 == field_data_lo_2 ? _field_data_T_37 : _GEN_842; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_844 = 14'h22 == field_data_lo_2 ? _field_data_T_38 : _GEN_843; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_845 = 14'h23 == field_data_lo_2 ? _field_data_T_39 : _GEN_844; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_846 = 14'h24 == field_data_lo_2 ? _field_data_T_40 : _GEN_845; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_847 = 14'h25 == field_data_lo_2 ? _field_data_T_41 : _GEN_846; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_848 = 14'h26 == field_data_lo_2 ? _field_data_T_42 : _GEN_847; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_849 = 14'h27 == field_data_lo_2 ? _field_data_T_43 : _GEN_848; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_850 = 14'h28 == field_data_lo_2 ? _field_data_T_44 : _GEN_849; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_851 = 14'h29 == field_data_lo_2 ? _field_data_T_45 : _GEN_850; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_852 = 14'h2a == field_data_lo_2 ? _field_data_T_46 : _GEN_851; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_853 = 14'h2b == field_data_lo_2 ? _field_data_T_47 : _GEN_852; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_854 = 14'h2c == field_data_lo_2 ? _field_data_T_48 : _GEN_853; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_855 = 14'h2d == field_data_lo_2 ? _field_data_T_49 : _GEN_854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_856 = 14'h2e == field_data_lo_2 ? _field_data_T_50 : _GEN_855; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_857 = 14'h2f == field_data_lo_2 ? _field_data_T_51 : _GEN_856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_858 = 14'h30 == field_data_lo_2 ? _field_data_T_52 : _GEN_857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_859 = 14'h31 == field_data_lo_2 ? _field_data_T_53 : _GEN_858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_23 = vliw_23[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_3 = vliw_23[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_23 = field_data_lo_3[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_23 = field_data_lo_3[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_26 = {{1'd0}, args_offset_23}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_26 = _total_offset_T_26[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_863 = 3'h1 == total_offset_26 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_864 = 3'h2 == total_offset_26 ? args_2 : _GEN_863; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_865 = 3'h3 == total_offset_26 ? args_3 : _GEN_864; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_866 = 3'h4 == total_offset_26 ? args_4 : _GEN_865; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_867 = 3'h5 == total_offset_26 ? args_5 : _GEN_866; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_868 = 3'h6 == total_offset_26 ? args_6 : _GEN_867; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_869 = total_offset_26 < 3'h7 ? _GEN_868 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_23_1 = 3'h0 < args_length_23 ? _GEN_869 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_27 = args_offset_23 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_872 = 3'h1 == total_offset_27 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_873 = 3'h2 == total_offset_27 ? args_2 : _GEN_872; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_874 = 3'h3 == total_offset_27 ? args_3 : _GEN_873; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_875 = 3'h4 == total_offset_27 ? args_4 : _GEN_874; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_876 = 3'h5 == total_offset_27 ? args_5 : _GEN_875; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_877 = 3'h6 == total_offset_27 ? args_6 : _GEN_876; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_878 = total_offset_27 < 3'h7 ? _GEN_877 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_23_0 = 3'h1 < args_length_23 ? _GEN_878 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_122 = {field_bytes_23_0,field_bytes_23_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_880 = opcode_23 == 4'ha ? _field_data_T_122 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_881 = opcode_23 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_662 = opcode_23 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_3 = field_data_lo_3[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_125 = {field_data_hi_3,field_data_lo_3}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_47 = _T_662 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_882 = opcode_23 == 4'h8 | opcode_23 == 4'hb ? _field_data_T_125 : _GEN_880; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_883 = opcode_23 == 4'h8 | opcode_23 == 4'hb ? _field_tag_T_47 : _GEN_881; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_884 = 14'h14 == field_data_lo_3 ? _field_data_T_24 : _GEN_882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_885 = 14'h15 == field_data_lo_3 ? _field_data_T_25 : _GEN_884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_886 = 14'h16 == field_data_lo_3 ? _field_data_T_26 : _GEN_885; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_887 = 14'h17 == field_data_lo_3 ? _field_data_T_27 : _GEN_886; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_888 = 14'h18 == field_data_lo_3 ? _field_data_T_28 : _GEN_887; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_889 = 14'h19 == field_data_lo_3 ? _field_data_T_29 : _GEN_888; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_890 = 14'h1a == field_data_lo_3 ? _field_data_T_30 : _GEN_889; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_891 = 14'h1b == field_data_lo_3 ? _field_data_T_31 : _GEN_890; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_892 = 14'h1c == field_data_lo_3 ? _field_data_T_32 : _GEN_891; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_893 = 14'h1d == field_data_lo_3 ? _field_data_T_33 : _GEN_892; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_894 = 14'h1e == field_data_lo_3 ? _field_data_T_34 : _GEN_893; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_895 = 14'h1f == field_data_lo_3 ? _field_data_T_35 : _GEN_894; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_896 = 14'h20 == field_data_lo_3 ? _field_data_T_36 : _GEN_895; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_897 = 14'h21 == field_data_lo_3 ? _field_data_T_37 : _GEN_896; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_898 = 14'h22 == field_data_lo_3 ? _field_data_T_38 : _GEN_897; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_899 = 14'h23 == field_data_lo_3 ? _field_data_T_39 : _GEN_898; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_900 = 14'h24 == field_data_lo_3 ? _field_data_T_40 : _GEN_899; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_901 = 14'h25 == field_data_lo_3 ? _field_data_T_41 : _GEN_900; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_902 = 14'h26 == field_data_lo_3 ? _field_data_T_42 : _GEN_901; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_903 = 14'h27 == field_data_lo_3 ? _field_data_T_43 : _GEN_902; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_904 = 14'h28 == field_data_lo_3 ? _field_data_T_44 : _GEN_903; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_905 = 14'h29 == field_data_lo_3 ? _field_data_T_45 : _GEN_904; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_906 = 14'h2a == field_data_lo_3 ? _field_data_T_46 : _GEN_905; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_907 = 14'h2b == field_data_lo_3 ? _field_data_T_47 : _GEN_906; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_908 = 14'h2c == field_data_lo_3 ? _field_data_T_48 : _GEN_907; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_909 = 14'h2d == field_data_lo_3 ? _field_data_T_49 : _GEN_908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_910 = 14'h2e == field_data_lo_3 ? _field_data_T_50 : _GEN_909; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_911 = 14'h2f == field_data_lo_3 ? _field_data_T_51 : _GEN_910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_912 = 14'h30 == field_data_lo_3 ? _field_data_T_52 : _GEN_911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_913 = 14'h31 == field_data_lo_3 ? _field_data_T_53 : _GEN_912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_24 = vliw_24[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_4 = vliw_24[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_24 = field_data_lo_4[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_24 = field_data_lo_4[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_28 = {{1'd0}, args_offset_24}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_28 = _total_offset_T_28[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_917 = 3'h1 == total_offset_28 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_918 = 3'h2 == total_offset_28 ? args_2 : _GEN_917; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_919 = 3'h3 == total_offset_28 ? args_3 : _GEN_918; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_920 = 3'h4 == total_offset_28 ? args_4 : _GEN_919; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_921 = 3'h5 == total_offset_28 ? args_5 : _GEN_920; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_922 = 3'h6 == total_offset_28 ? args_6 : _GEN_921; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_923 = total_offset_28 < 3'h7 ? _GEN_922 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_24_1 = 3'h0 < args_length_24 ? _GEN_923 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_29 = args_offset_24 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_926 = 3'h1 == total_offset_29 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_927 = 3'h2 == total_offset_29 ? args_2 : _GEN_926; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_928 = 3'h3 == total_offset_29 ? args_3 : _GEN_927; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_929 = 3'h4 == total_offset_29 ? args_4 : _GEN_928; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_930 = 3'h5 == total_offset_29 ? args_5 : _GEN_929; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_931 = 3'h6 == total_offset_29 ? args_6 : _GEN_930; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_932 = total_offset_29 < 3'h7 ? _GEN_931 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_24_0 = 3'h1 < args_length_24 ? _GEN_932 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_156 = {field_bytes_24_0,field_bytes_24_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_934 = opcode_24 == 4'ha ? _field_data_T_156 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_935 = opcode_24 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_701 = opcode_24 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_4 = field_data_lo_4[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_159 = {field_data_hi_4,field_data_lo_4}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_49 = _T_701 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_936 = opcode_24 == 4'h8 | opcode_24 == 4'hb ? _field_data_T_159 : _GEN_934; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_937 = opcode_24 == 4'h8 | opcode_24 == 4'hb ? _field_tag_T_49 : _GEN_935; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_938 = 14'h14 == field_data_lo_4 ? _field_data_T_24 : _GEN_936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_939 = 14'h15 == field_data_lo_4 ? _field_data_T_25 : _GEN_938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_940 = 14'h16 == field_data_lo_4 ? _field_data_T_26 : _GEN_939; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_941 = 14'h17 == field_data_lo_4 ? _field_data_T_27 : _GEN_940; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_942 = 14'h18 == field_data_lo_4 ? _field_data_T_28 : _GEN_941; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_943 = 14'h19 == field_data_lo_4 ? _field_data_T_29 : _GEN_942; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_944 = 14'h1a == field_data_lo_4 ? _field_data_T_30 : _GEN_943; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_945 = 14'h1b == field_data_lo_4 ? _field_data_T_31 : _GEN_944; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_946 = 14'h1c == field_data_lo_4 ? _field_data_T_32 : _GEN_945; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_947 = 14'h1d == field_data_lo_4 ? _field_data_T_33 : _GEN_946; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_948 = 14'h1e == field_data_lo_4 ? _field_data_T_34 : _GEN_947; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_949 = 14'h1f == field_data_lo_4 ? _field_data_T_35 : _GEN_948; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_950 = 14'h20 == field_data_lo_4 ? _field_data_T_36 : _GEN_949; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_951 = 14'h21 == field_data_lo_4 ? _field_data_T_37 : _GEN_950; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_952 = 14'h22 == field_data_lo_4 ? _field_data_T_38 : _GEN_951; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_953 = 14'h23 == field_data_lo_4 ? _field_data_T_39 : _GEN_952; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_954 = 14'h24 == field_data_lo_4 ? _field_data_T_40 : _GEN_953; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_955 = 14'h25 == field_data_lo_4 ? _field_data_T_41 : _GEN_954; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_956 = 14'h26 == field_data_lo_4 ? _field_data_T_42 : _GEN_955; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_957 = 14'h27 == field_data_lo_4 ? _field_data_T_43 : _GEN_956; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_958 = 14'h28 == field_data_lo_4 ? _field_data_T_44 : _GEN_957; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_959 = 14'h29 == field_data_lo_4 ? _field_data_T_45 : _GEN_958; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_960 = 14'h2a == field_data_lo_4 ? _field_data_T_46 : _GEN_959; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_961 = 14'h2b == field_data_lo_4 ? _field_data_T_47 : _GEN_960; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_962 = 14'h2c == field_data_lo_4 ? _field_data_T_48 : _GEN_961; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_963 = 14'h2d == field_data_lo_4 ? _field_data_T_49 : _GEN_962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_964 = 14'h2e == field_data_lo_4 ? _field_data_T_50 : _GEN_963; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_965 = 14'h2f == field_data_lo_4 ? _field_data_T_51 : _GEN_964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_966 = 14'h30 == field_data_lo_4 ? _field_data_T_52 : _GEN_965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_967 = 14'h31 == field_data_lo_4 ? _field_data_T_53 : _GEN_966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_25 = vliw_25[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_5 = vliw_25[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_25 = field_data_lo_5[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_25 = field_data_lo_5[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_30 = {{1'd0}, args_offset_25}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_30 = _total_offset_T_30[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_971 = 3'h1 == total_offset_30 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_972 = 3'h2 == total_offset_30 ? args_2 : _GEN_971; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_973 = 3'h3 == total_offset_30 ? args_3 : _GEN_972; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_974 = 3'h4 == total_offset_30 ? args_4 : _GEN_973; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_975 = 3'h5 == total_offset_30 ? args_5 : _GEN_974; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_976 = 3'h6 == total_offset_30 ? args_6 : _GEN_975; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_977 = total_offset_30 < 3'h7 ? _GEN_976 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_25_1 = 3'h0 < args_length_25 ? _GEN_977 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_31 = args_offset_25 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_980 = 3'h1 == total_offset_31 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_981 = 3'h2 == total_offset_31 ? args_2 : _GEN_980; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_982 = 3'h3 == total_offset_31 ? args_3 : _GEN_981; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_983 = 3'h4 == total_offset_31 ? args_4 : _GEN_982; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_984 = 3'h5 == total_offset_31 ? args_5 : _GEN_983; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_985 = 3'h6 == total_offset_31 ? args_6 : _GEN_984; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_986 = total_offset_31 < 3'h7 ? _GEN_985 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_25_0 = 3'h1 < args_length_25 ? _GEN_986 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_190 = {field_bytes_25_0,field_bytes_25_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_988 = opcode_25 == 4'ha ? _field_data_T_190 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_989 = opcode_25 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_740 = opcode_25 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_5 = field_data_lo_5[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_193 = {field_data_hi_5,field_data_lo_5}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_51 = _T_740 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_990 = opcode_25 == 4'h8 | opcode_25 == 4'hb ? _field_data_T_193 : _GEN_988; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_991 = opcode_25 == 4'h8 | opcode_25 == 4'hb ? _field_tag_T_51 : _GEN_989; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_992 = 14'h14 == field_data_lo_5 ? _field_data_T_24 : _GEN_990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_993 = 14'h15 == field_data_lo_5 ? _field_data_T_25 : _GEN_992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_994 = 14'h16 == field_data_lo_5 ? _field_data_T_26 : _GEN_993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_995 = 14'h17 == field_data_lo_5 ? _field_data_T_27 : _GEN_994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_996 = 14'h18 == field_data_lo_5 ? _field_data_T_28 : _GEN_995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_997 = 14'h19 == field_data_lo_5 ? _field_data_T_29 : _GEN_996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_998 = 14'h1a == field_data_lo_5 ? _field_data_T_30 : _GEN_997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_999 = 14'h1b == field_data_lo_5 ? _field_data_T_31 : _GEN_998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1000 = 14'h1c == field_data_lo_5 ? _field_data_T_32 : _GEN_999; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1001 = 14'h1d == field_data_lo_5 ? _field_data_T_33 : _GEN_1000; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1002 = 14'h1e == field_data_lo_5 ? _field_data_T_34 : _GEN_1001; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1003 = 14'h1f == field_data_lo_5 ? _field_data_T_35 : _GEN_1002; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1004 = 14'h20 == field_data_lo_5 ? _field_data_T_36 : _GEN_1003; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1005 = 14'h21 == field_data_lo_5 ? _field_data_T_37 : _GEN_1004; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1006 = 14'h22 == field_data_lo_5 ? _field_data_T_38 : _GEN_1005; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1007 = 14'h23 == field_data_lo_5 ? _field_data_T_39 : _GEN_1006; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1008 = 14'h24 == field_data_lo_5 ? _field_data_T_40 : _GEN_1007; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1009 = 14'h25 == field_data_lo_5 ? _field_data_T_41 : _GEN_1008; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1010 = 14'h26 == field_data_lo_5 ? _field_data_T_42 : _GEN_1009; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1011 = 14'h27 == field_data_lo_5 ? _field_data_T_43 : _GEN_1010; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1012 = 14'h28 == field_data_lo_5 ? _field_data_T_44 : _GEN_1011; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1013 = 14'h29 == field_data_lo_5 ? _field_data_T_45 : _GEN_1012; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1014 = 14'h2a == field_data_lo_5 ? _field_data_T_46 : _GEN_1013; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1015 = 14'h2b == field_data_lo_5 ? _field_data_T_47 : _GEN_1014; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1016 = 14'h2c == field_data_lo_5 ? _field_data_T_48 : _GEN_1015; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1017 = 14'h2d == field_data_lo_5 ? _field_data_T_49 : _GEN_1016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1018 = 14'h2e == field_data_lo_5 ? _field_data_T_50 : _GEN_1017; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1019 = 14'h2f == field_data_lo_5 ? _field_data_T_51 : _GEN_1018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1020 = 14'h30 == field_data_lo_5 ? _field_data_T_52 : _GEN_1019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1021 = 14'h31 == field_data_lo_5 ? _field_data_T_53 : _GEN_1020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_26 = vliw_26[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_6 = vliw_26[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_26 = field_data_lo_6[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_26 = field_data_lo_6[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_32 = {{1'd0}, args_offset_26}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_32 = _total_offset_T_32[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1025 = 3'h1 == total_offset_32 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1026 = 3'h2 == total_offset_32 ? args_2 : _GEN_1025; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1027 = 3'h3 == total_offset_32 ? args_3 : _GEN_1026; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1028 = 3'h4 == total_offset_32 ? args_4 : _GEN_1027; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1029 = 3'h5 == total_offset_32 ? args_5 : _GEN_1028; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1030 = 3'h6 == total_offset_32 ? args_6 : _GEN_1029; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1031 = total_offset_32 < 3'h7 ? _GEN_1030 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_26_1 = 3'h0 < args_length_26 ? _GEN_1031 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_33 = args_offset_26 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1034 = 3'h1 == total_offset_33 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1035 = 3'h2 == total_offset_33 ? args_2 : _GEN_1034; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1036 = 3'h3 == total_offset_33 ? args_3 : _GEN_1035; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1037 = 3'h4 == total_offset_33 ? args_4 : _GEN_1036; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1038 = 3'h5 == total_offset_33 ? args_5 : _GEN_1037; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1039 = 3'h6 == total_offset_33 ? args_6 : _GEN_1038; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1040 = total_offset_33 < 3'h7 ? _GEN_1039 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_26_0 = 3'h1 < args_length_26 ? _GEN_1040 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_224 = {field_bytes_26_0,field_bytes_26_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1042 = opcode_26 == 4'ha ? _field_data_T_224 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1043 = opcode_26 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_779 = opcode_26 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_6 = field_data_lo_6[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_227 = {field_data_hi_6,field_data_lo_6}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_53 = _T_779 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1044 = opcode_26 == 4'h8 | opcode_26 == 4'hb ? _field_data_T_227 : _GEN_1042; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1045 = opcode_26 == 4'h8 | opcode_26 == 4'hb ? _field_tag_T_53 : _GEN_1043; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1046 = 14'h14 == field_data_lo_6 ? _field_data_T_24 : _GEN_1044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1047 = 14'h15 == field_data_lo_6 ? _field_data_T_25 : _GEN_1046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1048 = 14'h16 == field_data_lo_6 ? _field_data_T_26 : _GEN_1047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1049 = 14'h17 == field_data_lo_6 ? _field_data_T_27 : _GEN_1048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1050 = 14'h18 == field_data_lo_6 ? _field_data_T_28 : _GEN_1049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1051 = 14'h19 == field_data_lo_6 ? _field_data_T_29 : _GEN_1050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1052 = 14'h1a == field_data_lo_6 ? _field_data_T_30 : _GEN_1051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1053 = 14'h1b == field_data_lo_6 ? _field_data_T_31 : _GEN_1052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1054 = 14'h1c == field_data_lo_6 ? _field_data_T_32 : _GEN_1053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1055 = 14'h1d == field_data_lo_6 ? _field_data_T_33 : _GEN_1054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1056 = 14'h1e == field_data_lo_6 ? _field_data_T_34 : _GEN_1055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1057 = 14'h1f == field_data_lo_6 ? _field_data_T_35 : _GEN_1056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1058 = 14'h20 == field_data_lo_6 ? _field_data_T_36 : _GEN_1057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1059 = 14'h21 == field_data_lo_6 ? _field_data_T_37 : _GEN_1058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1060 = 14'h22 == field_data_lo_6 ? _field_data_T_38 : _GEN_1059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1061 = 14'h23 == field_data_lo_6 ? _field_data_T_39 : _GEN_1060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1062 = 14'h24 == field_data_lo_6 ? _field_data_T_40 : _GEN_1061; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1063 = 14'h25 == field_data_lo_6 ? _field_data_T_41 : _GEN_1062; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1064 = 14'h26 == field_data_lo_6 ? _field_data_T_42 : _GEN_1063; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1065 = 14'h27 == field_data_lo_6 ? _field_data_T_43 : _GEN_1064; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1066 = 14'h28 == field_data_lo_6 ? _field_data_T_44 : _GEN_1065; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1067 = 14'h29 == field_data_lo_6 ? _field_data_T_45 : _GEN_1066; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1068 = 14'h2a == field_data_lo_6 ? _field_data_T_46 : _GEN_1067; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1069 = 14'h2b == field_data_lo_6 ? _field_data_T_47 : _GEN_1068; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1070 = 14'h2c == field_data_lo_6 ? _field_data_T_48 : _GEN_1069; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1071 = 14'h2d == field_data_lo_6 ? _field_data_T_49 : _GEN_1070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1072 = 14'h2e == field_data_lo_6 ? _field_data_T_50 : _GEN_1071; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1073 = 14'h2f == field_data_lo_6 ? _field_data_T_51 : _GEN_1072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1074 = 14'h30 == field_data_lo_6 ? _field_data_T_52 : _GEN_1073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1075 = 14'h31 == field_data_lo_6 ? _field_data_T_53 : _GEN_1074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_27 = vliw_27[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_7 = vliw_27[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_27 = field_data_lo_7[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_27 = field_data_lo_7[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_34 = {{1'd0}, args_offset_27}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_34 = _total_offset_T_34[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1079 = 3'h1 == total_offset_34 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1080 = 3'h2 == total_offset_34 ? args_2 : _GEN_1079; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1081 = 3'h3 == total_offset_34 ? args_3 : _GEN_1080; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1082 = 3'h4 == total_offset_34 ? args_4 : _GEN_1081; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1083 = 3'h5 == total_offset_34 ? args_5 : _GEN_1082; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1084 = 3'h6 == total_offset_34 ? args_6 : _GEN_1083; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1085 = total_offset_34 < 3'h7 ? _GEN_1084 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_27_1 = 3'h0 < args_length_27 ? _GEN_1085 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_35 = args_offset_27 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1088 = 3'h1 == total_offset_35 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1089 = 3'h2 == total_offset_35 ? args_2 : _GEN_1088; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1090 = 3'h3 == total_offset_35 ? args_3 : _GEN_1089; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1091 = 3'h4 == total_offset_35 ? args_4 : _GEN_1090; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1092 = 3'h5 == total_offset_35 ? args_5 : _GEN_1091; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1093 = 3'h6 == total_offset_35 ? args_6 : _GEN_1092; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1094 = total_offset_35 < 3'h7 ? _GEN_1093 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_27_0 = 3'h1 < args_length_27 ? _GEN_1094 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_258 = {field_bytes_27_0,field_bytes_27_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1096 = opcode_27 == 4'ha ? _field_data_T_258 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1097 = opcode_27 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_818 = opcode_27 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_7 = field_data_lo_7[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_261 = {field_data_hi_7,field_data_lo_7}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_55 = _T_818 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1098 = opcode_27 == 4'h8 | opcode_27 == 4'hb ? _field_data_T_261 : _GEN_1096; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1099 = opcode_27 == 4'h8 | opcode_27 == 4'hb ? _field_tag_T_55 : _GEN_1097; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1100 = 14'h14 == field_data_lo_7 ? _field_data_T_24 : _GEN_1098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1101 = 14'h15 == field_data_lo_7 ? _field_data_T_25 : _GEN_1100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1102 = 14'h16 == field_data_lo_7 ? _field_data_T_26 : _GEN_1101; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1103 = 14'h17 == field_data_lo_7 ? _field_data_T_27 : _GEN_1102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1104 = 14'h18 == field_data_lo_7 ? _field_data_T_28 : _GEN_1103; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1105 = 14'h19 == field_data_lo_7 ? _field_data_T_29 : _GEN_1104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1106 = 14'h1a == field_data_lo_7 ? _field_data_T_30 : _GEN_1105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1107 = 14'h1b == field_data_lo_7 ? _field_data_T_31 : _GEN_1106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1108 = 14'h1c == field_data_lo_7 ? _field_data_T_32 : _GEN_1107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1109 = 14'h1d == field_data_lo_7 ? _field_data_T_33 : _GEN_1108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1110 = 14'h1e == field_data_lo_7 ? _field_data_T_34 : _GEN_1109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1111 = 14'h1f == field_data_lo_7 ? _field_data_T_35 : _GEN_1110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1112 = 14'h20 == field_data_lo_7 ? _field_data_T_36 : _GEN_1111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1113 = 14'h21 == field_data_lo_7 ? _field_data_T_37 : _GEN_1112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1114 = 14'h22 == field_data_lo_7 ? _field_data_T_38 : _GEN_1113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1115 = 14'h23 == field_data_lo_7 ? _field_data_T_39 : _GEN_1114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1116 = 14'h24 == field_data_lo_7 ? _field_data_T_40 : _GEN_1115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1117 = 14'h25 == field_data_lo_7 ? _field_data_T_41 : _GEN_1116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1118 = 14'h26 == field_data_lo_7 ? _field_data_T_42 : _GEN_1117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1119 = 14'h27 == field_data_lo_7 ? _field_data_T_43 : _GEN_1118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1120 = 14'h28 == field_data_lo_7 ? _field_data_T_44 : _GEN_1119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1121 = 14'h29 == field_data_lo_7 ? _field_data_T_45 : _GEN_1120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1122 = 14'h2a == field_data_lo_7 ? _field_data_T_46 : _GEN_1121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1123 = 14'h2b == field_data_lo_7 ? _field_data_T_47 : _GEN_1122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1124 = 14'h2c == field_data_lo_7 ? _field_data_T_48 : _GEN_1123; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1125 = 14'h2d == field_data_lo_7 ? _field_data_T_49 : _GEN_1124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1126 = 14'h2e == field_data_lo_7 ? _field_data_T_50 : _GEN_1125; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1127 = 14'h2f == field_data_lo_7 ? _field_data_T_51 : _GEN_1126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1128 = 14'h30 == field_data_lo_7 ? _field_data_T_52 : _GEN_1127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1129 = 14'h31 == field_data_lo_7 ? _field_data_T_53 : _GEN_1128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_28 = vliw_28[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_8 = vliw_28[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_28 = field_data_lo_8[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_28 = field_data_lo_8[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_36 = {{1'd0}, args_offset_28}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_36 = _total_offset_T_36[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1133 = 3'h1 == total_offset_36 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1134 = 3'h2 == total_offset_36 ? args_2 : _GEN_1133; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1135 = 3'h3 == total_offset_36 ? args_3 : _GEN_1134; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1136 = 3'h4 == total_offset_36 ? args_4 : _GEN_1135; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1137 = 3'h5 == total_offset_36 ? args_5 : _GEN_1136; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1138 = 3'h6 == total_offset_36 ? args_6 : _GEN_1137; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1139 = total_offset_36 < 3'h7 ? _GEN_1138 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_28_1 = 3'h0 < args_length_28 ? _GEN_1139 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_37 = args_offset_28 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1142 = 3'h1 == total_offset_37 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1143 = 3'h2 == total_offset_37 ? args_2 : _GEN_1142; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1144 = 3'h3 == total_offset_37 ? args_3 : _GEN_1143; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1145 = 3'h4 == total_offset_37 ? args_4 : _GEN_1144; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1146 = 3'h5 == total_offset_37 ? args_5 : _GEN_1145; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1147 = 3'h6 == total_offset_37 ? args_6 : _GEN_1146; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1148 = total_offset_37 < 3'h7 ? _GEN_1147 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_28_0 = 3'h1 < args_length_28 ? _GEN_1148 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_292 = {field_bytes_28_0,field_bytes_28_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1150 = opcode_28 == 4'ha ? _field_data_T_292 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1151 = opcode_28 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_857 = opcode_28 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_8 = field_data_lo_8[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_295 = {field_data_hi_8,field_data_lo_8}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_57 = _T_857 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1152 = opcode_28 == 4'h8 | opcode_28 == 4'hb ? _field_data_T_295 : _GEN_1150; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1153 = opcode_28 == 4'h8 | opcode_28 == 4'hb ? _field_tag_T_57 : _GEN_1151; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1154 = 14'h14 == field_data_lo_8 ? _field_data_T_24 : _GEN_1152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1155 = 14'h15 == field_data_lo_8 ? _field_data_T_25 : _GEN_1154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1156 = 14'h16 == field_data_lo_8 ? _field_data_T_26 : _GEN_1155; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1157 = 14'h17 == field_data_lo_8 ? _field_data_T_27 : _GEN_1156; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1158 = 14'h18 == field_data_lo_8 ? _field_data_T_28 : _GEN_1157; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1159 = 14'h19 == field_data_lo_8 ? _field_data_T_29 : _GEN_1158; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1160 = 14'h1a == field_data_lo_8 ? _field_data_T_30 : _GEN_1159; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1161 = 14'h1b == field_data_lo_8 ? _field_data_T_31 : _GEN_1160; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1162 = 14'h1c == field_data_lo_8 ? _field_data_T_32 : _GEN_1161; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1163 = 14'h1d == field_data_lo_8 ? _field_data_T_33 : _GEN_1162; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1164 = 14'h1e == field_data_lo_8 ? _field_data_T_34 : _GEN_1163; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1165 = 14'h1f == field_data_lo_8 ? _field_data_T_35 : _GEN_1164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1166 = 14'h20 == field_data_lo_8 ? _field_data_T_36 : _GEN_1165; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1167 = 14'h21 == field_data_lo_8 ? _field_data_T_37 : _GEN_1166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1168 = 14'h22 == field_data_lo_8 ? _field_data_T_38 : _GEN_1167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1169 = 14'h23 == field_data_lo_8 ? _field_data_T_39 : _GEN_1168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1170 = 14'h24 == field_data_lo_8 ? _field_data_T_40 : _GEN_1169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1171 = 14'h25 == field_data_lo_8 ? _field_data_T_41 : _GEN_1170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1172 = 14'h26 == field_data_lo_8 ? _field_data_T_42 : _GEN_1171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1173 = 14'h27 == field_data_lo_8 ? _field_data_T_43 : _GEN_1172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1174 = 14'h28 == field_data_lo_8 ? _field_data_T_44 : _GEN_1173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1175 = 14'h29 == field_data_lo_8 ? _field_data_T_45 : _GEN_1174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1176 = 14'h2a == field_data_lo_8 ? _field_data_T_46 : _GEN_1175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1177 = 14'h2b == field_data_lo_8 ? _field_data_T_47 : _GEN_1176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1178 = 14'h2c == field_data_lo_8 ? _field_data_T_48 : _GEN_1177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1179 = 14'h2d == field_data_lo_8 ? _field_data_T_49 : _GEN_1178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1180 = 14'h2e == field_data_lo_8 ? _field_data_T_50 : _GEN_1179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1181 = 14'h2f == field_data_lo_8 ? _field_data_T_51 : _GEN_1180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1182 = 14'h30 == field_data_lo_8 ? _field_data_T_52 : _GEN_1181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1183 = 14'h31 == field_data_lo_8 ? _field_data_T_53 : _GEN_1182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_29 = vliw_29[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_9 = vliw_29[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_29 = field_data_lo_9[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_29 = field_data_lo_9[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_38 = {{1'd0}, args_offset_29}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_38 = _total_offset_T_38[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1187 = 3'h1 == total_offset_38 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1188 = 3'h2 == total_offset_38 ? args_2 : _GEN_1187; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1189 = 3'h3 == total_offset_38 ? args_3 : _GEN_1188; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1190 = 3'h4 == total_offset_38 ? args_4 : _GEN_1189; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1191 = 3'h5 == total_offset_38 ? args_5 : _GEN_1190; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1192 = 3'h6 == total_offset_38 ? args_6 : _GEN_1191; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1193 = total_offset_38 < 3'h7 ? _GEN_1192 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_29_1 = 3'h0 < args_length_29 ? _GEN_1193 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_39 = args_offset_29 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1196 = 3'h1 == total_offset_39 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1197 = 3'h2 == total_offset_39 ? args_2 : _GEN_1196; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1198 = 3'h3 == total_offset_39 ? args_3 : _GEN_1197; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1199 = 3'h4 == total_offset_39 ? args_4 : _GEN_1198; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1200 = 3'h5 == total_offset_39 ? args_5 : _GEN_1199; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1201 = 3'h6 == total_offset_39 ? args_6 : _GEN_1200; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1202 = total_offset_39 < 3'h7 ? _GEN_1201 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_29_0 = 3'h1 < args_length_29 ? _GEN_1202 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_326 = {field_bytes_29_0,field_bytes_29_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1204 = opcode_29 == 4'ha ? _field_data_T_326 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1205 = opcode_29 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_896 = opcode_29 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_9 = field_data_lo_9[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_329 = {field_data_hi_9,field_data_lo_9}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_59 = _T_896 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1206 = opcode_29 == 4'h8 | opcode_29 == 4'hb ? _field_data_T_329 : _GEN_1204; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1207 = opcode_29 == 4'h8 | opcode_29 == 4'hb ? _field_tag_T_59 : _GEN_1205; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1208 = 14'h14 == field_data_lo_9 ? _field_data_T_24 : _GEN_1206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1209 = 14'h15 == field_data_lo_9 ? _field_data_T_25 : _GEN_1208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1210 = 14'h16 == field_data_lo_9 ? _field_data_T_26 : _GEN_1209; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1211 = 14'h17 == field_data_lo_9 ? _field_data_T_27 : _GEN_1210; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1212 = 14'h18 == field_data_lo_9 ? _field_data_T_28 : _GEN_1211; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1213 = 14'h19 == field_data_lo_9 ? _field_data_T_29 : _GEN_1212; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1214 = 14'h1a == field_data_lo_9 ? _field_data_T_30 : _GEN_1213; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1215 = 14'h1b == field_data_lo_9 ? _field_data_T_31 : _GEN_1214; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1216 = 14'h1c == field_data_lo_9 ? _field_data_T_32 : _GEN_1215; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1217 = 14'h1d == field_data_lo_9 ? _field_data_T_33 : _GEN_1216; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1218 = 14'h1e == field_data_lo_9 ? _field_data_T_34 : _GEN_1217; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1219 = 14'h1f == field_data_lo_9 ? _field_data_T_35 : _GEN_1218; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1220 = 14'h20 == field_data_lo_9 ? _field_data_T_36 : _GEN_1219; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1221 = 14'h21 == field_data_lo_9 ? _field_data_T_37 : _GEN_1220; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1222 = 14'h22 == field_data_lo_9 ? _field_data_T_38 : _GEN_1221; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1223 = 14'h23 == field_data_lo_9 ? _field_data_T_39 : _GEN_1222; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1224 = 14'h24 == field_data_lo_9 ? _field_data_T_40 : _GEN_1223; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1225 = 14'h25 == field_data_lo_9 ? _field_data_T_41 : _GEN_1224; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1226 = 14'h26 == field_data_lo_9 ? _field_data_T_42 : _GEN_1225; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1227 = 14'h27 == field_data_lo_9 ? _field_data_T_43 : _GEN_1226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1228 = 14'h28 == field_data_lo_9 ? _field_data_T_44 : _GEN_1227; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1229 = 14'h29 == field_data_lo_9 ? _field_data_T_45 : _GEN_1228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1230 = 14'h2a == field_data_lo_9 ? _field_data_T_46 : _GEN_1229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1231 = 14'h2b == field_data_lo_9 ? _field_data_T_47 : _GEN_1230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1232 = 14'h2c == field_data_lo_9 ? _field_data_T_48 : _GEN_1231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1233 = 14'h2d == field_data_lo_9 ? _field_data_T_49 : _GEN_1232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1234 = 14'h2e == field_data_lo_9 ? _field_data_T_50 : _GEN_1233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1235 = 14'h2f == field_data_lo_9 ? _field_data_T_51 : _GEN_1234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1236 = 14'h30 == field_data_lo_9 ? _field_data_T_52 : _GEN_1235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1237 = 14'h31 == field_data_lo_9 ? _field_data_T_53 : _GEN_1236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_30 = vliw_30[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_10 = vliw_30[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_30 = field_data_lo_10[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_30 = field_data_lo_10[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_40 = {{1'd0}, args_offset_30}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_40 = _total_offset_T_40[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1241 = 3'h1 == total_offset_40 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1242 = 3'h2 == total_offset_40 ? args_2 : _GEN_1241; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1243 = 3'h3 == total_offset_40 ? args_3 : _GEN_1242; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1244 = 3'h4 == total_offset_40 ? args_4 : _GEN_1243; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1245 = 3'h5 == total_offset_40 ? args_5 : _GEN_1244; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1246 = 3'h6 == total_offset_40 ? args_6 : _GEN_1245; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1247 = total_offset_40 < 3'h7 ? _GEN_1246 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_30_1 = 3'h0 < args_length_30 ? _GEN_1247 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_41 = args_offset_30 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1250 = 3'h1 == total_offset_41 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1251 = 3'h2 == total_offset_41 ? args_2 : _GEN_1250; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1252 = 3'h3 == total_offset_41 ? args_3 : _GEN_1251; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1253 = 3'h4 == total_offset_41 ? args_4 : _GEN_1252; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1254 = 3'h5 == total_offset_41 ? args_5 : _GEN_1253; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1255 = 3'h6 == total_offset_41 ? args_6 : _GEN_1254; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1256 = total_offset_41 < 3'h7 ? _GEN_1255 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_30_0 = 3'h1 < args_length_30 ? _GEN_1256 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_360 = {field_bytes_30_0,field_bytes_30_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1258 = opcode_30 == 4'ha ? _field_data_T_360 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1259 = opcode_30 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_935 = opcode_30 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_10 = field_data_lo_10[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_363 = {field_data_hi_10,field_data_lo_10}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_61 = _T_935 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1260 = opcode_30 == 4'h8 | opcode_30 == 4'hb ? _field_data_T_363 : _GEN_1258; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1261 = opcode_30 == 4'h8 | opcode_30 == 4'hb ? _field_tag_T_61 : _GEN_1259; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1262 = 14'h14 == field_data_lo_10 ? _field_data_T_24 : _GEN_1260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1263 = 14'h15 == field_data_lo_10 ? _field_data_T_25 : _GEN_1262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1264 = 14'h16 == field_data_lo_10 ? _field_data_T_26 : _GEN_1263; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1265 = 14'h17 == field_data_lo_10 ? _field_data_T_27 : _GEN_1264; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1266 = 14'h18 == field_data_lo_10 ? _field_data_T_28 : _GEN_1265; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1267 = 14'h19 == field_data_lo_10 ? _field_data_T_29 : _GEN_1266; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1268 = 14'h1a == field_data_lo_10 ? _field_data_T_30 : _GEN_1267; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1269 = 14'h1b == field_data_lo_10 ? _field_data_T_31 : _GEN_1268; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1270 = 14'h1c == field_data_lo_10 ? _field_data_T_32 : _GEN_1269; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1271 = 14'h1d == field_data_lo_10 ? _field_data_T_33 : _GEN_1270; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1272 = 14'h1e == field_data_lo_10 ? _field_data_T_34 : _GEN_1271; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1273 = 14'h1f == field_data_lo_10 ? _field_data_T_35 : _GEN_1272; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1274 = 14'h20 == field_data_lo_10 ? _field_data_T_36 : _GEN_1273; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1275 = 14'h21 == field_data_lo_10 ? _field_data_T_37 : _GEN_1274; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1276 = 14'h22 == field_data_lo_10 ? _field_data_T_38 : _GEN_1275; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1277 = 14'h23 == field_data_lo_10 ? _field_data_T_39 : _GEN_1276; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1278 = 14'h24 == field_data_lo_10 ? _field_data_T_40 : _GEN_1277; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1279 = 14'h25 == field_data_lo_10 ? _field_data_T_41 : _GEN_1278; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1280 = 14'h26 == field_data_lo_10 ? _field_data_T_42 : _GEN_1279; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1281 = 14'h27 == field_data_lo_10 ? _field_data_T_43 : _GEN_1280; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1282 = 14'h28 == field_data_lo_10 ? _field_data_T_44 : _GEN_1281; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1283 = 14'h29 == field_data_lo_10 ? _field_data_T_45 : _GEN_1282; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1284 = 14'h2a == field_data_lo_10 ? _field_data_T_46 : _GEN_1283; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1285 = 14'h2b == field_data_lo_10 ? _field_data_T_47 : _GEN_1284; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1286 = 14'h2c == field_data_lo_10 ? _field_data_T_48 : _GEN_1285; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1287 = 14'h2d == field_data_lo_10 ? _field_data_T_49 : _GEN_1286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1288 = 14'h2e == field_data_lo_10 ? _field_data_T_50 : _GEN_1287; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1289 = 14'h2f == field_data_lo_10 ? _field_data_T_51 : _GEN_1288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1290 = 14'h30 == field_data_lo_10 ? _field_data_T_52 : _GEN_1289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1291 = 14'h31 == field_data_lo_10 ? _field_data_T_53 : _GEN_1290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_31 = vliw_31[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_11 = vliw_31[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_31 = field_data_lo_11[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_31 = field_data_lo_11[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_42 = {{1'd0}, args_offset_31}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_42 = _total_offset_T_42[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1295 = 3'h1 == total_offset_42 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1296 = 3'h2 == total_offset_42 ? args_2 : _GEN_1295; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1297 = 3'h3 == total_offset_42 ? args_3 : _GEN_1296; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1298 = 3'h4 == total_offset_42 ? args_4 : _GEN_1297; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1299 = 3'h5 == total_offset_42 ? args_5 : _GEN_1298; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1300 = 3'h6 == total_offset_42 ? args_6 : _GEN_1299; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1301 = total_offset_42 < 3'h7 ? _GEN_1300 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_31_1 = 3'h0 < args_length_31 ? _GEN_1301 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_43 = args_offset_31 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1304 = 3'h1 == total_offset_43 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1305 = 3'h2 == total_offset_43 ? args_2 : _GEN_1304; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1306 = 3'h3 == total_offset_43 ? args_3 : _GEN_1305; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1307 = 3'h4 == total_offset_43 ? args_4 : _GEN_1306; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1308 = 3'h5 == total_offset_43 ? args_5 : _GEN_1307; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1309 = 3'h6 == total_offset_43 ? args_6 : _GEN_1308; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1310 = total_offset_43 < 3'h7 ? _GEN_1309 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_31_0 = 3'h1 < args_length_31 ? _GEN_1310 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_394 = {field_bytes_31_0,field_bytes_31_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1312 = opcode_31 == 4'ha ? _field_data_T_394 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1313 = opcode_31 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_974 = opcode_31 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_11 = field_data_lo_11[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_397 = {field_data_hi_11,field_data_lo_11}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_63 = _T_974 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1314 = opcode_31 == 4'h8 | opcode_31 == 4'hb ? _field_data_T_397 : _GEN_1312; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1315 = opcode_31 == 4'h8 | opcode_31 == 4'hb ? _field_tag_T_63 : _GEN_1313; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1316 = 14'h14 == field_data_lo_11 ? _field_data_T_24 : _GEN_1314; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1317 = 14'h15 == field_data_lo_11 ? _field_data_T_25 : _GEN_1316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1318 = 14'h16 == field_data_lo_11 ? _field_data_T_26 : _GEN_1317; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1319 = 14'h17 == field_data_lo_11 ? _field_data_T_27 : _GEN_1318; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1320 = 14'h18 == field_data_lo_11 ? _field_data_T_28 : _GEN_1319; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1321 = 14'h19 == field_data_lo_11 ? _field_data_T_29 : _GEN_1320; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1322 = 14'h1a == field_data_lo_11 ? _field_data_T_30 : _GEN_1321; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1323 = 14'h1b == field_data_lo_11 ? _field_data_T_31 : _GEN_1322; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1324 = 14'h1c == field_data_lo_11 ? _field_data_T_32 : _GEN_1323; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1325 = 14'h1d == field_data_lo_11 ? _field_data_T_33 : _GEN_1324; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1326 = 14'h1e == field_data_lo_11 ? _field_data_T_34 : _GEN_1325; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1327 = 14'h1f == field_data_lo_11 ? _field_data_T_35 : _GEN_1326; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1328 = 14'h20 == field_data_lo_11 ? _field_data_T_36 : _GEN_1327; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1329 = 14'h21 == field_data_lo_11 ? _field_data_T_37 : _GEN_1328; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1330 = 14'h22 == field_data_lo_11 ? _field_data_T_38 : _GEN_1329; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1331 = 14'h23 == field_data_lo_11 ? _field_data_T_39 : _GEN_1330; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1332 = 14'h24 == field_data_lo_11 ? _field_data_T_40 : _GEN_1331; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1333 = 14'h25 == field_data_lo_11 ? _field_data_T_41 : _GEN_1332; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1334 = 14'h26 == field_data_lo_11 ? _field_data_T_42 : _GEN_1333; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1335 = 14'h27 == field_data_lo_11 ? _field_data_T_43 : _GEN_1334; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1336 = 14'h28 == field_data_lo_11 ? _field_data_T_44 : _GEN_1335; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1337 = 14'h29 == field_data_lo_11 ? _field_data_T_45 : _GEN_1336; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1338 = 14'h2a == field_data_lo_11 ? _field_data_T_46 : _GEN_1337; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1339 = 14'h2b == field_data_lo_11 ? _field_data_T_47 : _GEN_1338; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1340 = 14'h2c == field_data_lo_11 ? _field_data_T_48 : _GEN_1339; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1341 = 14'h2d == field_data_lo_11 ? _field_data_T_49 : _GEN_1340; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1342 = 14'h2e == field_data_lo_11 ? _field_data_T_50 : _GEN_1341; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1343 = 14'h2f == field_data_lo_11 ? _field_data_T_51 : _GEN_1342; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1344 = 14'h30 == field_data_lo_11 ? _field_data_T_52 : _GEN_1343; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1345 = 14'h31 == field_data_lo_11 ? _field_data_T_53 : _GEN_1344; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_32 = vliw_32[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_12 = vliw_32[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_32 = field_data_lo_12[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_32 = field_data_lo_12[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_44 = {{1'd0}, args_offset_32}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_44 = _total_offset_T_44[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1349 = 3'h1 == total_offset_44 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1350 = 3'h2 == total_offset_44 ? args_2 : _GEN_1349; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1351 = 3'h3 == total_offset_44 ? args_3 : _GEN_1350; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1352 = 3'h4 == total_offset_44 ? args_4 : _GEN_1351; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1353 = 3'h5 == total_offset_44 ? args_5 : _GEN_1352; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1354 = 3'h6 == total_offset_44 ? args_6 : _GEN_1353; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1355 = total_offset_44 < 3'h7 ? _GEN_1354 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_32_1 = 3'h0 < args_length_32 ? _GEN_1355 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_45 = args_offset_32 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1358 = 3'h1 == total_offset_45 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1359 = 3'h2 == total_offset_45 ? args_2 : _GEN_1358; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1360 = 3'h3 == total_offset_45 ? args_3 : _GEN_1359; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1361 = 3'h4 == total_offset_45 ? args_4 : _GEN_1360; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1362 = 3'h5 == total_offset_45 ? args_5 : _GEN_1361; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1363 = 3'h6 == total_offset_45 ? args_6 : _GEN_1362; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1364 = total_offset_45 < 3'h7 ? _GEN_1363 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_32_0 = 3'h1 < args_length_32 ? _GEN_1364 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_428 = {field_bytes_32_0,field_bytes_32_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1366 = opcode_32 == 4'ha ? _field_data_T_428 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1367 = opcode_32 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1013 = opcode_32 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_12 = field_data_lo_12[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_431 = {field_data_hi_12,field_data_lo_12}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_65 = _T_1013 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1368 = opcode_32 == 4'h8 | opcode_32 == 4'hb ? _field_data_T_431 : _GEN_1366; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1369 = opcode_32 == 4'h8 | opcode_32 == 4'hb ? _field_tag_T_65 : _GEN_1367; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1370 = 14'h14 == field_data_lo_12 ? _field_data_T_24 : _GEN_1368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1371 = 14'h15 == field_data_lo_12 ? _field_data_T_25 : _GEN_1370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1372 = 14'h16 == field_data_lo_12 ? _field_data_T_26 : _GEN_1371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1373 = 14'h17 == field_data_lo_12 ? _field_data_T_27 : _GEN_1372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1374 = 14'h18 == field_data_lo_12 ? _field_data_T_28 : _GEN_1373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1375 = 14'h19 == field_data_lo_12 ? _field_data_T_29 : _GEN_1374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1376 = 14'h1a == field_data_lo_12 ? _field_data_T_30 : _GEN_1375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1377 = 14'h1b == field_data_lo_12 ? _field_data_T_31 : _GEN_1376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1378 = 14'h1c == field_data_lo_12 ? _field_data_T_32 : _GEN_1377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1379 = 14'h1d == field_data_lo_12 ? _field_data_T_33 : _GEN_1378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1380 = 14'h1e == field_data_lo_12 ? _field_data_T_34 : _GEN_1379; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1381 = 14'h1f == field_data_lo_12 ? _field_data_T_35 : _GEN_1380; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1382 = 14'h20 == field_data_lo_12 ? _field_data_T_36 : _GEN_1381; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1383 = 14'h21 == field_data_lo_12 ? _field_data_T_37 : _GEN_1382; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1384 = 14'h22 == field_data_lo_12 ? _field_data_T_38 : _GEN_1383; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1385 = 14'h23 == field_data_lo_12 ? _field_data_T_39 : _GEN_1384; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1386 = 14'h24 == field_data_lo_12 ? _field_data_T_40 : _GEN_1385; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1387 = 14'h25 == field_data_lo_12 ? _field_data_T_41 : _GEN_1386; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1388 = 14'h26 == field_data_lo_12 ? _field_data_T_42 : _GEN_1387; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1389 = 14'h27 == field_data_lo_12 ? _field_data_T_43 : _GEN_1388; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1390 = 14'h28 == field_data_lo_12 ? _field_data_T_44 : _GEN_1389; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1391 = 14'h29 == field_data_lo_12 ? _field_data_T_45 : _GEN_1390; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1392 = 14'h2a == field_data_lo_12 ? _field_data_T_46 : _GEN_1391; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1393 = 14'h2b == field_data_lo_12 ? _field_data_T_47 : _GEN_1392; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1394 = 14'h2c == field_data_lo_12 ? _field_data_T_48 : _GEN_1393; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1395 = 14'h2d == field_data_lo_12 ? _field_data_T_49 : _GEN_1394; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1396 = 14'h2e == field_data_lo_12 ? _field_data_T_50 : _GEN_1395; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1397 = 14'h2f == field_data_lo_12 ? _field_data_T_51 : _GEN_1396; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1398 = 14'h30 == field_data_lo_12 ? _field_data_T_52 : _GEN_1397; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1399 = 14'h31 == field_data_lo_12 ? _field_data_T_53 : _GEN_1398; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_33 = vliw_33[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_13 = vliw_33[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_33 = field_data_lo_13[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_33 = field_data_lo_13[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_46 = {{1'd0}, args_offset_33}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_46 = _total_offset_T_46[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1403 = 3'h1 == total_offset_46 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1404 = 3'h2 == total_offset_46 ? args_2 : _GEN_1403; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1405 = 3'h3 == total_offset_46 ? args_3 : _GEN_1404; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1406 = 3'h4 == total_offset_46 ? args_4 : _GEN_1405; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1407 = 3'h5 == total_offset_46 ? args_5 : _GEN_1406; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1408 = 3'h6 == total_offset_46 ? args_6 : _GEN_1407; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1409 = total_offset_46 < 3'h7 ? _GEN_1408 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_33_1 = 3'h0 < args_length_33 ? _GEN_1409 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_47 = args_offset_33 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1412 = 3'h1 == total_offset_47 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1413 = 3'h2 == total_offset_47 ? args_2 : _GEN_1412; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1414 = 3'h3 == total_offset_47 ? args_3 : _GEN_1413; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1415 = 3'h4 == total_offset_47 ? args_4 : _GEN_1414; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1416 = 3'h5 == total_offset_47 ? args_5 : _GEN_1415; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1417 = 3'h6 == total_offset_47 ? args_6 : _GEN_1416; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1418 = total_offset_47 < 3'h7 ? _GEN_1417 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_33_0 = 3'h1 < args_length_33 ? _GEN_1418 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_462 = {field_bytes_33_0,field_bytes_33_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1420 = opcode_33 == 4'ha ? _field_data_T_462 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1421 = opcode_33 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1052 = opcode_33 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_13 = field_data_lo_13[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_465 = {field_data_hi_13,field_data_lo_13}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_67 = _T_1052 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1422 = opcode_33 == 4'h8 | opcode_33 == 4'hb ? _field_data_T_465 : _GEN_1420; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1423 = opcode_33 == 4'h8 | opcode_33 == 4'hb ? _field_tag_T_67 : _GEN_1421; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1424 = 14'h14 == field_data_lo_13 ? _field_data_T_24 : _GEN_1422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1425 = 14'h15 == field_data_lo_13 ? _field_data_T_25 : _GEN_1424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1426 = 14'h16 == field_data_lo_13 ? _field_data_T_26 : _GEN_1425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1427 = 14'h17 == field_data_lo_13 ? _field_data_T_27 : _GEN_1426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1428 = 14'h18 == field_data_lo_13 ? _field_data_T_28 : _GEN_1427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1429 = 14'h19 == field_data_lo_13 ? _field_data_T_29 : _GEN_1428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1430 = 14'h1a == field_data_lo_13 ? _field_data_T_30 : _GEN_1429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1431 = 14'h1b == field_data_lo_13 ? _field_data_T_31 : _GEN_1430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1432 = 14'h1c == field_data_lo_13 ? _field_data_T_32 : _GEN_1431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1433 = 14'h1d == field_data_lo_13 ? _field_data_T_33 : _GEN_1432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1434 = 14'h1e == field_data_lo_13 ? _field_data_T_34 : _GEN_1433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1435 = 14'h1f == field_data_lo_13 ? _field_data_T_35 : _GEN_1434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1436 = 14'h20 == field_data_lo_13 ? _field_data_T_36 : _GEN_1435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1437 = 14'h21 == field_data_lo_13 ? _field_data_T_37 : _GEN_1436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1438 = 14'h22 == field_data_lo_13 ? _field_data_T_38 : _GEN_1437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1439 = 14'h23 == field_data_lo_13 ? _field_data_T_39 : _GEN_1438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1440 = 14'h24 == field_data_lo_13 ? _field_data_T_40 : _GEN_1439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1441 = 14'h25 == field_data_lo_13 ? _field_data_T_41 : _GEN_1440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1442 = 14'h26 == field_data_lo_13 ? _field_data_T_42 : _GEN_1441; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1443 = 14'h27 == field_data_lo_13 ? _field_data_T_43 : _GEN_1442; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1444 = 14'h28 == field_data_lo_13 ? _field_data_T_44 : _GEN_1443; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1445 = 14'h29 == field_data_lo_13 ? _field_data_T_45 : _GEN_1444; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1446 = 14'h2a == field_data_lo_13 ? _field_data_T_46 : _GEN_1445; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1447 = 14'h2b == field_data_lo_13 ? _field_data_T_47 : _GEN_1446; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1448 = 14'h2c == field_data_lo_13 ? _field_data_T_48 : _GEN_1447; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1449 = 14'h2d == field_data_lo_13 ? _field_data_T_49 : _GEN_1448; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1450 = 14'h2e == field_data_lo_13 ? _field_data_T_50 : _GEN_1449; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1451 = 14'h2f == field_data_lo_13 ? _field_data_T_51 : _GEN_1450; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1452 = 14'h30 == field_data_lo_13 ? _field_data_T_52 : _GEN_1451; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1453 = 14'h31 == field_data_lo_13 ? _field_data_T_53 : _GEN_1452; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_34 = vliw_34[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_14 = vliw_34[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_34 = field_data_lo_14[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_34 = field_data_lo_14[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_48 = {{1'd0}, args_offset_34}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_48 = _total_offset_T_48[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1457 = 3'h1 == total_offset_48 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1458 = 3'h2 == total_offset_48 ? args_2 : _GEN_1457; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1459 = 3'h3 == total_offset_48 ? args_3 : _GEN_1458; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1460 = 3'h4 == total_offset_48 ? args_4 : _GEN_1459; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1461 = 3'h5 == total_offset_48 ? args_5 : _GEN_1460; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1462 = 3'h6 == total_offset_48 ? args_6 : _GEN_1461; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1463 = total_offset_48 < 3'h7 ? _GEN_1462 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_34_1 = 3'h0 < args_length_34 ? _GEN_1463 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_49 = args_offset_34 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1466 = 3'h1 == total_offset_49 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1467 = 3'h2 == total_offset_49 ? args_2 : _GEN_1466; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1468 = 3'h3 == total_offset_49 ? args_3 : _GEN_1467; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1469 = 3'h4 == total_offset_49 ? args_4 : _GEN_1468; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1470 = 3'h5 == total_offset_49 ? args_5 : _GEN_1469; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1471 = 3'h6 == total_offset_49 ? args_6 : _GEN_1470; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1472 = total_offset_49 < 3'h7 ? _GEN_1471 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_34_0 = 3'h1 < args_length_34 ? _GEN_1472 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_496 = {field_bytes_34_0,field_bytes_34_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1474 = opcode_34 == 4'ha ? _field_data_T_496 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1475 = opcode_34 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1091 = opcode_34 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_14 = field_data_lo_14[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_499 = {field_data_hi_14,field_data_lo_14}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_69 = _T_1091 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1476 = opcode_34 == 4'h8 | opcode_34 == 4'hb ? _field_data_T_499 : _GEN_1474; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1477 = opcode_34 == 4'h8 | opcode_34 == 4'hb ? _field_tag_T_69 : _GEN_1475; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1478 = 14'h14 == field_data_lo_14 ? _field_data_T_24 : _GEN_1476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1479 = 14'h15 == field_data_lo_14 ? _field_data_T_25 : _GEN_1478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1480 = 14'h16 == field_data_lo_14 ? _field_data_T_26 : _GEN_1479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1481 = 14'h17 == field_data_lo_14 ? _field_data_T_27 : _GEN_1480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1482 = 14'h18 == field_data_lo_14 ? _field_data_T_28 : _GEN_1481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1483 = 14'h19 == field_data_lo_14 ? _field_data_T_29 : _GEN_1482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1484 = 14'h1a == field_data_lo_14 ? _field_data_T_30 : _GEN_1483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1485 = 14'h1b == field_data_lo_14 ? _field_data_T_31 : _GEN_1484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1486 = 14'h1c == field_data_lo_14 ? _field_data_T_32 : _GEN_1485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1487 = 14'h1d == field_data_lo_14 ? _field_data_T_33 : _GEN_1486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1488 = 14'h1e == field_data_lo_14 ? _field_data_T_34 : _GEN_1487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1489 = 14'h1f == field_data_lo_14 ? _field_data_T_35 : _GEN_1488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1490 = 14'h20 == field_data_lo_14 ? _field_data_T_36 : _GEN_1489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1491 = 14'h21 == field_data_lo_14 ? _field_data_T_37 : _GEN_1490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1492 = 14'h22 == field_data_lo_14 ? _field_data_T_38 : _GEN_1491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1493 = 14'h23 == field_data_lo_14 ? _field_data_T_39 : _GEN_1492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1494 = 14'h24 == field_data_lo_14 ? _field_data_T_40 : _GEN_1493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1495 = 14'h25 == field_data_lo_14 ? _field_data_T_41 : _GEN_1494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1496 = 14'h26 == field_data_lo_14 ? _field_data_T_42 : _GEN_1495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1497 = 14'h27 == field_data_lo_14 ? _field_data_T_43 : _GEN_1496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1498 = 14'h28 == field_data_lo_14 ? _field_data_T_44 : _GEN_1497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1499 = 14'h29 == field_data_lo_14 ? _field_data_T_45 : _GEN_1498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1500 = 14'h2a == field_data_lo_14 ? _field_data_T_46 : _GEN_1499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1501 = 14'h2b == field_data_lo_14 ? _field_data_T_47 : _GEN_1500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1502 = 14'h2c == field_data_lo_14 ? _field_data_T_48 : _GEN_1501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1503 = 14'h2d == field_data_lo_14 ? _field_data_T_49 : _GEN_1502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1504 = 14'h2e == field_data_lo_14 ? _field_data_T_50 : _GEN_1503; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1505 = 14'h2f == field_data_lo_14 ? _field_data_T_51 : _GEN_1504; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1506 = 14'h30 == field_data_lo_14 ? _field_data_T_52 : _GEN_1505; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1507 = 14'h31 == field_data_lo_14 ? _field_data_T_53 : _GEN_1506; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_35 = vliw_35[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_15 = vliw_35[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_35 = field_data_lo_15[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_35 = field_data_lo_15[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_50 = {{1'd0}, args_offset_35}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_50 = _total_offset_T_50[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1511 = 3'h1 == total_offset_50 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1512 = 3'h2 == total_offset_50 ? args_2 : _GEN_1511; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1513 = 3'h3 == total_offset_50 ? args_3 : _GEN_1512; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1514 = 3'h4 == total_offset_50 ? args_4 : _GEN_1513; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1515 = 3'h5 == total_offset_50 ? args_5 : _GEN_1514; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1516 = 3'h6 == total_offset_50 ? args_6 : _GEN_1515; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1517 = total_offset_50 < 3'h7 ? _GEN_1516 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_35_1 = 3'h0 < args_length_35 ? _GEN_1517 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_51 = args_offset_35 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1520 = 3'h1 == total_offset_51 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1521 = 3'h2 == total_offset_51 ? args_2 : _GEN_1520; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1522 = 3'h3 == total_offset_51 ? args_3 : _GEN_1521; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1523 = 3'h4 == total_offset_51 ? args_4 : _GEN_1522; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1524 = 3'h5 == total_offset_51 ? args_5 : _GEN_1523; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1525 = 3'h6 == total_offset_51 ? args_6 : _GEN_1524; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1526 = total_offset_51 < 3'h7 ? _GEN_1525 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_35_0 = 3'h1 < args_length_35 ? _GEN_1526 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_530 = {field_bytes_35_0,field_bytes_35_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1528 = opcode_35 == 4'ha ? _field_data_T_530 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1529 = opcode_35 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1130 = opcode_35 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_15 = field_data_lo_15[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_533 = {field_data_hi_15,field_data_lo_15}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_71 = _T_1130 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1530 = opcode_35 == 4'h8 | opcode_35 == 4'hb ? _field_data_T_533 : _GEN_1528; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1531 = opcode_35 == 4'h8 | opcode_35 == 4'hb ? _field_tag_T_71 : _GEN_1529; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1532 = 14'h14 == field_data_lo_15 ? _field_data_T_24 : _GEN_1530; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1533 = 14'h15 == field_data_lo_15 ? _field_data_T_25 : _GEN_1532; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1534 = 14'h16 == field_data_lo_15 ? _field_data_T_26 : _GEN_1533; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1535 = 14'h17 == field_data_lo_15 ? _field_data_T_27 : _GEN_1534; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1536 = 14'h18 == field_data_lo_15 ? _field_data_T_28 : _GEN_1535; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1537 = 14'h19 == field_data_lo_15 ? _field_data_T_29 : _GEN_1536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1538 = 14'h1a == field_data_lo_15 ? _field_data_T_30 : _GEN_1537; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1539 = 14'h1b == field_data_lo_15 ? _field_data_T_31 : _GEN_1538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1540 = 14'h1c == field_data_lo_15 ? _field_data_T_32 : _GEN_1539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1541 = 14'h1d == field_data_lo_15 ? _field_data_T_33 : _GEN_1540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1542 = 14'h1e == field_data_lo_15 ? _field_data_T_34 : _GEN_1541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1543 = 14'h1f == field_data_lo_15 ? _field_data_T_35 : _GEN_1542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1544 = 14'h20 == field_data_lo_15 ? _field_data_T_36 : _GEN_1543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1545 = 14'h21 == field_data_lo_15 ? _field_data_T_37 : _GEN_1544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1546 = 14'h22 == field_data_lo_15 ? _field_data_T_38 : _GEN_1545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1547 = 14'h23 == field_data_lo_15 ? _field_data_T_39 : _GEN_1546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1548 = 14'h24 == field_data_lo_15 ? _field_data_T_40 : _GEN_1547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1549 = 14'h25 == field_data_lo_15 ? _field_data_T_41 : _GEN_1548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1550 = 14'h26 == field_data_lo_15 ? _field_data_T_42 : _GEN_1549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1551 = 14'h27 == field_data_lo_15 ? _field_data_T_43 : _GEN_1550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1552 = 14'h28 == field_data_lo_15 ? _field_data_T_44 : _GEN_1551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1553 = 14'h29 == field_data_lo_15 ? _field_data_T_45 : _GEN_1552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1554 = 14'h2a == field_data_lo_15 ? _field_data_T_46 : _GEN_1553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1555 = 14'h2b == field_data_lo_15 ? _field_data_T_47 : _GEN_1554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1556 = 14'h2c == field_data_lo_15 ? _field_data_T_48 : _GEN_1555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1557 = 14'h2d == field_data_lo_15 ? _field_data_T_49 : _GEN_1556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1558 = 14'h2e == field_data_lo_15 ? _field_data_T_50 : _GEN_1557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1559 = 14'h2f == field_data_lo_15 ? _field_data_T_51 : _GEN_1558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1560 = 14'h30 == field_data_lo_15 ? _field_data_T_52 : _GEN_1559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1561 = 14'h31 == field_data_lo_15 ? _field_data_T_53 : _GEN_1560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_36 = vliw_36[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_16 = vliw_36[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_36 = field_data_lo_16[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_36 = field_data_lo_16[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_52 = {{1'd0}, args_offset_36}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_52 = _total_offset_T_52[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1565 = 3'h1 == total_offset_52 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1566 = 3'h2 == total_offset_52 ? args_2 : _GEN_1565; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1567 = 3'h3 == total_offset_52 ? args_3 : _GEN_1566; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1568 = 3'h4 == total_offset_52 ? args_4 : _GEN_1567; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1569 = 3'h5 == total_offset_52 ? args_5 : _GEN_1568; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1570 = 3'h6 == total_offset_52 ? args_6 : _GEN_1569; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1571 = total_offset_52 < 3'h7 ? _GEN_1570 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_36_1 = 3'h0 < args_length_36 ? _GEN_1571 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_53 = args_offset_36 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1574 = 3'h1 == total_offset_53 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1575 = 3'h2 == total_offset_53 ? args_2 : _GEN_1574; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1576 = 3'h3 == total_offset_53 ? args_3 : _GEN_1575; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1577 = 3'h4 == total_offset_53 ? args_4 : _GEN_1576; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1578 = 3'h5 == total_offset_53 ? args_5 : _GEN_1577; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1579 = 3'h6 == total_offset_53 ? args_6 : _GEN_1578; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1580 = total_offset_53 < 3'h7 ? _GEN_1579 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_36_0 = 3'h1 < args_length_36 ? _GEN_1580 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_564 = {field_bytes_36_0,field_bytes_36_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1582 = opcode_36 == 4'ha ? _field_data_T_564 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1583 = opcode_36 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1169 = opcode_36 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_16 = field_data_lo_16[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_567 = {field_data_hi_16,field_data_lo_16}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_73 = _T_1169 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1584 = opcode_36 == 4'h8 | opcode_36 == 4'hb ? _field_data_T_567 : _GEN_1582; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1585 = opcode_36 == 4'h8 | opcode_36 == 4'hb ? _field_tag_T_73 : _GEN_1583; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1586 = 14'h14 == field_data_lo_16 ? _field_data_T_24 : _GEN_1584; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1587 = 14'h15 == field_data_lo_16 ? _field_data_T_25 : _GEN_1586; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1588 = 14'h16 == field_data_lo_16 ? _field_data_T_26 : _GEN_1587; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1589 = 14'h17 == field_data_lo_16 ? _field_data_T_27 : _GEN_1588; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1590 = 14'h18 == field_data_lo_16 ? _field_data_T_28 : _GEN_1589; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1591 = 14'h19 == field_data_lo_16 ? _field_data_T_29 : _GEN_1590; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1592 = 14'h1a == field_data_lo_16 ? _field_data_T_30 : _GEN_1591; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1593 = 14'h1b == field_data_lo_16 ? _field_data_T_31 : _GEN_1592; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1594 = 14'h1c == field_data_lo_16 ? _field_data_T_32 : _GEN_1593; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1595 = 14'h1d == field_data_lo_16 ? _field_data_T_33 : _GEN_1594; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1596 = 14'h1e == field_data_lo_16 ? _field_data_T_34 : _GEN_1595; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1597 = 14'h1f == field_data_lo_16 ? _field_data_T_35 : _GEN_1596; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1598 = 14'h20 == field_data_lo_16 ? _field_data_T_36 : _GEN_1597; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1599 = 14'h21 == field_data_lo_16 ? _field_data_T_37 : _GEN_1598; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1600 = 14'h22 == field_data_lo_16 ? _field_data_T_38 : _GEN_1599; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1601 = 14'h23 == field_data_lo_16 ? _field_data_T_39 : _GEN_1600; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1602 = 14'h24 == field_data_lo_16 ? _field_data_T_40 : _GEN_1601; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1603 = 14'h25 == field_data_lo_16 ? _field_data_T_41 : _GEN_1602; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1604 = 14'h26 == field_data_lo_16 ? _field_data_T_42 : _GEN_1603; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1605 = 14'h27 == field_data_lo_16 ? _field_data_T_43 : _GEN_1604; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1606 = 14'h28 == field_data_lo_16 ? _field_data_T_44 : _GEN_1605; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1607 = 14'h29 == field_data_lo_16 ? _field_data_T_45 : _GEN_1606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1608 = 14'h2a == field_data_lo_16 ? _field_data_T_46 : _GEN_1607; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1609 = 14'h2b == field_data_lo_16 ? _field_data_T_47 : _GEN_1608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1610 = 14'h2c == field_data_lo_16 ? _field_data_T_48 : _GEN_1609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1611 = 14'h2d == field_data_lo_16 ? _field_data_T_49 : _GEN_1610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1612 = 14'h2e == field_data_lo_16 ? _field_data_T_50 : _GEN_1611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1613 = 14'h2f == field_data_lo_16 ? _field_data_T_51 : _GEN_1612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1614 = 14'h30 == field_data_lo_16 ? _field_data_T_52 : _GEN_1613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1615 = 14'h31 == field_data_lo_16 ? _field_data_T_53 : _GEN_1614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_37 = vliw_37[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_17 = vliw_37[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_37 = field_data_lo_17[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_37 = field_data_lo_17[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_54 = {{1'd0}, args_offset_37}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_54 = _total_offset_T_54[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1619 = 3'h1 == total_offset_54 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1620 = 3'h2 == total_offset_54 ? args_2 : _GEN_1619; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1621 = 3'h3 == total_offset_54 ? args_3 : _GEN_1620; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1622 = 3'h4 == total_offset_54 ? args_4 : _GEN_1621; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1623 = 3'h5 == total_offset_54 ? args_5 : _GEN_1622; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1624 = 3'h6 == total_offset_54 ? args_6 : _GEN_1623; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1625 = total_offset_54 < 3'h7 ? _GEN_1624 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_37_1 = 3'h0 < args_length_37 ? _GEN_1625 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_55 = args_offset_37 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1628 = 3'h1 == total_offset_55 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1629 = 3'h2 == total_offset_55 ? args_2 : _GEN_1628; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1630 = 3'h3 == total_offset_55 ? args_3 : _GEN_1629; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1631 = 3'h4 == total_offset_55 ? args_4 : _GEN_1630; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1632 = 3'h5 == total_offset_55 ? args_5 : _GEN_1631; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1633 = 3'h6 == total_offset_55 ? args_6 : _GEN_1632; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1634 = total_offset_55 < 3'h7 ? _GEN_1633 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_37_0 = 3'h1 < args_length_37 ? _GEN_1634 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_598 = {field_bytes_37_0,field_bytes_37_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1636 = opcode_37 == 4'ha ? _field_data_T_598 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1637 = opcode_37 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1208 = opcode_37 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_17 = field_data_lo_17[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_601 = {field_data_hi_17,field_data_lo_17}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_75 = _T_1208 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1638 = opcode_37 == 4'h8 | opcode_37 == 4'hb ? _field_data_T_601 : _GEN_1636; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1639 = opcode_37 == 4'h8 | opcode_37 == 4'hb ? _field_tag_T_75 : _GEN_1637; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1640 = 14'h14 == field_data_lo_17 ? _field_data_T_24 : _GEN_1638; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1641 = 14'h15 == field_data_lo_17 ? _field_data_T_25 : _GEN_1640; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1642 = 14'h16 == field_data_lo_17 ? _field_data_T_26 : _GEN_1641; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1643 = 14'h17 == field_data_lo_17 ? _field_data_T_27 : _GEN_1642; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1644 = 14'h18 == field_data_lo_17 ? _field_data_T_28 : _GEN_1643; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1645 = 14'h19 == field_data_lo_17 ? _field_data_T_29 : _GEN_1644; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1646 = 14'h1a == field_data_lo_17 ? _field_data_T_30 : _GEN_1645; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1647 = 14'h1b == field_data_lo_17 ? _field_data_T_31 : _GEN_1646; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1648 = 14'h1c == field_data_lo_17 ? _field_data_T_32 : _GEN_1647; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1649 = 14'h1d == field_data_lo_17 ? _field_data_T_33 : _GEN_1648; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1650 = 14'h1e == field_data_lo_17 ? _field_data_T_34 : _GEN_1649; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1651 = 14'h1f == field_data_lo_17 ? _field_data_T_35 : _GEN_1650; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1652 = 14'h20 == field_data_lo_17 ? _field_data_T_36 : _GEN_1651; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1653 = 14'h21 == field_data_lo_17 ? _field_data_T_37 : _GEN_1652; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1654 = 14'h22 == field_data_lo_17 ? _field_data_T_38 : _GEN_1653; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1655 = 14'h23 == field_data_lo_17 ? _field_data_T_39 : _GEN_1654; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1656 = 14'h24 == field_data_lo_17 ? _field_data_T_40 : _GEN_1655; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1657 = 14'h25 == field_data_lo_17 ? _field_data_T_41 : _GEN_1656; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1658 = 14'h26 == field_data_lo_17 ? _field_data_T_42 : _GEN_1657; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1659 = 14'h27 == field_data_lo_17 ? _field_data_T_43 : _GEN_1658; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1660 = 14'h28 == field_data_lo_17 ? _field_data_T_44 : _GEN_1659; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1661 = 14'h29 == field_data_lo_17 ? _field_data_T_45 : _GEN_1660; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1662 = 14'h2a == field_data_lo_17 ? _field_data_T_46 : _GEN_1661; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1663 = 14'h2b == field_data_lo_17 ? _field_data_T_47 : _GEN_1662; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1664 = 14'h2c == field_data_lo_17 ? _field_data_T_48 : _GEN_1663; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1665 = 14'h2d == field_data_lo_17 ? _field_data_T_49 : _GEN_1664; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1666 = 14'h2e == field_data_lo_17 ? _field_data_T_50 : _GEN_1665; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1667 = 14'h2f == field_data_lo_17 ? _field_data_T_51 : _GEN_1666; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1668 = 14'h30 == field_data_lo_17 ? _field_data_T_52 : _GEN_1667; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1669 = 14'h31 == field_data_lo_17 ? _field_data_T_53 : _GEN_1668; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_38 = vliw_38[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_18 = vliw_38[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_38 = field_data_lo_18[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_38 = field_data_lo_18[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_56 = {{1'd0}, args_offset_38}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_56 = _total_offset_T_56[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1673 = 3'h1 == total_offset_56 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1674 = 3'h2 == total_offset_56 ? args_2 : _GEN_1673; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1675 = 3'h3 == total_offset_56 ? args_3 : _GEN_1674; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1676 = 3'h4 == total_offset_56 ? args_4 : _GEN_1675; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1677 = 3'h5 == total_offset_56 ? args_5 : _GEN_1676; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1678 = 3'h6 == total_offset_56 ? args_6 : _GEN_1677; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1679 = total_offset_56 < 3'h7 ? _GEN_1678 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_38_1 = 3'h0 < args_length_38 ? _GEN_1679 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_57 = args_offset_38 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1682 = 3'h1 == total_offset_57 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1683 = 3'h2 == total_offset_57 ? args_2 : _GEN_1682; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1684 = 3'h3 == total_offset_57 ? args_3 : _GEN_1683; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1685 = 3'h4 == total_offset_57 ? args_4 : _GEN_1684; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1686 = 3'h5 == total_offset_57 ? args_5 : _GEN_1685; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1687 = 3'h6 == total_offset_57 ? args_6 : _GEN_1686; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1688 = total_offset_57 < 3'h7 ? _GEN_1687 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_38_0 = 3'h1 < args_length_38 ? _GEN_1688 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_632 = {field_bytes_38_0,field_bytes_38_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1690 = opcode_38 == 4'ha ? _field_data_T_632 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1691 = opcode_38 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1247 = opcode_38 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_18 = field_data_lo_18[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_635 = {field_data_hi_18,field_data_lo_18}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_77 = _T_1247 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1692 = opcode_38 == 4'h8 | opcode_38 == 4'hb ? _field_data_T_635 : _GEN_1690; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1693 = opcode_38 == 4'h8 | opcode_38 == 4'hb ? _field_tag_T_77 : _GEN_1691; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1694 = 14'h14 == field_data_lo_18 ? _field_data_T_24 : _GEN_1692; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1695 = 14'h15 == field_data_lo_18 ? _field_data_T_25 : _GEN_1694; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1696 = 14'h16 == field_data_lo_18 ? _field_data_T_26 : _GEN_1695; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1697 = 14'h17 == field_data_lo_18 ? _field_data_T_27 : _GEN_1696; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1698 = 14'h18 == field_data_lo_18 ? _field_data_T_28 : _GEN_1697; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1699 = 14'h19 == field_data_lo_18 ? _field_data_T_29 : _GEN_1698; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1700 = 14'h1a == field_data_lo_18 ? _field_data_T_30 : _GEN_1699; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1701 = 14'h1b == field_data_lo_18 ? _field_data_T_31 : _GEN_1700; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1702 = 14'h1c == field_data_lo_18 ? _field_data_T_32 : _GEN_1701; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1703 = 14'h1d == field_data_lo_18 ? _field_data_T_33 : _GEN_1702; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1704 = 14'h1e == field_data_lo_18 ? _field_data_T_34 : _GEN_1703; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1705 = 14'h1f == field_data_lo_18 ? _field_data_T_35 : _GEN_1704; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1706 = 14'h20 == field_data_lo_18 ? _field_data_T_36 : _GEN_1705; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1707 = 14'h21 == field_data_lo_18 ? _field_data_T_37 : _GEN_1706; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1708 = 14'h22 == field_data_lo_18 ? _field_data_T_38 : _GEN_1707; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1709 = 14'h23 == field_data_lo_18 ? _field_data_T_39 : _GEN_1708; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1710 = 14'h24 == field_data_lo_18 ? _field_data_T_40 : _GEN_1709; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1711 = 14'h25 == field_data_lo_18 ? _field_data_T_41 : _GEN_1710; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1712 = 14'h26 == field_data_lo_18 ? _field_data_T_42 : _GEN_1711; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1713 = 14'h27 == field_data_lo_18 ? _field_data_T_43 : _GEN_1712; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1714 = 14'h28 == field_data_lo_18 ? _field_data_T_44 : _GEN_1713; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1715 = 14'h29 == field_data_lo_18 ? _field_data_T_45 : _GEN_1714; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1716 = 14'h2a == field_data_lo_18 ? _field_data_T_46 : _GEN_1715; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1717 = 14'h2b == field_data_lo_18 ? _field_data_T_47 : _GEN_1716; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1718 = 14'h2c == field_data_lo_18 ? _field_data_T_48 : _GEN_1717; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1719 = 14'h2d == field_data_lo_18 ? _field_data_T_49 : _GEN_1718; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1720 = 14'h2e == field_data_lo_18 ? _field_data_T_50 : _GEN_1719; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1721 = 14'h2f == field_data_lo_18 ? _field_data_T_51 : _GEN_1720; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1722 = 14'h30 == field_data_lo_18 ? _field_data_T_52 : _GEN_1721; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1723 = 14'h31 == field_data_lo_18 ? _field_data_T_53 : _GEN_1722; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_39 = vliw_39[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_19 = vliw_39[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_39 = field_data_lo_19[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_39 = field_data_lo_19[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_58 = {{1'd0}, args_offset_39}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_58 = _total_offset_T_58[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1727 = 3'h1 == total_offset_58 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1728 = 3'h2 == total_offset_58 ? args_2 : _GEN_1727; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1729 = 3'h3 == total_offset_58 ? args_3 : _GEN_1728; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1730 = 3'h4 == total_offset_58 ? args_4 : _GEN_1729; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1731 = 3'h5 == total_offset_58 ? args_5 : _GEN_1730; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1732 = 3'h6 == total_offset_58 ? args_6 : _GEN_1731; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1733 = total_offset_58 < 3'h7 ? _GEN_1732 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_39_1 = 3'h0 < args_length_39 ? _GEN_1733 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_59 = args_offset_39 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1736 = 3'h1 == total_offset_59 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1737 = 3'h2 == total_offset_59 ? args_2 : _GEN_1736; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1738 = 3'h3 == total_offset_59 ? args_3 : _GEN_1737; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1739 = 3'h4 == total_offset_59 ? args_4 : _GEN_1738; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1740 = 3'h5 == total_offset_59 ? args_5 : _GEN_1739; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1741 = 3'h6 == total_offset_59 ? args_6 : _GEN_1740; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1742 = total_offset_59 < 3'h7 ? _GEN_1741 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_39_0 = 3'h1 < args_length_39 ? _GEN_1742 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_666 = {field_bytes_39_0,field_bytes_39_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1744 = opcode_39 == 4'ha ? _field_data_T_666 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1745 = opcode_39 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1286 = opcode_39 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_19 = field_data_lo_19[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_669 = {field_data_hi_19,field_data_lo_19}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_79 = _T_1286 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1746 = opcode_39 == 4'h8 | opcode_39 == 4'hb ? _field_data_T_669 : _GEN_1744; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1747 = opcode_39 == 4'h8 | opcode_39 == 4'hb ? _field_tag_T_79 : _GEN_1745; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1748 = 14'h14 == field_data_lo_19 ? _field_data_T_24 : _GEN_1746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1749 = 14'h15 == field_data_lo_19 ? _field_data_T_25 : _GEN_1748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1750 = 14'h16 == field_data_lo_19 ? _field_data_T_26 : _GEN_1749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1751 = 14'h17 == field_data_lo_19 ? _field_data_T_27 : _GEN_1750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1752 = 14'h18 == field_data_lo_19 ? _field_data_T_28 : _GEN_1751; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1753 = 14'h19 == field_data_lo_19 ? _field_data_T_29 : _GEN_1752; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1754 = 14'h1a == field_data_lo_19 ? _field_data_T_30 : _GEN_1753; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1755 = 14'h1b == field_data_lo_19 ? _field_data_T_31 : _GEN_1754; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1756 = 14'h1c == field_data_lo_19 ? _field_data_T_32 : _GEN_1755; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1757 = 14'h1d == field_data_lo_19 ? _field_data_T_33 : _GEN_1756; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1758 = 14'h1e == field_data_lo_19 ? _field_data_T_34 : _GEN_1757; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1759 = 14'h1f == field_data_lo_19 ? _field_data_T_35 : _GEN_1758; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1760 = 14'h20 == field_data_lo_19 ? _field_data_T_36 : _GEN_1759; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1761 = 14'h21 == field_data_lo_19 ? _field_data_T_37 : _GEN_1760; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1762 = 14'h22 == field_data_lo_19 ? _field_data_T_38 : _GEN_1761; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1763 = 14'h23 == field_data_lo_19 ? _field_data_T_39 : _GEN_1762; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1764 = 14'h24 == field_data_lo_19 ? _field_data_T_40 : _GEN_1763; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1765 = 14'h25 == field_data_lo_19 ? _field_data_T_41 : _GEN_1764; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1766 = 14'h26 == field_data_lo_19 ? _field_data_T_42 : _GEN_1765; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1767 = 14'h27 == field_data_lo_19 ? _field_data_T_43 : _GEN_1766; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1768 = 14'h28 == field_data_lo_19 ? _field_data_T_44 : _GEN_1767; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1769 = 14'h29 == field_data_lo_19 ? _field_data_T_45 : _GEN_1768; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1770 = 14'h2a == field_data_lo_19 ? _field_data_T_46 : _GEN_1769; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1771 = 14'h2b == field_data_lo_19 ? _field_data_T_47 : _GEN_1770; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1772 = 14'h2c == field_data_lo_19 ? _field_data_T_48 : _GEN_1771; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1773 = 14'h2d == field_data_lo_19 ? _field_data_T_49 : _GEN_1772; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1774 = 14'h2e == field_data_lo_19 ? _field_data_T_50 : _GEN_1773; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1775 = 14'h2f == field_data_lo_19 ? _field_data_T_51 : _GEN_1774; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1776 = 14'h30 == field_data_lo_19 ? _field_data_T_52 : _GEN_1775; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1777 = 14'h31 == field_data_lo_19 ? _field_data_T_53 : _GEN_1776; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_40 = vliw_40[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_20 = vliw_40[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_40 = field_data_lo_20[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_40 = field_data_lo_20[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_60 = {{1'd0}, args_offset_40}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_60 = _total_offset_T_60[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1781 = 3'h1 == total_offset_60 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1782 = 3'h2 == total_offset_60 ? args_2 : _GEN_1781; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1783 = 3'h3 == total_offset_60 ? args_3 : _GEN_1782; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1784 = 3'h4 == total_offset_60 ? args_4 : _GEN_1783; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1785 = 3'h5 == total_offset_60 ? args_5 : _GEN_1784; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1786 = 3'h6 == total_offset_60 ? args_6 : _GEN_1785; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1787 = total_offset_60 < 3'h7 ? _GEN_1786 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_40_1 = 3'h0 < args_length_40 ? _GEN_1787 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_61 = args_offset_40 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1790 = 3'h1 == total_offset_61 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1791 = 3'h2 == total_offset_61 ? args_2 : _GEN_1790; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1792 = 3'h3 == total_offset_61 ? args_3 : _GEN_1791; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1793 = 3'h4 == total_offset_61 ? args_4 : _GEN_1792; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1794 = 3'h5 == total_offset_61 ? args_5 : _GEN_1793; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1795 = 3'h6 == total_offset_61 ? args_6 : _GEN_1794; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1796 = total_offset_61 < 3'h7 ? _GEN_1795 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_40_0 = 3'h1 < args_length_40 ? _GEN_1796 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_700 = {field_bytes_40_0,field_bytes_40_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1798 = opcode_40 == 4'ha ? _field_data_T_700 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1799 = opcode_40 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1325 = opcode_40 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_20 = field_data_lo_20[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_703 = {field_data_hi_20,field_data_lo_20}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_81 = _T_1325 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1800 = opcode_40 == 4'h8 | opcode_40 == 4'hb ? _field_data_T_703 : _GEN_1798; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1801 = opcode_40 == 4'h8 | opcode_40 == 4'hb ? _field_tag_T_81 : _GEN_1799; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1802 = 14'h14 == field_data_lo_20 ? _field_data_T_24 : _GEN_1800; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1803 = 14'h15 == field_data_lo_20 ? _field_data_T_25 : _GEN_1802; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1804 = 14'h16 == field_data_lo_20 ? _field_data_T_26 : _GEN_1803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1805 = 14'h17 == field_data_lo_20 ? _field_data_T_27 : _GEN_1804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1806 = 14'h18 == field_data_lo_20 ? _field_data_T_28 : _GEN_1805; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1807 = 14'h19 == field_data_lo_20 ? _field_data_T_29 : _GEN_1806; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1808 = 14'h1a == field_data_lo_20 ? _field_data_T_30 : _GEN_1807; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1809 = 14'h1b == field_data_lo_20 ? _field_data_T_31 : _GEN_1808; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1810 = 14'h1c == field_data_lo_20 ? _field_data_T_32 : _GEN_1809; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1811 = 14'h1d == field_data_lo_20 ? _field_data_T_33 : _GEN_1810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1812 = 14'h1e == field_data_lo_20 ? _field_data_T_34 : _GEN_1811; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1813 = 14'h1f == field_data_lo_20 ? _field_data_T_35 : _GEN_1812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1814 = 14'h20 == field_data_lo_20 ? _field_data_T_36 : _GEN_1813; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1815 = 14'h21 == field_data_lo_20 ? _field_data_T_37 : _GEN_1814; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1816 = 14'h22 == field_data_lo_20 ? _field_data_T_38 : _GEN_1815; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1817 = 14'h23 == field_data_lo_20 ? _field_data_T_39 : _GEN_1816; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1818 = 14'h24 == field_data_lo_20 ? _field_data_T_40 : _GEN_1817; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1819 = 14'h25 == field_data_lo_20 ? _field_data_T_41 : _GEN_1818; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1820 = 14'h26 == field_data_lo_20 ? _field_data_T_42 : _GEN_1819; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1821 = 14'h27 == field_data_lo_20 ? _field_data_T_43 : _GEN_1820; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1822 = 14'h28 == field_data_lo_20 ? _field_data_T_44 : _GEN_1821; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1823 = 14'h29 == field_data_lo_20 ? _field_data_T_45 : _GEN_1822; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1824 = 14'h2a == field_data_lo_20 ? _field_data_T_46 : _GEN_1823; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1825 = 14'h2b == field_data_lo_20 ? _field_data_T_47 : _GEN_1824; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1826 = 14'h2c == field_data_lo_20 ? _field_data_T_48 : _GEN_1825; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1827 = 14'h2d == field_data_lo_20 ? _field_data_T_49 : _GEN_1826; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1828 = 14'h2e == field_data_lo_20 ? _field_data_T_50 : _GEN_1827; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1829 = 14'h2f == field_data_lo_20 ? _field_data_T_51 : _GEN_1828; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1830 = 14'h30 == field_data_lo_20 ? _field_data_T_52 : _GEN_1829; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1831 = 14'h31 == field_data_lo_20 ? _field_data_T_53 : _GEN_1830; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_41 = vliw_41[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_21 = vliw_41[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_41 = field_data_lo_21[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_41 = field_data_lo_21[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_62 = {{1'd0}, args_offset_41}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_62 = _total_offset_T_62[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1835 = 3'h1 == total_offset_62 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1836 = 3'h2 == total_offset_62 ? args_2 : _GEN_1835; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1837 = 3'h3 == total_offset_62 ? args_3 : _GEN_1836; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1838 = 3'h4 == total_offset_62 ? args_4 : _GEN_1837; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1839 = 3'h5 == total_offset_62 ? args_5 : _GEN_1838; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1840 = 3'h6 == total_offset_62 ? args_6 : _GEN_1839; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1841 = total_offset_62 < 3'h7 ? _GEN_1840 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_41_1 = 3'h0 < args_length_41 ? _GEN_1841 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_63 = args_offset_41 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1844 = 3'h1 == total_offset_63 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1845 = 3'h2 == total_offset_63 ? args_2 : _GEN_1844; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1846 = 3'h3 == total_offset_63 ? args_3 : _GEN_1845; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1847 = 3'h4 == total_offset_63 ? args_4 : _GEN_1846; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1848 = 3'h5 == total_offset_63 ? args_5 : _GEN_1847; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1849 = 3'h6 == total_offset_63 ? args_6 : _GEN_1848; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1850 = total_offset_63 < 3'h7 ? _GEN_1849 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_41_0 = 3'h1 < args_length_41 ? _GEN_1850 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_734 = {field_bytes_41_0,field_bytes_41_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1852 = opcode_41 == 4'ha ? _field_data_T_734 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1853 = opcode_41 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1364 = opcode_41 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_21 = field_data_lo_21[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_737 = {field_data_hi_21,field_data_lo_21}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_83 = _T_1364 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1854 = opcode_41 == 4'h8 | opcode_41 == 4'hb ? _field_data_T_737 : _GEN_1852; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1855 = opcode_41 == 4'h8 | opcode_41 == 4'hb ? _field_tag_T_83 : _GEN_1853; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1856 = 14'h14 == field_data_lo_21 ? _field_data_T_24 : _GEN_1854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1857 = 14'h15 == field_data_lo_21 ? _field_data_T_25 : _GEN_1856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1858 = 14'h16 == field_data_lo_21 ? _field_data_T_26 : _GEN_1857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1859 = 14'h17 == field_data_lo_21 ? _field_data_T_27 : _GEN_1858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1860 = 14'h18 == field_data_lo_21 ? _field_data_T_28 : _GEN_1859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1861 = 14'h19 == field_data_lo_21 ? _field_data_T_29 : _GEN_1860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1862 = 14'h1a == field_data_lo_21 ? _field_data_T_30 : _GEN_1861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1863 = 14'h1b == field_data_lo_21 ? _field_data_T_31 : _GEN_1862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1864 = 14'h1c == field_data_lo_21 ? _field_data_T_32 : _GEN_1863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1865 = 14'h1d == field_data_lo_21 ? _field_data_T_33 : _GEN_1864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1866 = 14'h1e == field_data_lo_21 ? _field_data_T_34 : _GEN_1865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1867 = 14'h1f == field_data_lo_21 ? _field_data_T_35 : _GEN_1866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1868 = 14'h20 == field_data_lo_21 ? _field_data_T_36 : _GEN_1867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1869 = 14'h21 == field_data_lo_21 ? _field_data_T_37 : _GEN_1868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1870 = 14'h22 == field_data_lo_21 ? _field_data_T_38 : _GEN_1869; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1871 = 14'h23 == field_data_lo_21 ? _field_data_T_39 : _GEN_1870; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1872 = 14'h24 == field_data_lo_21 ? _field_data_T_40 : _GEN_1871; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1873 = 14'h25 == field_data_lo_21 ? _field_data_T_41 : _GEN_1872; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1874 = 14'h26 == field_data_lo_21 ? _field_data_T_42 : _GEN_1873; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1875 = 14'h27 == field_data_lo_21 ? _field_data_T_43 : _GEN_1874; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1876 = 14'h28 == field_data_lo_21 ? _field_data_T_44 : _GEN_1875; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1877 = 14'h29 == field_data_lo_21 ? _field_data_T_45 : _GEN_1876; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1878 = 14'h2a == field_data_lo_21 ? _field_data_T_46 : _GEN_1877; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1879 = 14'h2b == field_data_lo_21 ? _field_data_T_47 : _GEN_1878; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1880 = 14'h2c == field_data_lo_21 ? _field_data_T_48 : _GEN_1879; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1881 = 14'h2d == field_data_lo_21 ? _field_data_T_49 : _GEN_1880; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1882 = 14'h2e == field_data_lo_21 ? _field_data_T_50 : _GEN_1881; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1883 = 14'h2f == field_data_lo_21 ? _field_data_T_51 : _GEN_1882; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1884 = 14'h30 == field_data_lo_21 ? _field_data_T_52 : _GEN_1883; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1885 = 14'h31 == field_data_lo_21 ? _field_data_T_53 : _GEN_1884; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_42 = vliw_42[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_22 = vliw_42[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_42 = field_data_lo_22[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_42 = field_data_lo_22[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_64 = {{1'd0}, args_offset_42}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_64 = _total_offset_T_64[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1889 = 3'h1 == total_offset_64 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1890 = 3'h2 == total_offset_64 ? args_2 : _GEN_1889; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1891 = 3'h3 == total_offset_64 ? args_3 : _GEN_1890; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1892 = 3'h4 == total_offset_64 ? args_4 : _GEN_1891; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1893 = 3'h5 == total_offset_64 ? args_5 : _GEN_1892; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1894 = 3'h6 == total_offset_64 ? args_6 : _GEN_1893; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1895 = total_offset_64 < 3'h7 ? _GEN_1894 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_42_1 = 3'h0 < args_length_42 ? _GEN_1895 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_65 = args_offset_42 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1898 = 3'h1 == total_offset_65 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1899 = 3'h2 == total_offset_65 ? args_2 : _GEN_1898; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1900 = 3'h3 == total_offset_65 ? args_3 : _GEN_1899; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1901 = 3'h4 == total_offset_65 ? args_4 : _GEN_1900; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1902 = 3'h5 == total_offset_65 ? args_5 : _GEN_1901; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1903 = 3'h6 == total_offset_65 ? args_6 : _GEN_1902; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1904 = total_offset_65 < 3'h7 ? _GEN_1903 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_42_0 = 3'h1 < args_length_42 ? _GEN_1904 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_768 = {field_bytes_42_0,field_bytes_42_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1906 = opcode_42 == 4'ha ? _field_data_T_768 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1907 = opcode_42 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1403 = opcode_42 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_22 = field_data_lo_22[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_771 = {field_data_hi_22,field_data_lo_22}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_85 = _T_1403 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1908 = opcode_42 == 4'h8 | opcode_42 == 4'hb ? _field_data_T_771 : _GEN_1906; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1909 = opcode_42 == 4'h8 | opcode_42 == 4'hb ? _field_tag_T_85 : _GEN_1907; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1910 = 14'h14 == field_data_lo_22 ? _field_data_T_24 : _GEN_1908; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1911 = 14'h15 == field_data_lo_22 ? _field_data_T_25 : _GEN_1910; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1912 = 14'h16 == field_data_lo_22 ? _field_data_T_26 : _GEN_1911; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1913 = 14'h17 == field_data_lo_22 ? _field_data_T_27 : _GEN_1912; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1914 = 14'h18 == field_data_lo_22 ? _field_data_T_28 : _GEN_1913; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1915 = 14'h19 == field_data_lo_22 ? _field_data_T_29 : _GEN_1914; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1916 = 14'h1a == field_data_lo_22 ? _field_data_T_30 : _GEN_1915; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1917 = 14'h1b == field_data_lo_22 ? _field_data_T_31 : _GEN_1916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1918 = 14'h1c == field_data_lo_22 ? _field_data_T_32 : _GEN_1917; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1919 = 14'h1d == field_data_lo_22 ? _field_data_T_33 : _GEN_1918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1920 = 14'h1e == field_data_lo_22 ? _field_data_T_34 : _GEN_1919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1921 = 14'h1f == field_data_lo_22 ? _field_data_T_35 : _GEN_1920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1922 = 14'h20 == field_data_lo_22 ? _field_data_T_36 : _GEN_1921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1923 = 14'h21 == field_data_lo_22 ? _field_data_T_37 : _GEN_1922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1924 = 14'h22 == field_data_lo_22 ? _field_data_T_38 : _GEN_1923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1925 = 14'h23 == field_data_lo_22 ? _field_data_T_39 : _GEN_1924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1926 = 14'h24 == field_data_lo_22 ? _field_data_T_40 : _GEN_1925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1927 = 14'h25 == field_data_lo_22 ? _field_data_T_41 : _GEN_1926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1928 = 14'h26 == field_data_lo_22 ? _field_data_T_42 : _GEN_1927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1929 = 14'h27 == field_data_lo_22 ? _field_data_T_43 : _GEN_1928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1930 = 14'h28 == field_data_lo_22 ? _field_data_T_44 : _GEN_1929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1931 = 14'h29 == field_data_lo_22 ? _field_data_T_45 : _GEN_1930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1932 = 14'h2a == field_data_lo_22 ? _field_data_T_46 : _GEN_1931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1933 = 14'h2b == field_data_lo_22 ? _field_data_T_47 : _GEN_1932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1934 = 14'h2c == field_data_lo_22 ? _field_data_T_48 : _GEN_1933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1935 = 14'h2d == field_data_lo_22 ? _field_data_T_49 : _GEN_1934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1936 = 14'h2e == field_data_lo_22 ? _field_data_T_50 : _GEN_1935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1937 = 14'h2f == field_data_lo_22 ? _field_data_T_51 : _GEN_1936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1938 = 14'h30 == field_data_lo_22 ? _field_data_T_52 : _GEN_1937; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1939 = 14'h31 == field_data_lo_22 ? _field_data_T_53 : _GEN_1938; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_43 = vliw_43[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_23 = vliw_43[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_43 = field_data_lo_23[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_43 = field_data_lo_23[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_66 = {{1'd0}, args_offset_43}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_66 = _total_offset_T_66[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1943 = 3'h1 == total_offset_66 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1944 = 3'h2 == total_offset_66 ? args_2 : _GEN_1943; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1945 = 3'h3 == total_offset_66 ? args_3 : _GEN_1944; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1946 = 3'h4 == total_offset_66 ? args_4 : _GEN_1945; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1947 = 3'h5 == total_offset_66 ? args_5 : _GEN_1946; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1948 = 3'h6 == total_offset_66 ? args_6 : _GEN_1947; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1949 = total_offset_66 < 3'h7 ? _GEN_1948 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_43_1 = 3'h0 < args_length_43 ? _GEN_1949 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_67 = args_offset_43 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1952 = 3'h1 == total_offset_67 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1953 = 3'h2 == total_offset_67 ? args_2 : _GEN_1952; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1954 = 3'h3 == total_offset_67 ? args_3 : _GEN_1953; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1955 = 3'h4 == total_offset_67 ? args_4 : _GEN_1954; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1956 = 3'h5 == total_offset_67 ? args_5 : _GEN_1955; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1957 = 3'h6 == total_offset_67 ? args_6 : _GEN_1956; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1958 = total_offset_67 < 3'h7 ? _GEN_1957 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_43_0 = 3'h1 < args_length_43 ? _GEN_1958 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_802 = {field_bytes_43_0,field_bytes_43_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_1960 = opcode_43 == 4'ha ? _field_data_T_802 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_1961 = opcode_43 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1442 = opcode_43 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_23 = field_data_lo_23[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_805 = {field_data_hi_23,field_data_lo_23}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_87 = _T_1442 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_1962 = opcode_43 == 4'h8 | opcode_43 == 4'hb ? _field_data_T_805 : _GEN_1960; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_1963 = opcode_43 == 4'h8 | opcode_43 == 4'hb ? _field_tag_T_87 : _GEN_1961; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_1964 = 14'h14 == field_data_lo_23 ? _field_data_T_24 : _GEN_1962; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1965 = 14'h15 == field_data_lo_23 ? _field_data_T_25 : _GEN_1964; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1966 = 14'h16 == field_data_lo_23 ? _field_data_T_26 : _GEN_1965; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1967 = 14'h17 == field_data_lo_23 ? _field_data_T_27 : _GEN_1966; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1968 = 14'h18 == field_data_lo_23 ? _field_data_T_28 : _GEN_1967; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1969 = 14'h19 == field_data_lo_23 ? _field_data_T_29 : _GEN_1968; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1970 = 14'h1a == field_data_lo_23 ? _field_data_T_30 : _GEN_1969; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1971 = 14'h1b == field_data_lo_23 ? _field_data_T_31 : _GEN_1970; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1972 = 14'h1c == field_data_lo_23 ? _field_data_T_32 : _GEN_1971; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1973 = 14'h1d == field_data_lo_23 ? _field_data_T_33 : _GEN_1972; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1974 = 14'h1e == field_data_lo_23 ? _field_data_T_34 : _GEN_1973; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1975 = 14'h1f == field_data_lo_23 ? _field_data_T_35 : _GEN_1974; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1976 = 14'h20 == field_data_lo_23 ? _field_data_T_36 : _GEN_1975; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1977 = 14'h21 == field_data_lo_23 ? _field_data_T_37 : _GEN_1976; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1978 = 14'h22 == field_data_lo_23 ? _field_data_T_38 : _GEN_1977; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1979 = 14'h23 == field_data_lo_23 ? _field_data_T_39 : _GEN_1978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1980 = 14'h24 == field_data_lo_23 ? _field_data_T_40 : _GEN_1979; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1981 = 14'h25 == field_data_lo_23 ? _field_data_T_41 : _GEN_1980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1982 = 14'h26 == field_data_lo_23 ? _field_data_T_42 : _GEN_1981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1983 = 14'h27 == field_data_lo_23 ? _field_data_T_43 : _GEN_1982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1984 = 14'h28 == field_data_lo_23 ? _field_data_T_44 : _GEN_1983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1985 = 14'h29 == field_data_lo_23 ? _field_data_T_45 : _GEN_1984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1986 = 14'h2a == field_data_lo_23 ? _field_data_T_46 : _GEN_1985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1987 = 14'h2b == field_data_lo_23 ? _field_data_T_47 : _GEN_1986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1988 = 14'h2c == field_data_lo_23 ? _field_data_T_48 : _GEN_1987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1989 = 14'h2d == field_data_lo_23 ? _field_data_T_49 : _GEN_1988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1990 = 14'h2e == field_data_lo_23 ? _field_data_T_50 : _GEN_1989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1991 = 14'h2f == field_data_lo_23 ? _field_data_T_51 : _GEN_1990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1992 = 14'h30 == field_data_lo_23 ? _field_data_T_52 : _GEN_1991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_1993 = 14'h31 == field_data_lo_23 ? _field_data_T_53 : _GEN_1992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_44 = vliw_44[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_24 = vliw_44[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_44 = field_data_lo_24[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_44 = field_data_lo_24[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_68 = {{1'd0}, args_offset_44}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_68 = _total_offset_T_68[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_1997 = 3'h1 == total_offset_68 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1998 = 3'h2 == total_offset_68 ? args_2 : _GEN_1997; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_1999 = 3'h3 == total_offset_68 ? args_3 : _GEN_1998; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2000 = 3'h4 == total_offset_68 ? args_4 : _GEN_1999; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2001 = 3'h5 == total_offset_68 ? args_5 : _GEN_2000; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2002 = 3'h6 == total_offset_68 ? args_6 : _GEN_2001; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2003 = total_offset_68 < 3'h7 ? _GEN_2002 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_44_1 = 3'h0 < args_length_44 ? _GEN_2003 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_69 = args_offset_44 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2006 = 3'h1 == total_offset_69 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2007 = 3'h2 == total_offset_69 ? args_2 : _GEN_2006; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2008 = 3'h3 == total_offset_69 ? args_3 : _GEN_2007; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2009 = 3'h4 == total_offset_69 ? args_4 : _GEN_2008; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2010 = 3'h5 == total_offset_69 ? args_5 : _GEN_2009; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2011 = 3'h6 == total_offset_69 ? args_6 : _GEN_2010; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2012 = total_offset_69 < 3'h7 ? _GEN_2011 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_44_0 = 3'h1 < args_length_44 ? _GEN_2012 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_836 = {field_bytes_44_0,field_bytes_44_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2014 = opcode_44 == 4'ha ? _field_data_T_836 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2015 = opcode_44 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1481 = opcode_44 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_24 = field_data_lo_24[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_839 = {field_data_hi_24,field_data_lo_24}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_89 = _T_1481 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2016 = opcode_44 == 4'h8 | opcode_44 == 4'hb ? _field_data_T_839 : _GEN_2014; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2017 = opcode_44 == 4'h8 | opcode_44 == 4'hb ? _field_tag_T_89 : _GEN_2015; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2018 = 14'h14 == field_data_lo_24 ? _field_data_T_24 : _GEN_2016; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2019 = 14'h15 == field_data_lo_24 ? _field_data_T_25 : _GEN_2018; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2020 = 14'h16 == field_data_lo_24 ? _field_data_T_26 : _GEN_2019; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2021 = 14'h17 == field_data_lo_24 ? _field_data_T_27 : _GEN_2020; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2022 = 14'h18 == field_data_lo_24 ? _field_data_T_28 : _GEN_2021; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2023 = 14'h19 == field_data_lo_24 ? _field_data_T_29 : _GEN_2022; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2024 = 14'h1a == field_data_lo_24 ? _field_data_T_30 : _GEN_2023; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2025 = 14'h1b == field_data_lo_24 ? _field_data_T_31 : _GEN_2024; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2026 = 14'h1c == field_data_lo_24 ? _field_data_T_32 : _GEN_2025; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2027 = 14'h1d == field_data_lo_24 ? _field_data_T_33 : _GEN_2026; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2028 = 14'h1e == field_data_lo_24 ? _field_data_T_34 : _GEN_2027; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2029 = 14'h1f == field_data_lo_24 ? _field_data_T_35 : _GEN_2028; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2030 = 14'h20 == field_data_lo_24 ? _field_data_T_36 : _GEN_2029; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2031 = 14'h21 == field_data_lo_24 ? _field_data_T_37 : _GEN_2030; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2032 = 14'h22 == field_data_lo_24 ? _field_data_T_38 : _GEN_2031; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2033 = 14'h23 == field_data_lo_24 ? _field_data_T_39 : _GEN_2032; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2034 = 14'h24 == field_data_lo_24 ? _field_data_T_40 : _GEN_2033; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2035 = 14'h25 == field_data_lo_24 ? _field_data_T_41 : _GEN_2034; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2036 = 14'h26 == field_data_lo_24 ? _field_data_T_42 : _GEN_2035; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2037 = 14'h27 == field_data_lo_24 ? _field_data_T_43 : _GEN_2036; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2038 = 14'h28 == field_data_lo_24 ? _field_data_T_44 : _GEN_2037; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2039 = 14'h29 == field_data_lo_24 ? _field_data_T_45 : _GEN_2038; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2040 = 14'h2a == field_data_lo_24 ? _field_data_T_46 : _GEN_2039; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2041 = 14'h2b == field_data_lo_24 ? _field_data_T_47 : _GEN_2040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2042 = 14'h2c == field_data_lo_24 ? _field_data_T_48 : _GEN_2041; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2043 = 14'h2d == field_data_lo_24 ? _field_data_T_49 : _GEN_2042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2044 = 14'h2e == field_data_lo_24 ? _field_data_T_50 : _GEN_2043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2045 = 14'h2f == field_data_lo_24 ? _field_data_T_51 : _GEN_2044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2046 = 14'h30 == field_data_lo_24 ? _field_data_T_52 : _GEN_2045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2047 = 14'h31 == field_data_lo_24 ? _field_data_T_53 : _GEN_2046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_45 = vliw_45[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_25 = vliw_45[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_45 = field_data_lo_25[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_45 = field_data_lo_25[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_70 = {{1'd0}, args_offset_45}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_70 = _total_offset_T_70[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2051 = 3'h1 == total_offset_70 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2052 = 3'h2 == total_offset_70 ? args_2 : _GEN_2051; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2053 = 3'h3 == total_offset_70 ? args_3 : _GEN_2052; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2054 = 3'h4 == total_offset_70 ? args_4 : _GEN_2053; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2055 = 3'h5 == total_offset_70 ? args_5 : _GEN_2054; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2056 = 3'h6 == total_offset_70 ? args_6 : _GEN_2055; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2057 = total_offset_70 < 3'h7 ? _GEN_2056 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_45_1 = 3'h0 < args_length_45 ? _GEN_2057 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_71 = args_offset_45 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2060 = 3'h1 == total_offset_71 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2061 = 3'h2 == total_offset_71 ? args_2 : _GEN_2060; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2062 = 3'h3 == total_offset_71 ? args_3 : _GEN_2061; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2063 = 3'h4 == total_offset_71 ? args_4 : _GEN_2062; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2064 = 3'h5 == total_offset_71 ? args_5 : _GEN_2063; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2065 = 3'h6 == total_offset_71 ? args_6 : _GEN_2064; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2066 = total_offset_71 < 3'h7 ? _GEN_2065 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_45_0 = 3'h1 < args_length_45 ? _GEN_2066 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_870 = {field_bytes_45_0,field_bytes_45_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2068 = opcode_45 == 4'ha ? _field_data_T_870 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2069 = opcode_45 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1520 = opcode_45 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_25 = field_data_lo_25[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_873 = {field_data_hi_25,field_data_lo_25}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_91 = _T_1520 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2070 = opcode_45 == 4'h8 | opcode_45 == 4'hb ? _field_data_T_873 : _GEN_2068; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2071 = opcode_45 == 4'h8 | opcode_45 == 4'hb ? _field_tag_T_91 : _GEN_2069; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2072 = 14'h14 == field_data_lo_25 ? _field_data_T_24 : _GEN_2070; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2073 = 14'h15 == field_data_lo_25 ? _field_data_T_25 : _GEN_2072; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2074 = 14'h16 == field_data_lo_25 ? _field_data_T_26 : _GEN_2073; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2075 = 14'h17 == field_data_lo_25 ? _field_data_T_27 : _GEN_2074; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2076 = 14'h18 == field_data_lo_25 ? _field_data_T_28 : _GEN_2075; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2077 = 14'h19 == field_data_lo_25 ? _field_data_T_29 : _GEN_2076; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2078 = 14'h1a == field_data_lo_25 ? _field_data_T_30 : _GEN_2077; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2079 = 14'h1b == field_data_lo_25 ? _field_data_T_31 : _GEN_2078; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2080 = 14'h1c == field_data_lo_25 ? _field_data_T_32 : _GEN_2079; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2081 = 14'h1d == field_data_lo_25 ? _field_data_T_33 : _GEN_2080; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2082 = 14'h1e == field_data_lo_25 ? _field_data_T_34 : _GEN_2081; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2083 = 14'h1f == field_data_lo_25 ? _field_data_T_35 : _GEN_2082; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2084 = 14'h20 == field_data_lo_25 ? _field_data_T_36 : _GEN_2083; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2085 = 14'h21 == field_data_lo_25 ? _field_data_T_37 : _GEN_2084; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2086 = 14'h22 == field_data_lo_25 ? _field_data_T_38 : _GEN_2085; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2087 = 14'h23 == field_data_lo_25 ? _field_data_T_39 : _GEN_2086; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2088 = 14'h24 == field_data_lo_25 ? _field_data_T_40 : _GEN_2087; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2089 = 14'h25 == field_data_lo_25 ? _field_data_T_41 : _GEN_2088; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2090 = 14'h26 == field_data_lo_25 ? _field_data_T_42 : _GEN_2089; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2091 = 14'h27 == field_data_lo_25 ? _field_data_T_43 : _GEN_2090; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2092 = 14'h28 == field_data_lo_25 ? _field_data_T_44 : _GEN_2091; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2093 = 14'h29 == field_data_lo_25 ? _field_data_T_45 : _GEN_2092; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2094 = 14'h2a == field_data_lo_25 ? _field_data_T_46 : _GEN_2093; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2095 = 14'h2b == field_data_lo_25 ? _field_data_T_47 : _GEN_2094; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2096 = 14'h2c == field_data_lo_25 ? _field_data_T_48 : _GEN_2095; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2097 = 14'h2d == field_data_lo_25 ? _field_data_T_49 : _GEN_2096; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2098 = 14'h2e == field_data_lo_25 ? _field_data_T_50 : _GEN_2097; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2099 = 14'h2f == field_data_lo_25 ? _field_data_T_51 : _GEN_2098; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2100 = 14'h30 == field_data_lo_25 ? _field_data_T_52 : _GEN_2099; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2101 = 14'h31 == field_data_lo_25 ? _field_data_T_53 : _GEN_2100; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_46 = vliw_46[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_26 = vliw_46[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_46 = field_data_lo_26[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_46 = field_data_lo_26[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_72 = {{1'd0}, args_offset_46}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_72 = _total_offset_T_72[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2105 = 3'h1 == total_offset_72 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2106 = 3'h2 == total_offset_72 ? args_2 : _GEN_2105; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2107 = 3'h3 == total_offset_72 ? args_3 : _GEN_2106; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2108 = 3'h4 == total_offset_72 ? args_4 : _GEN_2107; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2109 = 3'h5 == total_offset_72 ? args_5 : _GEN_2108; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2110 = 3'h6 == total_offset_72 ? args_6 : _GEN_2109; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2111 = total_offset_72 < 3'h7 ? _GEN_2110 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_46_1 = 3'h0 < args_length_46 ? _GEN_2111 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_73 = args_offset_46 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2114 = 3'h1 == total_offset_73 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2115 = 3'h2 == total_offset_73 ? args_2 : _GEN_2114; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2116 = 3'h3 == total_offset_73 ? args_3 : _GEN_2115; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2117 = 3'h4 == total_offset_73 ? args_4 : _GEN_2116; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2118 = 3'h5 == total_offset_73 ? args_5 : _GEN_2117; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2119 = 3'h6 == total_offset_73 ? args_6 : _GEN_2118; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2120 = total_offset_73 < 3'h7 ? _GEN_2119 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_46_0 = 3'h1 < args_length_46 ? _GEN_2120 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_904 = {field_bytes_46_0,field_bytes_46_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2122 = opcode_46 == 4'ha ? _field_data_T_904 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2123 = opcode_46 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1559 = opcode_46 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_26 = field_data_lo_26[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_907 = {field_data_hi_26,field_data_lo_26}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_93 = _T_1559 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2124 = opcode_46 == 4'h8 | opcode_46 == 4'hb ? _field_data_T_907 : _GEN_2122; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2125 = opcode_46 == 4'h8 | opcode_46 == 4'hb ? _field_tag_T_93 : _GEN_2123; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2126 = 14'h14 == field_data_lo_26 ? _field_data_T_24 : _GEN_2124; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2127 = 14'h15 == field_data_lo_26 ? _field_data_T_25 : _GEN_2126; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2128 = 14'h16 == field_data_lo_26 ? _field_data_T_26 : _GEN_2127; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2129 = 14'h17 == field_data_lo_26 ? _field_data_T_27 : _GEN_2128; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2130 = 14'h18 == field_data_lo_26 ? _field_data_T_28 : _GEN_2129; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2131 = 14'h19 == field_data_lo_26 ? _field_data_T_29 : _GEN_2130; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2132 = 14'h1a == field_data_lo_26 ? _field_data_T_30 : _GEN_2131; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2133 = 14'h1b == field_data_lo_26 ? _field_data_T_31 : _GEN_2132; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2134 = 14'h1c == field_data_lo_26 ? _field_data_T_32 : _GEN_2133; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2135 = 14'h1d == field_data_lo_26 ? _field_data_T_33 : _GEN_2134; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2136 = 14'h1e == field_data_lo_26 ? _field_data_T_34 : _GEN_2135; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2137 = 14'h1f == field_data_lo_26 ? _field_data_T_35 : _GEN_2136; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2138 = 14'h20 == field_data_lo_26 ? _field_data_T_36 : _GEN_2137; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2139 = 14'h21 == field_data_lo_26 ? _field_data_T_37 : _GEN_2138; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2140 = 14'h22 == field_data_lo_26 ? _field_data_T_38 : _GEN_2139; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2141 = 14'h23 == field_data_lo_26 ? _field_data_T_39 : _GEN_2140; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2142 = 14'h24 == field_data_lo_26 ? _field_data_T_40 : _GEN_2141; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2143 = 14'h25 == field_data_lo_26 ? _field_data_T_41 : _GEN_2142; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2144 = 14'h26 == field_data_lo_26 ? _field_data_T_42 : _GEN_2143; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2145 = 14'h27 == field_data_lo_26 ? _field_data_T_43 : _GEN_2144; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2146 = 14'h28 == field_data_lo_26 ? _field_data_T_44 : _GEN_2145; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2147 = 14'h29 == field_data_lo_26 ? _field_data_T_45 : _GEN_2146; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2148 = 14'h2a == field_data_lo_26 ? _field_data_T_46 : _GEN_2147; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2149 = 14'h2b == field_data_lo_26 ? _field_data_T_47 : _GEN_2148; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2150 = 14'h2c == field_data_lo_26 ? _field_data_T_48 : _GEN_2149; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2151 = 14'h2d == field_data_lo_26 ? _field_data_T_49 : _GEN_2150; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2152 = 14'h2e == field_data_lo_26 ? _field_data_T_50 : _GEN_2151; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2153 = 14'h2f == field_data_lo_26 ? _field_data_T_51 : _GEN_2152; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2154 = 14'h30 == field_data_lo_26 ? _field_data_T_52 : _GEN_2153; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2155 = 14'h31 == field_data_lo_26 ? _field_data_T_53 : _GEN_2154; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_47 = vliw_47[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_27 = vliw_47[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_47 = field_data_lo_27[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_47 = field_data_lo_27[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_74 = {{1'd0}, args_offset_47}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_74 = _total_offset_T_74[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2159 = 3'h1 == total_offset_74 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2160 = 3'h2 == total_offset_74 ? args_2 : _GEN_2159; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2161 = 3'h3 == total_offset_74 ? args_3 : _GEN_2160; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2162 = 3'h4 == total_offset_74 ? args_4 : _GEN_2161; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2163 = 3'h5 == total_offset_74 ? args_5 : _GEN_2162; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2164 = 3'h6 == total_offset_74 ? args_6 : _GEN_2163; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2165 = total_offset_74 < 3'h7 ? _GEN_2164 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_47_1 = 3'h0 < args_length_47 ? _GEN_2165 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_75 = args_offset_47 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2168 = 3'h1 == total_offset_75 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2169 = 3'h2 == total_offset_75 ? args_2 : _GEN_2168; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2170 = 3'h3 == total_offset_75 ? args_3 : _GEN_2169; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2171 = 3'h4 == total_offset_75 ? args_4 : _GEN_2170; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2172 = 3'h5 == total_offset_75 ? args_5 : _GEN_2171; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2173 = 3'h6 == total_offset_75 ? args_6 : _GEN_2172; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2174 = total_offset_75 < 3'h7 ? _GEN_2173 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_47_0 = 3'h1 < args_length_47 ? _GEN_2174 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_938 = {field_bytes_47_0,field_bytes_47_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2176 = opcode_47 == 4'ha ? _field_data_T_938 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2177 = opcode_47 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1598 = opcode_47 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_27 = field_data_lo_27[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_941 = {field_data_hi_27,field_data_lo_27}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_95 = _T_1598 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2178 = opcode_47 == 4'h8 | opcode_47 == 4'hb ? _field_data_T_941 : _GEN_2176; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2179 = opcode_47 == 4'h8 | opcode_47 == 4'hb ? _field_tag_T_95 : _GEN_2177; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2180 = 14'h14 == field_data_lo_27 ? _field_data_T_24 : _GEN_2178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2181 = 14'h15 == field_data_lo_27 ? _field_data_T_25 : _GEN_2180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2182 = 14'h16 == field_data_lo_27 ? _field_data_T_26 : _GEN_2181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2183 = 14'h17 == field_data_lo_27 ? _field_data_T_27 : _GEN_2182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2184 = 14'h18 == field_data_lo_27 ? _field_data_T_28 : _GEN_2183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2185 = 14'h19 == field_data_lo_27 ? _field_data_T_29 : _GEN_2184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2186 = 14'h1a == field_data_lo_27 ? _field_data_T_30 : _GEN_2185; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2187 = 14'h1b == field_data_lo_27 ? _field_data_T_31 : _GEN_2186; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2188 = 14'h1c == field_data_lo_27 ? _field_data_T_32 : _GEN_2187; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2189 = 14'h1d == field_data_lo_27 ? _field_data_T_33 : _GEN_2188; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2190 = 14'h1e == field_data_lo_27 ? _field_data_T_34 : _GEN_2189; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2191 = 14'h1f == field_data_lo_27 ? _field_data_T_35 : _GEN_2190; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2192 = 14'h20 == field_data_lo_27 ? _field_data_T_36 : _GEN_2191; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2193 = 14'h21 == field_data_lo_27 ? _field_data_T_37 : _GEN_2192; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2194 = 14'h22 == field_data_lo_27 ? _field_data_T_38 : _GEN_2193; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2195 = 14'h23 == field_data_lo_27 ? _field_data_T_39 : _GEN_2194; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2196 = 14'h24 == field_data_lo_27 ? _field_data_T_40 : _GEN_2195; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2197 = 14'h25 == field_data_lo_27 ? _field_data_T_41 : _GEN_2196; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2198 = 14'h26 == field_data_lo_27 ? _field_data_T_42 : _GEN_2197; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2199 = 14'h27 == field_data_lo_27 ? _field_data_T_43 : _GEN_2198; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2200 = 14'h28 == field_data_lo_27 ? _field_data_T_44 : _GEN_2199; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2201 = 14'h29 == field_data_lo_27 ? _field_data_T_45 : _GEN_2200; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2202 = 14'h2a == field_data_lo_27 ? _field_data_T_46 : _GEN_2201; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2203 = 14'h2b == field_data_lo_27 ? _field_data_T_47 : _GEN_2202; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2204 = 14'h2c == field_data_lo_27 ? _field_data_T_48 : _GEN_2203; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2205 = 14'h2d == field_data_lo_27 ? _field_data_T_49 : _GEN_2204; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2206 = 14'h2e == field_data_lo_27 ? _field_data_T_50 : _GEN_2205; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2207 = 14'h2f == field_data_lo_27 ? _field_data_T_51 : _GEN_2206; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2208 = 14'h30 == field_data_lo_27 ? _field_data_T_52 : _GEN_2207; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2209 = 14'h31 == field_data_lo_27 ? _field_data_T_53 : _GEN_2208; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_48 = vliw_48[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_28 = vliw_48[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_48 = field_data_lo_28[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_48 = field_data_lo_28[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_76 = {{1'd0}, args_offset_48}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_76 = _total_offset_T_76[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2213 = 3'h1 == total_offset_76 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2214 = 3'h2 == total_offset_76 ? args_2 : _GEN_2213; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2215 = 3'h3 == total_offset_76 ? args_3 : _GEN_2214; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2216 = 3'h4 == total_offset_76 ? args_4 : _GEN_2215; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2217 = 3'h5 == total_offset_76 ? args_5 : _GEN_2216; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2218 = 3'h6 == total_offset_76 ? args_6 : _GEN_2217; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2219 = total_offset_76 < 3'h7 ? _GEN_2218 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_48_1 = 3'h0 < args_length_48 ? _GEN_2219 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_77 = args_offset_48 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2222 = 3'h1 == total_offset_77 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2223 = 3'h2 == total_offset_77 ? args_2 : _GEN_2222; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2224 = 3'h3 == total_offset_77 ? args_3 : _GEN_2223; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2225 = 3'h4 == total_offset_77 ? args_4 : _GEN_2224; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2226 = 3'h5 == total_offset_77 ? args_5 : _GEN_2225; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2227 = 3'h6 == total_offset_77 ? args_6 : _GEN_2226; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2228 = total_offset_77 < 3'h7 ? _GEN_2227 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_48_0 = 3'h1 < args_length_48 ? _GEN_2228 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_972 = {field_bytes_48_0,field_bytes_48_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2230 = opcode_48 == 4'ha ? _field_data_T_972 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2231 = opcode_48 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1637 = opcode_48 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_28 = field_data_lo_28[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_975 = {field_data_hi_28,field_data_lo_28}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_97 = _T_1637 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2232 = opcode_48 == 4'h8 | opcode_48 == 4'hb ? _field_data_T_975 : _GEN_2230; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2233 = opcode_48 == 4'h8 | opcode_48 == 4'hb ? _field_tag_T_97 : _GEN_2231; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2234 = 14'h14 == field_data_lo_28 ? _field_data_T_24 : _GEN_2232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2235 = 14'h15 == field_data_lo_28 ? _field_data_T_25 : _GEN_2234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2236 = 14'h16 == field_data_lo_28 ? _field_data_T_26 : _GEN_2235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2237 = 14'h17 == field_data_lo_28 ? _field_data_T_27 : _GEN_2236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2238 = 14'h18 == field_data_lo_28 ? _field_data_T_28 : _GEN_2237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2239 = 14'h19 == field_data_lo_28 ? _field_data_T_29 : _GEN_2238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2240 = 14'h1a == field_data_lo_28 ? _field_data_T_30 : _GEN_2239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2241 = 14'h1b == field_data_lo_28 ? _field_data_T_31 : _GEN_2240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2242 = 14'h1c == field_data_lo_28 ? _field_data_T_32 : _GEN_2241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2243 = 14'h1d == field_data_lo_28 ? _field_data_T_33 : _GEN_2242; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2244 = 14'h1e == field_data_lo_28 ? _field_data_T_34 : _GEN_2243; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2245 = 14'h1f == field_data_lo_28 ? _field_data_T_35 : _GEN_2244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2246 = 14'h20 == field_data_lo_28 ? _field_data_T_36 : _GEN_2245; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2247 = 14'h21 == field_data_lo_28 ? _field_data_T_37 : _GEN_2246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2248 = 14'h22 == field_data_lo_28 ? _field_data_T_38 : _GEN_2247; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2249 = 14'h23 == field_data_lo_28 ? _field_data_T_39 : _GEN_2248; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2250 = 14'h24 == field_data_lo_28 ? _field_data_T_40 : _GEN_2249; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2251 = 14'h25 == field_data_lo_28 ? _field_data_T_41 : _GEN_2250; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2252 = 14'h26 == field_data_lo_28 ? _field_data_T_42 : _GEN_2251; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2253 = 14'h27 == field_data_lo_28 ? _field_data_T_43 : _GEN_2252; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2254 = 14'h28 == field_data_lo_28 ? _field_data_T_44 : _GEN_2253; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2255 = 14'h29 == field_data_lo_28 ? _field_data_T_45 : _GEN_2254; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2256 = 14'h2a == field_data_lo_28 ? _field_data_T_46 : _GEN_2255; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2257 = 14'h2b == field_data_lo_28 ? _field_data_T_47 : _GEN_2256; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2258 = 14'h2c == field_data_lo_28 ? _field_data_T_48 : _GEN_2257; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2259 = 14'h2d == field_data_lo_28 ? _field_data_T_49 : _GEN_2258; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2260 = 14'h2e == field_data_lo_28 ? _field_data_T_50 : _GEN_2259; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2261 = 14'h2f == field_data_lo_28 ? _field_data_T_51 : _GEN_2260; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2262 = 14'h30 == field_data_lo_28 ? _field_data_T_52 : _GEN_2261; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2263 = 14'h31 == field_data_lo_28 ? _field_data_T_53 : _GEN_2262; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_49 = vliw_49[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_29 = vliw_49[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_49 = field_data_lo_29[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_49 = field_data_lo_29[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_78 = {{1'd0}, args_offset_49}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_78 = _total_offset_T_78[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2267 = 3'h1 == total_offset_78 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2268 = 3'h2 == total_offset_78 ? args_2 : _GEN_2267; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2269 = 3'h3 == total_offset_78 ? args_3 : _GEN_2268; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2270 = 3'h4 == total_offset_78 ? args_4 : _GEN_2269; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2271 = 3'h5 == total_offset_78 ? args_5 : _GEN_2270; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2272 = 3'h6 == total_offset_78 ? args_6 : _GEN_2271; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2273 = total_offset_78 < 3'h7 ? _GEN_2272 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_49_1 = 3'h0 < args_length_49 ? _GEN_2273 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_79 = args_offset_49 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2276 = 3'h1 == total_offset_79 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2277 = 3'h2 == total_offset_79 ? args_2 : _GEN_2276; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2278 = 3'h3 == total_offset_79 ? args_3 : _GEN_2277; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2279 = 3'h4 == total_offset_79 ? args_4 : _GEN_2278; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2280 = 3'h5 == total_offset_79 ? args_5 : _GEN_2279; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2281 = 3'h6 == total_offset_79 ? args_6 : _GEN_2280; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2282 = total_offset_79 < 3'h7 ? _GEN_2281 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_49_0 = 3'h1 < args_length_49 ? _GEN_2282 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [15:0] _field_data_T_1006 = {field_bytes_49_0,field_bytes_49_1}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_2284 = opcode_49 == 4'ha ? _field_data_T_1006 : 16'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2285 = opcode_49 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1676 = opcode_49 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [1:0] field_data_hi_29 = field_data_lo_29[13] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _field_data_T_1009 = {field_data_hi_29,field_data_lo_29}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_99 = _T_1676 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [15:0] _GEN_2286 = opcode_49 == 4'h8 | opcode_49 == 4'hb ? _field_data_T_1009 : _GEN_2284; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2287 = opcode_49 == 4'h8 | opcode_49 == 4'hb ? _field_tag_T_99 : _GEN_2285; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [15:0] _GEN_2288 = 14'h14 == field_data_lo_29 ? _field_data_T_24 : _GEN_2286; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2289 = 14'h15 == field_data_lo_29 ? _field_data_T_25 : _GEN_2288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2290 = 14'h16 == field_data_lo_29 ? _field_data_T_26 : _GEN_2289; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2291 = 14'h17 == field_data_lo_29 ? _field_data_T_27 : _GEN_2290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2292 = 14'h18 == field_data_lo_29 ? _field_data_T_28 : _GEN_2291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2293 = 14'h19 == field_data_lo_29 ? _field_data_T_29 : _GEN_2292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2294 = 14'h1a == field_data_lo_29 ? _field_data_T_30 : _GEN_2293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2295 = 14'h1b == field_data_lo_29 ? _field_data_T_31 : _GEN_2294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2296 = 14'h1c == field_data_lo_29 ? _field_data_T_32 : _GEN_2295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2297 = 14'h1d == field_data_lo_29 ? _field_data_T_33 : _GEN_2296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2298 = 14'h1e == field_data_lo_29 ? _field_data_T_34 : _GEN_2297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2299 = 14'h1f == field_data_lo_29 ? _field_data_T_35 : _GEN_2298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2300 = 14'h20 == field_data_lo_29 ? _field_data_T_36 : _GEN_2299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2301 = 14'h21 == field_data_lo_29 ? _field_data_T_37 : _GEN_2300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2302 = 14'h22 == field_data_lo_29 ? _field_data_T_38 : _GEN_2301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2303 = 14'h23 == field_data_lo_29 ? _field_data_T_39 : _GEN_2302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2304 = 14'h24 == field_data_lo_29 ? _field_data_T_40 : _GEN_2303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2305 = 14'h25 == field_data_lo_29 ? _field_data_T_41 : _GEN_2304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2306 = 14'h26 == field_data_lo_29 ? _field_data_T_42 : _GEN_2305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2307 = 14'h27 == field_data_lo_29 ? _field_data_T_43 : _GEN_2306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2308 = 14'h28 == field_data_lo_29 ? _field_data_T_44 : _GEN_2307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2309 = 14'h29 == field_data_lo_29 ? _field_data_T_45 : _GEN_2308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2310 = 14'h2a == field_data_lo_29 ? _field_data_T_46 : _GEN_2309; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2311 = 14'h2b == field_data_lo_29 ? _field_data_T_47 : _GEN_2310; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2312 = 14'h2c == field_data_lo_29 ? _field_data_T_48 : _GEN_2311; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2313 = 14'h2d == field_data_lo_29 ? _field_data_T_49 : _GEN_2312; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2314 = 14'h2e == field_data_lo_29 ? _field_data_T_50 : _GEN_2313; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2315 = 14'h2f == field_data_lo_29 ? _field_data_T_51 : _GEN_2314; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2316 = 14'h30 == field_data_lo_29 ? _field_data_T_52 : _GEN_2315; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [15:0] _GEN_2317 = 14'h31 == field_data_lo_29 ? _field_data_T_53 : _GEN_2316; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_50 = vliw_50[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_30 = vliw_50[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_50 = field_data_lo_30[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_50 = field_data_lo_30[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_80 = {{1'd0}, args_offset_50}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_80 = _total_offset_T_80[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2321 = 3'h1 == total_offset_80 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2322 = 3'h2 == total_offset_80 ? args_2 : _GEN_2321; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2323 = 3'h3 == total_offset_80 ? args_3 : _GEN_2322; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2324 = 3'h4 == total_offset_80 ? args_4 : _GEN_2323; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2325 = 3'h5 == total_offset_80 ? args_5 : _GEN_2324; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2326 = 3'h6 == total_offset_80 ? args_6 : _GEN_2325; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2327 = total_offset_80 < 3'h7 ? _GEN_2326 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_50_3 = 3'h0 < args_length_50 ? _GEN_2327 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_81 = args_offset_50 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2330 = 3'h1 == total_offset_81 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2331 = 3'h2 == total_offset_81 ? args_2 : _GEN_2330; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2332 = 3'h3 == total_offset_81 ? args_3 : _GEN_2331; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2333 = 3'h4 == total_offset_81 ? args_4 : _GEN_2332; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2334 = 3'h5 == total_offset_81 ? args_5 : _GEN_2333; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2335 = 3'h6 == total_offset_81 ? args_6 : _GEN_2334; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2336 = total_offset_81 < 3'h7 ? _GEN_2335 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_50_2 = 3'h1 < args_length_50 ? _GEN_2336 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_82 = args_offset_50 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2339 = 3'h1 == total_offset_82 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2340 = 3'h2 == total_offset_82 ? args_2 : _GEN_2339; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2341 = 3'h3 == total_offset_82 ? args_3 : _GEN_2340; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2342 = 3'h4 == total_offset_82 ? args_4 : _GEN_2341; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2343 = 3'h5 == total_offset_82 ? args_5 : _GEN_2342; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2344 = 3'h6 == total_offset_82 ? args_6 : _GEN_2343; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2345 = total_offset_82 < 3'h7 ? _GEN_2344 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_50_1 = 3'h2 < args_length_50 ? _GEN_2345 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_83 = args_offset_50 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2348 = 3'h1 == total_offset_83 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2349 = 3'h2 == total_offset_83 ? args_2 : _GEN_2348; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2350 = 3'h3 == total_offset_83 ? args_3 : _GEN_2349; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2351 = 3'h4 == total_offset_83 ? args_4 : _GEN_2350; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2352 = 3'h5 == total_offset_83 ? args_5 : _GEN_2351; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2353 = 3'h6 == total_offset_83 ? args_6 : _GEN_2352; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2354 = total_offset_83 < 3'h7 ? _GEN_2353 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_50_0 = 3'h3 < args_length_50 ? _GEN_2354 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1040 = {field_bytes_50_0,field_bytes_50_1,field_bytes_50_2,field_bytes_50_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2356 = opcode_50 == 4'ha ? _field_data_T_1040 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2357 = opcode_50 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1719 = opcode_50 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_32 = field_data_lo_30[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1043 = {field_data_hi_32,field_data_lo_30}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_101 = _T_1719 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2358 = opcode_50 == 4'h8 | opcode_50 == 4'hb ? _field_data_T_1043 : _GEN_2356; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2359 = opcode_50 == 4'h8 | opcode_50 == 4'hb ? _field_tag_T_101 : _GEN_2357; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _field_data_T_1044 = {phv_data_80,phv_data_81,phv_data_82,phv_data_83}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2360 = 14'h32 == field_data_lo_30 ? _field_data_T_1044 : _GEN_2358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1045 = {phv_data_84,phv_data_85,phv_data_86,phv_data_87}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2361 = 14'h33 == field_data_lo_30 ? _field_data_T_1045 : _GEN_2360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1046 = {phv_data_88,phv_data_89,phv_data_90,phv_data_91}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2362 = 14'h34 == field_data_lo_30 ? _field_data_T_1046 : _GEN_2361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1047 = {phv_data_92,phv_data_93,phv_data_94,phv_data_95}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2363 = 14'h35 == field_data_lo_30 ? _field_data_T_1047 : _GEN_2362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1048 = {phv_data_96,phv_data_97,phv_data_98,phv_data_99}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2364 = 14'h36 == field_data_lo_30 ? _field_data_T_1048 : _GEN_2363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1049 = {phv_data_100,phv_data_101,phv_data_102,phv_data_103}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2365 = 14'h37 == field_data_lo_30 ? _field_data_T_1049 : _GEN_2364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1050 = {phv_data_104,phv_data_105,phv_data_106,phv_data_107}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2366 = 14'h38 == field_data_lo_30 ? _field_data_T_1050 : _GEN_2365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1051 = {phv_data_108,phv_data_109,phv_data_110,phv_data_111}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2367 = 14'h39 == field_data_lo_30 ? _field_data_T_1051 : _GEN_2366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1052 = {phv_data_112,phv_data_113,phv_data_114,phv_data_115}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2368 = 14'h3a == field_data_lo_30 ? _field_data_T_1052 : _GEN_2367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1053 = {phv_data_116,phv_data_117,phv_data_118,phv_data_119}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2369 = 14'h3b == field_data_lo_30 ? _field_data_T_1053 : _GEN_2368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1054 = {phv_data_120,phv_data_121,phv_data_122,phv_data_123}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2370 = 14'h3c == field_data_lo_30 ? _field_data_T_1054 : _GEN_2369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1055 = {phv_data_124,phv_data_125,phv_data_126,phv_data_127}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2371 = 14'h3d == field_data_lo_30 ? _field_data_T_1055 : _GEN_2370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1056 = {phv_data_128,phv_data_129,phv_data_130,phv_data_131}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2372 = 14'h3e == field_data_lo_30 ? _field_data_T_1056 : _GEN_2371; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1057 = {phv_data_132,phv_data_133,phv_data_134,phv_data_135}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2373 = 14'h3f == field_data_lo_30 ? _field_data_T_1057 : _GEN_2372; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1058 = {phv_data_136,phv_data_137,phv_data_138,phv_data_139}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2374 = 14'h40 == field_data_lo_30 ? _field_data_T_1058 : _GEN_2373; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1059 = {phv_data_140,phv_data_141,phv_data_142,phv_data_143}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2375 = 14'h41 == field_data_lo_30 ? _field_data_T_1059 : _GEN_2374; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1060 = {phv_data_144,phv_data_145,phv_data_146,phv_data_147}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2376 = 14'h42 == field_data_lo_30 ? _field_data_T_1060 : _GEN_2375; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1061 = {phv_data_148,phv_data_149,phv_data_150,phv_data_151}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2377 = 14'h43 == field_data_lo_30 ? _field_data_T_1061 : _GEN_2376; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1062 = {phv_data_152,phv_data_153,phv_data_154,phv_data_155}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2378 = 14'h44 == field_data_lo_30 ? _field_data_T_1062 : _GEN_2377; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _field_data_T_1063 = {phv_data_156,phv_data_157,phv_data_158,phv_data_159}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2379 = 14'h45 == field_data_lo_30 ? _field_data_T_1063 : _GEN_2378; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_51 = vliw_51[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_51 = vliw_51[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_51 = field_data_lo_51[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_51 = field_data_lo_51[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_84 = {{1'd0}, args_offset_51}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_84 = _total_offset_T_84[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2383 = 3'h1 == total_offset_84 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2384 = 3'h2 == total_offset_84 ? args_2 : _GEN_2383; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2385 = 3'h3 == total_offset_84 ? args_3 : _GEN_2384; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2386 = 3'h4 == total_offset_84 ? args_4 : _GEN_2385; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2387 = 3'h5 == total_offset_84 ? args_5 : _GEN_2386; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2388 = 3'h6 == total_offset_84 ? args_6 : _GEN_2387; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2389 = total_offset_84 < 3'h7 ? _GEN_2388 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_51_3 = 3'h0 < args_length_51 ? _GEN_2389 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_85 = args_offset_51 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2392 = 3'h1 == total_offset_85 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2393 = 3'h2 == total_offset_85 ? args_2 : _GEN_2392; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2394 = 3'h3 == total_offset_85 ? args_3 : _GEN_2393; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2395 = 3'h4 == total_offset_85 ? args_4 : _GEN_2394; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2396 = 3'h5 == total_offset_85 ? args_5 : _GEN_2395; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2397 = 3'h6 == total_offset_85 ? args_6 : _GEN_2396; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2398 = total_offset_85 < 3'h7 ? _GEN_2397 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_51_2 = 3'h1 < args_length_51 ? _GEN_2398 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_86 = args_offset_51 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2401 = 3'h1 == total_offset_86 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2402 = 3'h2 == total_offset_86 ? args_2 : _GEN_2401; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2403 = 3'h3 == total_offset_86 ? args_3 : _GEN_2402; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2404 = 3'h4 == total_offset_86 ? args_4 : _GEN_2403; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2405 = 3'h5 == total_offset_86 ? args_5 : _GEN_2404; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2406 = 3'h6 == total_offset_86 ? args_6 : _GEN_2405; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2407 = total_offset_86 < 3'h7 ? _GEN_2406 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_51_1 = 3'h2 < args_length_51 ? _GEN_2407 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_87 = args_offset_51 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2410 = 3'h1 == total_offset_87 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2411 = 3'h2 == total_offset_87 ? args_2 : _GEN_2410; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2412 = 3'h3 == total_offset_87 ? args_3 : _GEN_2411; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2413 = 3'h4 == total_offset_87 ? args_4 : _GEN_2412; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2414 = 3'h5 == total_offset_87 ? args_5 : _GEN_2413; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2415 = 3'h6 == total_offset_87 ? args_6 : _GEN_2414; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2416 = total_offset_87 < 3'h7 ? _GEN_2415 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_51_0 = 3'h3 < args_length_51 ? _GEN_2416 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1064 = {field_bytes_51_0,field_bytes_51_1,field_bytes_51_2,field_bytes_51_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2418 = opcode_51 == 4'ha ? _field_data_T_1064 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2419 = opcode_51 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1752 = opcode_51 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_55 = field_data_lo_51[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1067 = {field_data_hi_55,field_data_lo_51}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_103 = _T_1752 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2420 = opcode_51 == 4'h8 | opcode_51 == 4'hb ? _field_data_T_1067 : _GEN_2418; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2421 = opcode_51 == 4'h8 | opcode_51 == 4'hb ? _field_tag_T_103 : _GEN_2419; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2422 = 14'h32 == field_data_lo_51 ? _field_data_T_1044 : _GEN_2420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2423 = 14'h33 == field_data_lo_51 ? _field_data_T_1045 : _GEN_2422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2424 = 14'h34 == field_data_lo_51 ? _field_data_T_1046 : _GEN_2423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2425 = 14'h35 == field_data_lo_51 ? _field_data_T_1047 : _GEN_2424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2426 = 14'h36 == field_data_lo_51 ? _field_data_T_1048 : _GEN_2425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2427 = 14'h37 == field_data_lo_51 ? _field_data_T_1049 : _GEN_2426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2428 = 14'h38 == field_data_lo_51 ? _field_data_T_1050 : _GEN_2427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2429 = 14'h39 == field_data_lo_51 ? _field_data_T_1051 : _GEN_2428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2430 = 14'h3a == field_data_lo_51 ? _field_data_T_1052 : _GEN_2429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2431 = 14'h3b == field_data_lo_51 ? _field_data_T_1053 : _GEN_2430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2432 = 14'h3c == field_data_lo_51 ? _field_data_T_1054 : _GEN_2431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2433 = 14'h3d == field_data_lo_51 ? _field_data_T_1055 : _GEN_2432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2434 = 14'h3e == field_data_lo_51 ? _field_data_T_1056 : _GEN_2433; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2435 = 14'h3f == field_data_lo_51 ? _field_data_T_1057 : _GEN_2434; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2436 = 14'h40 == field_data_lo_51 ? _field_data_T_1058 : _GEN_2435; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2437 = 14'h41 == field_data_lo_51 ? _field_data_T_1059 : _GEN_2436; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2438 = 14'h42 == field_data_lo_51 ? _field_data_T_1060 : _GEN_2437; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2439 = 14'h43 == field_data_lo_51 ? _field_data_T_1061 : _GEN_2438; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2440 = 14'h44 == field_data_lo_51 ? _field_data_T_1062 : _GEN_2439; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2441 = 14'h45 == field_data_lo_51 ? _field_data_T_1063 : _GEN_2440; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_52 = vliw_52[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_72 = vliw_52[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_52 = field_data_lo_72[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_52 = field_data_lo_72[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_88 = {{1'd0}, args_offset_52}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_88 = _total_offset_T_88[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2445 = 3'h1 == total_offset_88 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2446 = 3'h2 == total_offset_88 ? args_2 : _GEN_2445; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2447 = 3'h3 == total_offset_88 ? args_3 : _GEN_2446; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2448 = 3'h4 == total_offset_88 ? args_4 : _GEN_2447; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2449 = 3'h5 == total_offset_88 ? args_5 : _GEN_2448; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2450 = 3'h6 == total_offset_88 ? args_6 : _GEN_2449; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2451 = total_offset_88 < 3'h7 ? _GEN_2450 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_52_3 = 3'h0 < args_length_52 ? _GEN_2451 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_89 = args_offset_52 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2454 = 3'h1 == total_offset_89 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2455 = 3'h2 == total_offset_89 ? args_2 : _GEN_2454; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2456 = 3'h3 == total_offset_89 ? args_3 : _GEN_2455; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2457 = 3'h4 == total_offset_89 ? args_4 : _GEN_2456; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2458 = 3'h5 == total_offset_89 ? args_5 : _GEN_2457; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2459 = 3'h6 == total_offset_89 ? args_6 : _GEN_2458; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2460 = total_offset_89 < 3'h7 ? _GEN_2459 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_52_2 = 3'h1 < args_length_52 ? _GEN_2460 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_90 = args_offset_52 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2463 = 3'h1 == total_offset_90 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2464 = 3'h2 == total_offset_90 ? args_2 : _GEN_2463; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2465 = 3'h3 == total_offset_90 ? args_3 : _GEN_2464; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2466 = 3'h4 == total_offset_90 ? args_4 : _GEN_2465; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2467 = 3'h5 == total_offset_90 ? args_5 : _GEN_2466; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2468 = 3'h6 == total_offset_90 ? args_6 : _GEN_2467; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2469 = total_offset_90 < 3'h7 ? _GEN_2468 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_52_1 = 3'h2 < args_length_52 ? _GEN_2469 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_91 = args_offset_52 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2472 = 3'h1 == total_offset_91 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2473 = 3'h2 == total_offset_91 ? args_2 : _GEN_2472; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2474 = 3'h3 == total_offset_91 ? args_3 : _GEN_2473; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2475 = 3'h4 == total_offset_91 ? args_4 : _GEN_2474; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2476 = 3'h5 == total_offset_91 ? args_5 : _GEN_2475; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2477 = 3'h6 == total_offset_91 ? args_6 : _GEN_2476; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2478 = total_offset_91 < 3'h7 ? _GEN_2477 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_52_0 = 3'h3 < args_length_52 ? _GEN_2478 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1088 = {field_bytes_52_0,field_bytes_52_1,field_bytes_52_2,field_bytes_52_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2480 = opcode_52 == 4'ha ? _field_data_T_1088 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2481 = opcode_52 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1785 = opcode_52 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_78 = field_data_lo_72[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1091 = {field_data_hi_78,field_data_lo_72}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_105 = _T_1785 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2482 = opcode_52 == 4'h8 | opcode_52 == 4'hb ? _field_data_T_1091 : _GEN_2480; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2483 = opcode_52 == 4'h8 | opcode_52 == 4'hb ? _field_tag_T_105 : _GEN_2481; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2484 = 14'h32 == field_data_lo_72 ? _field_data_T_1044 : _GEN_2482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2485 = 14'h33 == field_data_lo_72 ? _field_data_T_1045 : _GEN_2484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2486 = 14'h34 == field_data_lo_72 ? _field_data_T_1046 : _GEN_2485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2487 = 14'h35 == field_data_lo_72 ? _field_data_T_1047 : _GEN_2486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2488 = 14'h36 == field_data_lo_72 ? _field_data_T_1048 : _GEN_2487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2489 = 14'h37 == field_data_lo_72 ? _field_data_T_1049 : _GEN_2488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2490 = 14'h38 == field_data_lo_72 ? _field_data_T_1050 : _GEN_2489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2491 = 14'h39 == field_data_lo_72 ? _field_data_T_1051 : _GEN_2490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2492 = 14'h3a == field_data_lo_72 ? _field_data_T_1052 : _GEN_2491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2493 = 14'h3b == field_data_lo_72 ? _field_data_T_1053 : _GEN_2492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2494 = 14'h3c == field_data_lo_72 ? _field_data_T_1054 : _GEN_2493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2495 = 14'h3d == field_data_lo_72 ? _field_data_T_1055 : _GEN_2494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2496 = 14'h3e == field_data_lo_72 ? _field_data_T_1056 : _GEN_2495; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2497 = 14'h3f == field_data_lo_72 ? _field_data_T_1057 : _GEN_2496; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2498 = 14'h40 == field_data_lo_72 ? _field_data_T_1058 : _GEN_2497; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2499 = 14'h41 == field_data_lo_72 ? _field_data_T_1059 : _GEN_2498; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2500 = 14'h42 == field_data_lo_72 ? _field_data_T_1060 : _GEN_2499; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2501 = 14'h43 == field_data_lo_72 ? _field_data_T_1061 : _GEN_2500; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2502 = 14'h44 == field_data_lo_72 ? _field_data_T_1062 : _GEN_2501; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2503 = 14'h45 == field_data_lo_72 ? _field_data_T_1063 : _GEN_2502; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_53 = vliw_53[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_93 = vliw_53[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_53 = field_data_lo_93[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_53 = field_data_lo_93[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_92 = {{1'd0}, args_offset_53}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_92 = _total_offset_T_92[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2507 = 3'h1 == total_offset_92 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2508 = 3'h2 == total_offset_92 ? args_2 : _GEN_2507; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2509 = 3'h3 == total_offset_92 ? args_3 : _GEN_2508; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2510 = 3'h4 == total_offset_92 ? args_4 : _GEN_2509; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2511 = 3'h5 == total_offset_92 ? args_5 : _GEN_2510; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2512 = 3'h6 == total_offset_92 ? args_6 : _GEN_2511; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2513 = total_offset_92 < 3'h7 ? _GEN_2512 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_53_3 = 3'h0 < args_length_53 ? _GEN_2513 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_93 = args_offset_53 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2516 = 3'h1 == total_offset_93 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2517 = 3'h2 == total_offset_93 ? args_2 : _GEN_2516; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2518 = 3'h3 == total_offset_93 ? args_3 : _GEN_2517; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2519 = 3'h4 == total_offset_93 ? args_4 : _GEN_2518; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2520 = 3'h5 == total_offset_93 ? args_5 : _GEN_2519; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2521 = 3'h6 == total_offset_93 ? args_6 : _GEN_2520; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2522 = total_offset_93 < 3'h7 ? _GEN_2521 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_53_2 = 3'h1 < args_length_53 ? _GEN_2522 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_94 = args_offset_53 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2525 = 3'h1 == total_offset_94 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2526 = 3'h2 == total_offset_94 ? args_2 : _GEN_2525; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2527 = 3'h3 == total_offset_94 ? args_3 : _GEN_2526; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2528 = 3'h4 == total_offset_94 ? args_4 : _GEN_2527; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2529 = 3'h5 == total_offset_94 ? args_5 : _GEN_2528; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2530 = 3'h6 == total_offset_94 ? args_6 : _GEN_2529; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2531 = total_offset_94 < 3'h7 ? _GEN_2530 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_53_1 = 3'h2 < args_length_53 ? _GEN_2531 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_95 = args_offset_53 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2534 = 3'h1 == total_offset_95 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2535 = 3'h2 == total_offset_95 ? args_2 : _GEN_2534; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2536 = 3'h3 == total_offset_95 ? args_3 : _GEN_2535; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2537 = 3'h4 == total_offset_95 ? args_4 : _GEN_2536; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2538 = 3'h5 == total_offset_95 ? args_5 : _GEN_2537; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2539 = 3'h6 == total_offset_95 ? args_6 : _GEN_2538; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2540 = total_offset_95 < 3'h7 ? _GEN_2539 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_53_0 = 3'h3 < args_length_53 ? _GEN_2540 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1112 = {field_bytes_53_0,field_bytes_53_1,field_bytes_53_2,field_bytes_53_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2542 = opcode_53 == 4'ha ? _field_data_T_1112 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2543 = opcode_53 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1818 = opcode_53 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_101 = field_data_lo_93[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1115 = {field_data_hi_101,field_data_lo_93}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_107 = _T_1818 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2544 = opcode_53 == 4'h8 | opcode_53 == 4'hb ? _field_data_T_1115 : _GEN_2542; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2545 = opcode_53 == 4'h8 | opcode_53 == 4'hb ? _field_tag_T_107 : _GEN_2543; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2546 = 14'h32 == field_data_lo_93 ? _field_data_T_1044 : _GEN_2544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2547 = 14'h33 == field_data_lo_93 ? _field_data_T_1045 : _GEN_2546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2548 = 14'h34 == field_data_lo_93 ? _field_data_T_1046 : _GEN_2547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2549 = 14'h35 == field_data_lo_93 ? _field_data_T_1047 : _GEN_2548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2550 = 14'h36 == field_data_lo_93 ? _field_data_T_1048 : _GEN_2549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2551 = 14'h37 == field_data_lo_93 ? _field_data_T_1049 : _GEN_2550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2552 = 14'h38 == field_data_lo_93 ? _field_data_T_1050 : _GEN_2551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2553 = 14'h39 == field_data_lo_93 ? _field_data_T_1051 : _GEN_2552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2554 = 14'h3a == field_data_lo_93 ? _field_data_T_1052 : _GEN_2553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2555 = 14'h3b == field_data_lo_93 ? _field_data_T_1053 : _GEN_2554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2556 = 14'h3c == field_data_lo_93 ? _field_data_T_1054 : _GEN_2555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2557 = 14'h3d == field_data_lo_93 ? _field_data_T_1055 : _GEN_2556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2558 = 14'h3e == field_data_lo_93 ? _field_data_T_1056 : _GEN_2557; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2559 = 14'h3f == field_data_lo_93 ? _field_data_T_1057 : _GEN_2558; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2560 = 14'h40 == field_data_lo_93 ? _field_data_T_1058 : _GEN_2559; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2561 = 14'h41 == field_data_lo_93 ? _field_data_T_1059 : _GEN_2560; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2562 = 14'h42 == field_data_lo_93 ? _field_data_T_1060 : _GEN_2561; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2563 = 14'h43 == field_data_lo_93 ? _field_data_T_1061 : _GEN_2562; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2564 = 14'h44 == field_data_lo_93 ? _field_data_T_1062 : _GEN_2563; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2565 = 14'h45 == field_data_lo_93 ? _field_data_T_1063 : _GEN_2564; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_54 = vliw_54[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_114 = vliw_54[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_54 = field_data_lo_114[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_54 = field_data_lo_114[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_96 = {{1'd0}, args_offset_54}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_96 = _total_offset_T_96[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2569 = 3'h1 == total_offset_96 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2570 = 3'h2 == total_offset_96 ? args_2 : _GEN_2569; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2571 = 3'h3 == total_offset_96 ? args_3 : _GEN_2570; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2572 = 3'h4 == total_offset_96 ? args_4 : _GEN_2571; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2573 = 3'h5 == total_offset_96 ? args_5 : _GEN_2572; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2574 = 3'h6 == total_offset_96 ? args_6 : _GEN_2573; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2575 = total_offset_96 < 3'h7 ? _GEN_2574 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_54_3 = 3'h0 < args_length_54 ? _GEN_2575 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_97 = args_offset_54 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2578 = 3'h1 == total_offset_97 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2579 = 3'h2 == total_offset_97 ? args_2 : _GEN_2578; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2580 = 3'h3 == total_offset_97 ? args_3 : _GEN_2579; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2581 = 3'h4 == total_offset_97 ? args_4 : _GEN_2580; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2582 = 3'h5 == total_offset_97 ? args_5 : _GEN_2581; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2583 = 3'h6 == total_offset_97 ? args_6 : _GEN_2582; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2584 = total_offset_97 < 3'h7 ? _GEN_2583 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_54_2 = 3'h1 < args_length_54 ? _GEN_2584 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_98 = args_offset_54 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2587 = 3'h1 == total_offset_98 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2588 = 3'h2 == total_offset_98 ? args_2 : _GEN_2587; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2589 = 3'h3 == total_offset_98 ? args_3 : _GEN_2588; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2590 = 3'h4 == total_offset_98 ? args_4 : _GEN_2589; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2591 = 3'h5 == total_offset_98 ? args_5 : _GEN_2590; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2592 = 3'h6 == total_offset_98 ? args_6 : _GEN_2591; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2593 = total_offset_98 < 3'h7 ? _GEN_2592 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_54_1 = 3'h2 < args_length_54 ? _GEN_2593 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_99 = args_offset_54 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2596 = 3'h1 == total_offset_99 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2597 = 3'h2 == total_offset_99 ? args_2 : _GEN_2596; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2598 = 3'h3 == total_offset_99 ? args_3 : _GEN_2597; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2599 = 3'h4 == total_offset_99 ? args_4 : _GEN_2598; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2600 = 3'h5 == total_offset_99 ? args_5 : _GEN_2599; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2601 = 3'h6 == total_offset_99 ? args_6 : _GEN_2600; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2602 = total_offset_99 < 3'h7 ? _GEN_2601 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_54_0 = 3'h3 < args_length_54 ? _GEN_2602 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1136 = {field_bytes_54_0,field_bytes_54_1,field_bytes_54_2,field_bytes_54_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2604 = opcode_54 == 4'ha ? _field_data_T_1136 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2605 = opcode_54 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1851 = opcode_54 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_124 = field_data_lo_114[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1139 = {field_data_hi_124,field_data_lo_114}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_109 = _T_1851 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2606 = opcode_54 == 4'h8 | opcode_54 == 4'hb ? _field_data_T_1139 : _GEN_2604; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2607 = opcode_54 == 4'h8 | opcode_54 == 4'hb ? _field_tag_T_109 : _GEN_2605; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2608 = 14'h32 == field_data_lo_114 ? _field_data_T_1044 : _GEN_2606; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2609 = 14'h33 == field_data_lo_114 ? _field_data_T_1045 : _GEN_2608; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2610 = 14'h34 == field_data_lo_114 ? _field_data_T_1046 : _GEN_2609; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2611 = 14'h35 == field_data_lo_114 ? _field_data_T_1047 : _GEN_2610; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2612 = 14'h36 == field_data_lo_114 ? _field_data_T_1048 : _GEN_2611; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2613 = 14'h37 == field_data_lo_114 ? _field_data_T_1049 : _GEN_2612; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2614 = 14'h38 == field_data_lo_114 ? _field_data_T_1050 : _GEN_2613; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2615 = 14'h39 == field_data_lo_114 ? _field_data_T_1051 : _GEN_2614; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2616 = 14'h3a == field_data_lo_114 ? _field_data_T_1052 : _GEN_2615; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2617 = 14'h3b == field_data_lo_114 ? _field_data_T_1053 : _GEN_2616; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2618 = 14'h3c == field_data_lo_114 ? _field_data_T_1054 : _GEN_2617; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2619 = 14'h3d == field_data_lo_114 ? _field_data_T_1055 : _GEN_2618; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2620 = 14'h3e == field_data_lo_114 ? _field_data_T_1056 : _GEN_2619; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2621 = 14'h3f == field_data_lo_114 ? _field_data_T_1057 : _GEN_2620; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2622 = 14'h40 == field_data_lo_114 ? _field_data_T_1058 : _GEN_2621; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2623 = 14'h41 == field_data_lo_114 ? _field_data_T_1059 : _GEN_2622; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2624 = 14'h42 == field_data_lo_114 ? _field_data_T_1060 : _GEN_2623; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2625 = 14'h43 == field_data_lo_114 ? _field_data_T_1061 : _GEN_2624; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2626 = 14'h44 == field_data_lo_114 ? _field_data_T_1062 : _GEN_2625; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2627 = 14'h45 == field_data_lo_114 ? _field_data_T_1063 : _GEN_2626; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_55 = vliw_55[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_135 = vliw_55[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_55 = field_data_lo_135[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_55 = field_data_lo_135[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_100 = {{1'd0}, args_offset_55}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_100 = _total_offset_T_100[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2631 = 3'h1 == total_offset_100 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2632 = 3'h2 == total_offset_100 ? args_2 : _GEN_2631; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2633 = 3'h3 == total_offset_100 ? args_3 : _GEN_2632; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2634 = 3'h4 == total_offset_100 ? args_4 : _GEN_2633; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2635 = 3'h5 == total_offset_100 ? args_5 : _GEN_2634; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2636 = 3'h6 == total_offset_100 ? args_6 : _GEN_2635; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2637 = total_offset_100 < 3'h7 ? _GEN_2636 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_55_3 = 3'h0 < args_length_55 ? _GEN_2637 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_101 = args_offset_55 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2640 = 3'h1 == total_offset_101 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2641 = 3'h2 == total_offset_101 ? args_2 : _GEN_2640; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2642 = 3'h3 == total_offset_101 ? args_3 : _GEN_2641; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2643 = 3'h4 == total_offset_101 ? args_4 : _GEN_2642; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2644 = 3'h5 == total_offset_101 ? args_5 : _GEN_2643; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2645 = 3'h6 == total_offset_101 ? args_6 : _GEN_2644; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2646 = total_offset_101 < 3'h7 ? _GEN_2645 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_55_2 = 3'h1 < args_length_55 ? _GEN_2646 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_102 = args_offset_55 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2649 = 3'h1 == total_offset_102 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2650 = 3'h2 == total_offset_102 ? args_2 : _GEN_2649; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2651 = 3'h3 == total_offset_102 ? args_3 : _GEN_2650; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2652 = 3'h4 == total_offset_102 ? args_4 : _GEN_2651; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2653 = 3'h5 == total_offset_102 ? args_5 : _GEN_2652; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2654 = 3'h6 == total_offset_102 ? args_6 : _GEN_2653; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2655 = total_offset_102 < 3'h7 ? _GEN_2654 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_55_1 = 3'h2 < args_length_55 ? _GEN_2655 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_103 = args_offset_55 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2658 = 3'h1 == total_offset_103 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2659 = 3'h2 == total_offset_103 ? args_2 : _GEN_2658; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2660 = 3'h3 == total_offset_103 ? args_3 : _GEN_2659; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2661 = 3'h4 == total_offset_103 ? args_4 : _GEN_2660; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2662 = 3'h5 == total_offset_103 ? args_5 : _GEN_2661; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2663 = 3'h6 == total_offset_103 ? args_6 : _GEN_2662; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2664 = total_offset_103 < 3'h7 ? _GEN_2663 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_55_0 = 3'h3 < args_length_55 ? _GEN_2664 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1160 = {field_bytes_55_0,field_bytes_55_1,field_bytes_55_2,field_bytes_55_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2666 = opcode_55 == 4'ha ? _field_data_T_1160 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2667 = opcode_55 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1884 = opcode_55 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_147 = field_data_lo_135[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1163 = {field_data_hi_147,field_data_lo_135}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_111 = _T_1884 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2668 = opcode_55 == 4'h8 | opcode_55 == 4'hb ? _field_data_T_1163 : _GEN_2666; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2669 = opcode_55 == 4'h8 | opcode_55 == 4'hb ? _field_tag_T_111 : _GEN_2667; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2670 = 14'h32 == field_data_lo_135 ? _field_data_T_1044 : _GEN_2668; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2671 = 14'h33 == field_data_lo_135 ? _field_data_T_1045 : _GEN_2670; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2672 = 14'h34 == field_data_lo_135 ? _field_data_T_1046 : _GEN_2671; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2673 = 14'h35 == field_data_lo_135 ? _field_data_T_1047 : _GEN_2672; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2674 = 14'h36 == field_data_lo_135 ? _field_data_T_1048 : _GEN_2673; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2675 = 14'h37 == field_data_lo_135 ? _field_data_T_1049 : _GEN_2674; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2676 = 14'h38 == field_data_lo_135 ? _field_data_T_1050 : _GEN_2675; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2677 = 14'h39 == field_data_lo_135 ? _field_data_T_1051 : _GEN_2676; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2678 = 14'h3a == field_data_lo_135 ? _field_data_T_1052 : _GEN_2677; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2679 = 14'h3b == field_data_lo_135 ? _field_data_T_1053 : _GEN_2678; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2680 = 14'h3c == field_data_lo_135 ? _field_data_T_1054 : _GEN_2679; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2681 = 14'h3d == field_data_lo_135 ? _field_data_T_1055 : _GEN_2680; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2682 = 14'h3e == field_data_lo_135 ? _field_data_T_1056 : _GEN_2681; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2683 = 14'h3f == field_data_lo_135 ? _field_data_T_1057 : _GEN_2682; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2684 = 14'h40 == field_data_lo_135 ? _field_data_T_1058 : _GEN_2683; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2685 = 14'h41 == field_data_lo_135 ? _field_data_T_1059 : _GEN_2684; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2686 = 14'h42 == field_data_lo_135 ? _field_data_T_1060 : _GEN_2685; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2687 = 14'h43 == field_data_lo_135 ? _field_data_T_1061 : _GEN_2686; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2688 = 14'h44 == field_data_lo_135 ? _field_data_T_1062 : _GEN_2687; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2689 = 14'h45 == field_data_lo_135 ? _field_data_T_1063 : _GEN_2688; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_56 = vliw_56[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_156 = vliw_56[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_56 = field_data_lo_156[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_56 = field_data_lo_156[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_104 = {{1'd0}, args_offset_56}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_104 = _total_offset_T_104[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2693 = 3'h1 == total_offset_104 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2694 = 3'h2 == total_offset_104 ? args_2 : _GEN_2693; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2695 = 3'h3 == total_offset_104 ? args_3 : _GEN_2694; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2696 = 3'h4 == total_offset_104 ? args_4 : _GEN_2695; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2697 = 3'h5 == total_offset_104 ? args_5 : _GEN_2696; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2698 = 3'h6 == total_offset_104 ? args_6 : _GEN_2697; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2699 = total_offset_104 < 3'h7 ? _GEN_2698 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_56_3 = 3'h0 < args_length_56 ? _GEN_2699 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_105 = args_offset_56 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2702 = 3'h1 == total_offset_105 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2703 = 3'h2 == total_offset_105 ? args_2 : _GEN_2702; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2704 = 3'h3 == total_offset_105 ? args_3 : _GEN_2703; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2705 = 3'h4 == total_offset_105 ? args_4 : _GEN_2704; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2706 = 3'h5 == total_offset_105 ? args_5 : _GEN_2705; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2707 = 3'h6 == total_offset_105 ? args_6 : _GEN_2706; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2708 = total_offset_105 < 3'h7 ? _GEN_2707 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_56_2 = 3'h1 < args_length_56 ? _GEN_2708 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_106 = args_offset_56 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2711 = 3'h1 == total_offset_106 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2712 = 3'h2 == total_offset_106 ? args_2 : _GEN_2711; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2713 = 3'h3 == total_offset_106 ? args_3 : _GEN_2712; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2714 = 3'h4 == total_offset_106 ? args_4 : _GEN_2713; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2715 = 3'h5 == total_offset_106 ? args_5 : _GEN_2714; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2716 = 3'h6 == total_offset_106 ? args_6 : _GEN_2715; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2717 = total_offset_106 < 3'h7 ? _GEN_2716 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_56_1 = 3'h2 < args_length_56 ? _GEN_2717 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_107 = args_offset_56 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2720 = 3'h1 == total_offset_107 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2721 = 3'h2 == total_offset_107 ? args_2 : _GEN_2720; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2722 = 3'h3 == total_offset_107 ? args_3 : _GEN_2721; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2723 = 3'h4 == total_offset_107 ? args_4 : _GEN_2722; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2724 = 3'h5 == total_offset_107 ? args_5 : _GEN_2723; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2725 = 3'h6 == total_offset_107 ? args_6 : _GEN_2724; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2726 = total_offset_107 < 3'h7 ? _GEN_2725 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_56_0 = 3'h3 < args_length_56 ? _GEN_2726 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1184 = {field_bytes_56_0,field_bytes_56_1,field_bytes_56_2,field_bytes_56_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2728 = opcode_56 == 4'ha ? _field_data_T_1184 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2729 = opcode_56 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1917 = opcode_56 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_170 = field_data_lo_156[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1187 = {field_data_hi_170,field_data_lo_156}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_113 = _T_1917 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2730 = opcode_56 == 4'h8 | opcode_56 == 4'hb ? _field_data_T_1187 : _GEN_2728; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2731 = opcode_56 == 4'h8 | opcode_56 == 4'hb ? _field_tag_T_113 : _GEN_2729; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2732 = 14'h32 == field_data_lo_156 ? _field_data_T_1044 : _GEN_2730; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2733 = 14'h33 == field_data_lo_156 ? _field_data_T_1045 : _GEN_2732; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2734 = 14'h34 == field_data_lo_156 ? _field_data_T_1046 : _GEN_2733; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2735 = 14'h35 == field_data_lo_156 ? _field_data_T_1047 : _GEN_2734; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2736 = 14'h36 == field_data_lo_156 ? _field_data_T_1048 : _GEN_2735; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2737 = 14'h37 == field_data_lo_156 ? _field_data_T_1049 : _GEN_2736; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2738 = 14'h38 == field_data_lo_156 ? _field_data_T_1050 : _GEN_2737; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2739 = 14'h39 == field_data_lo_156 ? _field_data_T_1051 : _GEN_2738; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2740 = 14'h3a == field_data_lo_156 ? _field_data_T_1052 : _GEN_2739; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2741 = 14'h3b == field_data_lo_156 ? _field_data_T_1053 : _GEN_2740; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2742 = 14'h3c == field_data_lo_156 ? _field_data_T_1054 : _GEN_2741; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2743 = 14'h3d == field_data_lo_156 ? _field_data_T_1055 : _GEN_2742; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2744 = 14'h3e == field_data_lo_156 ? _field_data_T_1056 : _GEN_2743; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2745 = 14'h3f == field_data_lo_156 ? _field_data_T_1057 : _GEN_2744; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2746 = 14'h40 == field_data_lo_156 ? _field_data_T_1058 : _GEN_2745; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2747 = 14'h41 == field_data_lo_156 ? _field_data_T_1059 : _GEN_2746; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2748 = 14'h42 == field_data_lo_156 ? _field_data_T_1060 : _GEN_2747; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2749 = 14'h43 == field_data_lo_156 ? _field_data_T_1061 : _GEN_2748; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2750 = 14'h44 == field_data_lo_156 ? _field_data_T_1062 : _GEN_2749; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2751 = 14'h45 == field_data_lo_156 ? _field_data_T_1063 : _GEN_2750; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_57 = vliw_57[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_177 = vliw_57[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_57 = field_data_lo_177[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_57 = field_data_lo_177[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_108 = {{1'd0}, args_offset_57}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_108 = _total_offset_T_108[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2755 = 3'h1 == total_offset_108 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2756 = 3'h2 == total_offset_108 ? args_2 : _GEN_2755; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2757 = 3'h3 == total_offset_108 ? args_3 : _GEN_2756; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2758 = 3'h4 == total_offset_108 ? args_4 : _GEN_2757; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2759 = 3'h5 == total_offset_108 ? args_5 : _GEN_2758; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2760 = 3'h6 == total_offset_108 ? args_6 : _GEN_2759; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2761 = total_offset_108 < 3'h7 ? _GEN_2760 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_57_3 = 3'h0 < args_length_57 ? _GEN_2761 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_109 = args_offset_57 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2764 = 3'h1 == total_offset_109 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2765 = 3'h2 == total_offset_109 ? args_2 : _GEN_2764; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2766 = 3'h3 == total_offset_109 ? args_3 : _GEN_2765; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2767 = 3'h4 == total_offset_109 ? args_4 : _GEN_2766; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2768 = 3'h5 == total_offset_109 ? args_5 : _GEN_2767; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2769 = 3'h6 == total_offset_109 ? args_6 : _GEN_2768; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2770 = total_offset_109 < 3'h7 ? _GEN_2769 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_57_2 = 3'h1 < args_length_57 ? _GEN_2770 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_110 = args_offset_57 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2773 = 3'h1 == total_offset_110 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2774 = 3'h2 == total_offset_110 ? args_2 : _GEN_2773; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2775 = 3'h3 == total_offset_110 ? args_3 : _GEN_2774; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2776 = 3'h4 == total_offset_110 ? args_4 : _GEN_2775; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2777 = 3'h5 == total_offset_110 ? args_5 : _GEN_2776; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2778 = 3'h6 == total_offset_110 ? args_6 : _GEN_2777; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2779 = total_offset_110 < 3'h7 ? _GEN_2778 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_57_1 = 3'h2 < args_length_57 ? _GEN_2779 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_111 = args_offset_57 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2782 = 3'h1 == total_offset_111 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2783 = 3'h2 == total_offset_111 ? args_2 : _GEN_2782; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2784 = 3'h3 == total_offset_111 ? args_3 : _GEN_2783; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2785 = 3'h4 == total_offset_111 ? args_4 : _GEN_2784; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2786 = 3'h5 == total_offset_111 ? args_5 : _GEN_2785; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2787 = 3'h6 == total_offset_111 ? args_6 : _GEN_2786; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2788 = total_offset_111 < 3'h7 ? _GEN_2787 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_57_0 = 3'h3 < args_length_57 ? _GEN_2788 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1208 = {field_bytes_57_0,field_bytes_57_1,field_bytes_57_2,field_bytes_57_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2790 = opcode_57 == 4'ha ? _field_data_T_1208 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2791 = opcode_57 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1950 = opcode_57 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_193 = field_data_lo_177[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1211 = {field_data_hi_193,field_data_lo_177}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_115 = _T_1950 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2792 = opcode_57 == 4'h8 | opcode_57 == 4'hb ? _field_data_T_1211 : _GEN_2790; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2793 = opcode_57 == 4'h8 | opcode_57 == 4'hb ? _field_tag_T_115 : _GEN_2791; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2794 = 14'h32 == field_data_lo_177 ? _field_data_T_1044 : _GEN_2792; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2795 = 14'h33 == field_data_lo_177 ? _field_data_T_1045 : _GEN_2794; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2796 = 14'h34 == field_data_lo_177 ? _field_data_T_1046 : _GEN_2795; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2797 = 14'h35 == field_data_lo_177 ? _field_data_T_1047 : _GEN_2796; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2798 = 14'h36 == field_data_lo_177 ? _field_data_T_1048 : _GEN_2797; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2799 = 14'h37 == field_data_lo_177 ? _field_data_T_1049 : _GEN_2798; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2800 = 14'h38 == field_data_lo_177 ? _field_data_T_1050 : _GEN_2799; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2801 = 14'h39 == field_data_lo_177 ? _field_data_T_1051 : _GEN_2800; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2802 = 14'h3a == field_data_lo_177 ? _field_data_T_1052 : _GEN_2801; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2803 = 14'h3b == field_data_lo_177 ? _field_data_T_1053 : _GEN_2802; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2804 = 14'h3c == field_data_lo_177 ? _field_data_T_1054 : _GEN_2803; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2805 = 14'h3d == field_data_lo_177 ? _field_data_T_1055 : _GEN_2804; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2806 = 14'h3e == field_data_lo_177 ? _field_data_T_1056 : _GEN_2805; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2807 = 14'h3f == field_data_lo_177 ? _field_data_T_1057 : _GEN_2806; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2808 = 14'h40 == field_data_lo_177 ? _field_data_T_1058 : _GEN_2807; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2809 = 14'h41 == field_data_lo_177 ? _field_data_T_1059 : _GEN_2808; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2810 = 14'h42 == field_data_lo_177 ? _field_data_T_1060 : _GEN_2809; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2811 = 14'h43 == field_data_lo_177 ? _field_data_T_1061 : _GEN_2810; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2812 = 14'h44 == field_data_lo_177 ? _field_data_T_1062 : _GEN_2811; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2813 = 14'h45 == field_data_lo_177 ? _field_data_T_1063 : _GEN_2812; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_58 = vliw_58[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_198 = vliw_58[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_58 = field_data_lo_198[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_58 = field_data_lo_198[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_112 = {{1'd0}, args_offset_58}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_112 = _total_offset_T_112[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2817 = 3'h1 == total_offset_112 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2818 = 3'h2 == total_offset_112 ? args_2 : _GEN_2817; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2819 = 3'h3 == total_offset_112 ? args_3 : _GEN_2818; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2820 = 3'h4 == total_offset_112 ? args_4 : _GEN_2819; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2821 = 3'h5 == total_offset_112 ? args_5 : _GEN_2820; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2822 = 3'h6 == total_offset_112 ? args_6 : _GEN_2821; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2823 = total_offset_112 < 3'h7 ? _GEN_2822 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_58_3 = 3'h0 < args_length_58 ? _GEN_2823 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_113 = args_offset_58 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2826 = 3'h1 == total_offset_113 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2827 = 3'h2 == total_offset_113 ? args_2 : _GEN_2826; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2828 = 3'h3 == total_offset_113 ? args_3 : _GEN_2827; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2829 = 3'h4 == total_offset_113 ? args_4 : _GEN_2828; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2830 = 3'h5 == total_offset_113 ? args_5 : _GEN_2829; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2831 = 3'h6 == total_offset_113 ? args_6 : _GEN_2830; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2832 = total_offset_113 < 3'h7 ? _GEN_2831 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_58_2 = 3'h1 < args_length_58 ? _GEN_2832 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_114 = args_offset_58 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2835 = 3'h1 == total_offset_114 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2836 = 3'h2 == total_offset_114 ? args_2 : _GEN_2835; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2837 = 3'h3 == total_offset_114 ? args_3 : _GEN_2836; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2838 = 3'h4 == total_offset_114 ? args_4 : _GEN_2837; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2839 = 3'h5 == total_offset_114 ? args_5 : _GEN_2838; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2840 = 3'h6 == total_offset_114 ? args_6 : _GEN_2839; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2841 = total_offset_114 < 3'h7 ? _GEN_2840 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_58_1 = 3'h2 < args_length_58 ? _GEN_2841 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_115 = args_offset_58 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2844 = 3'h1 == total_offset_115 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2845 = 3'h2 == total_offset_115 ? args_2 : _GEN_2844; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2846 = 3'h3 == total_offset_115 ? args_3 : _GEN_2845; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2847 = 3'h4 == total_offset_115 ? args_4 : _GEN_2846; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2848 = 3'h5 == total_offset_115 ? args_5 : _GEN_2847; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2849 = 3'h6 == total_offset_115 ? args_6 : _GEN_2848; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2850 = total_offset_115 < 3'h7 ? _GEN_2849 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_58_0 = 3'h3 < args_length_58 ? _GEN_2850 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1232 = {field_bytes_58_0,field_bytes_58_1,field_bytes_58_2,field_bytes_58_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2852 = opcode_58 == 4'ha ? _field_data_T_1232 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2853 = opcode_58 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_1983 = opcode_58 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_216 = field_data_lo_198[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1235 = {field_data_hi_216,field_data_lo_198}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_117 = _T_1983 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2854 = opcode_58 == 4'h8 | opcode_58 == 4'hb ? _field_data_T_1235 : _GEN_2852; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2855 = opcode_58 == 4'h8 | opcode_58 == 4'hb ? _field_tag_T_117 : _GEN_2853; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2856 = 14'h32 == field_data_lo_198 ? _field_data_T_1044 : _GEN_2854; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2857 = 14'h33 == field_data_lo_198 ? _field_data_T_1045 : _GEN_2856; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2858 = 14'h34 == field_data_lo_198 ? _field_data_T_1046 : _GEN_2857; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2859 = 14'h35 == field_data_lo_198 ? _field_data_T_1047 : _GEN_2858; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2860 = 14'h36 == field_data_lo_198 ? _field_data_T_1048 : _GEN_2859; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2861 = 14'h37 == field_data_lo_198 ? _field_data_T_1049 : _GEN_2860; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2862 = 14'h38 == field_data_lo_198 ? _field_data_T_1050 : _GEN_2861; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2863 = 14'h39 == field_data_lo_198 ? _field_data_T_1051 : _GEN_2862; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2864 = 14'h3a == field_data_lo_198 ? _field_data_T_1052 : _GEN_2863; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2865 = 14'h3b == field_data_lo_198 ? _field_data_T_1053 : _GEN_2864; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2866 = 14'h3c == field_data_lo_198 ? _field_data_T_1054 : _GEN_2865; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2867 = 14'h3d == field_data_lo_198 ? _field_data_T_1055 : _GEN_2866; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2868 = 14'h3e == field_data_lo_198 ? _field_data_T_1056 : _GEN_2867; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2869 = 14'h3f == field_data_lo_198 ? _field_data_T_1057 : _GEN_2868; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2870 = 14'h40 == field_data_lo_198 ? _field_data_T_1058 : _GEN_2869; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2871 = 14'h41 == field_data_lo_198 ? _field_data_T_1059 : _GEN_2870; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2872 = 14'h42 == field_data_lo_198 ? _field_data_T_1060 : _GEN_2871; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2873 = 14'h43 == field_data_lo_198 ? _field_data_T_1061 : _GEN_2872; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2874 = 14'h44 == field_data_lo_198 ? _field_data_T_1062 : _GEN_2873; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2875 = 14'h45 == field_data_lo_198 ? _field_data_T_1063 : _GEN_2874; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_59 = vliw_59[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_219 = vliw_59[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_59 = field_data_lo_219[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_59 = field_data_lo_219[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_116 = {{1'd0}, args_offset_59}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_116 = _total_offset_T_116[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2879 = 3'h1 == total_offset_116 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2880 = 3'h2 == total_offset_116 ? args_2 : _GEN_2879; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2881 = 3'h3 == total_offset_116 ? args_3 : _GEN_2880; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2882 = 3'h4 == total_offset_116 ? args_4 : _GEN_2881; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2883 = 3'h5 == total_offset_116 ? args_5 : _GEN_2882; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2884 = 3'h6 == total_offset_116 ? args_6 : _GEN_2883; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2885 = total_offset_116 < 3'h7 ? _GEN_2884 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_59_3 = 3'h0 < args_length_59 ? _GEN_2885 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_117 = args_offset_59 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2888 = 3'h1 == total_offset_117 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2889 = 3'h2 == total_offset_117 ? args_2 : _GEN_2888; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2890 = 3'h3 == total_offset_117 ? args_3 : _GEN_2889; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2891 = 3'h4 == total_offset_117 ? args_4 : _GEN_2890; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2892 = 3'h5 == total_offset_117 ? args_5 : _GEN_2891; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2893 = 3'h6 == total_offset_117 ? args_6 : _GEN_2892; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2894 = total_offset_117 < 3'h7 ? _GEN_2893 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_59_2 = 3'h1 < args_length_59 ? _GEN_2894 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_118 = args_offset_59 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2897 = 3'h1 == total_offset_118 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2898 = 3'h2 == total_offset_118 ? args_2 : _GEN_2897; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2899 = 3'h3 == total_offset_118 ? args_3 : _GEN_2898; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2900 = 3'h4 == total_offset_118 ? args_4 : _GEN_2899; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2901 = 3'h5 == total_offset_118 ? args_5 : _GEN_2900; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2902 = 3'h6 == total_offset_118 ? args_6 : _GEN_2901; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2903 = total_offset_118 < 3'h7 ? _GEN_2902 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_59_1 = 3'h2 < args_length_59 ? _GEN_2903 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_119 = args_offset_59 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2906 = 3'h1 == total_offset_119 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2907 = 3'h2 == total_offset_119 ? args_2 : _GEN_2906; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2908 = 3'h3 == total_offset_119 ? args_3 : _GEN_2907; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2909 = 3'h4 == total_offset_119 ? args_4 : _GEN_2908; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2910 = 3'h5 == total_offset_119 ? args_5 : _GEN_2909; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2911 = 3'h6 == total_offset_119 ? args_6 : _GEN_2910; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2912 = total_offset_119 < 3'h7 ? _GEN_2911 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_59_0 = 3'h3 < args_length_59 ? _GEN_2912 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1256 = {field_bytes_59_0,field_bytes_59_1,field_bytes_59_2,field_bytes_59_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2914 = opcode_59 == 4'ha ? _field_data_T_1256 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2915 = opcode_59 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2016 = opcode_59 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_239 = field_data_lo_219[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1259 = {field_data_hi_239,field_data_lo_219}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_119 = _T_2016 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2916 = opcode_59 == 4'h8 | opcode_59 == 4'hb ? _field_data_T_1259 : _GEN_2914; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2917 = opcode_59 == 4'h8 | opcode_59 == 4'hb ? _field_tag_T_119 : _GEN_2915; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2918 = 14'h32 == field_data_lo_219 ? _field_data_T_1044 : _GEN_2916; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2919 = 14'h33 == field_data_lo_219 ? _field_data_T_1045 : _GEN_2918; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2920 = 14'h34 == field_data_lo_219 ? _field_data_T_1046 : _GEN_2919; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2921 = 14'h35 == field_data_lo_219 ? _field_data_T_1047 : _GEN_2920; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2922 = 14'h36 == field_data_lo_219 ? _field_data_T_1048 : _GEN_2921; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2923 = 14'h37 == field_data_lo_219 ? _field_data_T_1049 : _GEN_2922; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2924 = 14'h38 == field_data_lo_219 ? _field_data_T_1050 : _GEN_2923; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2925 = 14'h39 == field_data_lo_219 ? _field_data_T_1051 : _GEN_2924; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2926 = 14'h3a == field_data_lo_219 ? _field_data_T_1052 : _GEN_2925; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2927 = 14'h3b == field_data_lo_219 ? _field_data_T_1053 : _GEN_2926; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2928 = 14'h3c == field_data_lo_219 ? _field_data_T_1054 : _GEN_2927; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2929 = 14'h3d == field_data_lo_219 ? _field_data_T_1055 : _GEN_2928; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2930 = 14'h3e == field_data_lo_219 ? _field_data_T_1056 : _GEN_2929; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2931 = 14'h3f == field_data_lo_219 ? _field_data_T_1057 : _GEN_2930; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2932 = 14'h40 == field_data_lo_219 ? _field_data_T_1058 : _GEN_2931; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2933 = 14'h41 == field_data_lo_219 ? _field_data_T_1059 : _GEN_2932; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2934 = 14'h42 == field_data_lo_219 ? _field_data_T_1060 : _GEN_2933; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2935 = 14'h43 == field_data_lo_219 ? _field_data_T_1061 : _GEN_2934; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2936 = 14'h44 == field_data_lo_219 ? _field_data_T_1062 : _GEN_2935; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2937 = 14'h45 == field_data_lo_219 ? _field_data_T_1063 : _GEN_2936; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_60 = vliw_60[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_240 = vliw_60[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_60 = field_data_lo_240[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_60 = field_data_lo_240[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_120 = {{1'd0}, args_offset_60}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_120 = _total_offset_T_120[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2941 = 3'h1 == total_offset_120 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2942 = 3'h2 == total_offset_120 ? args_2 : _GEN_2941; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2943 = 3'h3 == total_offset_120 ? args_3 : _GEN_2942; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2944 = 3'h4 == total_offset_120 ? args_4 : _GEN_2943; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2945 = 3'h5 == total_offset_120 ? args_5 : _GEN_2944; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2946 = 3'h6 == total_offset_120 ? args_6 : _GEN_2945; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2947 = total_offset_120 < 3'h7 ? _GEN_2946 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_60_3 = 3'h0 < args_length_60 ? _GEN_2947 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_121 = args_offset_60 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2950 = 3'h1 == total_offset_121 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2951 = 3'h2 == total_offset_121 ? args_2 : _GEN_2950; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2952 = 3'h3 == total_offset_121 ? args_3 : _GEN_2951; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2953 = 3'h4 == total_offset_121 ? args_4 : _GEN_2952; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2954 = 3'h5 == total_offset_121 ? args_5 : _GEN_2953; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2955 = 3'h6 == total_offset_121 ? args_6 : _GEN_2954; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2956 = total_offset_121 < 3'h7 ? _GEN_2955 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_60_2 = 3'h1 < args_length_60 ? _GEN_2956 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_122 = args_offset_60 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2959 = 3'h1 == total_offset_122 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2960 = 3'h2 == total_offset_122 ? args_2 : _GEN_2959; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2961 = 3'h3 == total_offset_122 ? args_3 : _GEN_2960; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2962 = 3'h4 == total_offset_122 ? args_4 : _GEN_2961; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2963 = 3'h5 == total_offset_122 ? args_5 : _GEN_2962; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2964 = 3'h6 == total_offset_122 ? args_6 : _GEN_2963; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2965 = total_offset_122 < 3'h7 ? _GEN_2964 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_60_1 = 3'h2 < args_length_60 ? _GEN_2965 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_123 = args_offset_60 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_2968 = 3'h1 == total_offset_123 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2969 = 3'h2 == total_offset_123 ? args_2 : _GEN_2968; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2970 = 3'h3 == total_offset_123 ? args_3 : _GEN_2969; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2971 = 3'h4 == total_offset_123 ? args_4 : _GEN_2970; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2972 = 3'h5 == total_offset_123 ? args_5 : _GEN_2971; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2973 = 3'h6 == total_offset_123 ? args_6 : _GEN_2972; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_2974 = total_offset_123 < 3'h7 ? _GEN_2973 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_60_0 = 3'h3 < args_length_60 ? _GEN_2974 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1280 = {field_bytes_60_0,field_bytes_60_1,field_bytes_60_2,field_bytes_60_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2976 = opcode_60 == 4'ha ? _field_data_T_1280 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_2977 = opcode_60 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2049 = opcode_60 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_262 = field_data_lo_240[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1283 = {field_data_hi_262,field_data_lo_240}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_121 = _T_2049 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_2978 = opcode_60 == 4'h8 | opcode_60 == 4'hb ? _field_data_T_1283 : _GEN_2976; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_2979 = opcode_60 == 4'h8 | opcode_60 == 4'hb ? _field_tag_T_121 : _GEN_2977; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_2980 = 14'h32 == field_data_lo_240 ? _field_data_T_1044 : _GEN_2978; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2981 = 14'h33 == field_data_lo_240 ? _field_data_T_1045 : _GEN_2980; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2982 = 14'h34 == field_data_lo_240 ? _field_data_T_1046 : _GEN_2981; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2983 = 14'h35 == field_data_lo_240 ? _field_data_T_1047 : _GEN_2982; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2984 = 14'h36 == field_data_lo_240 ? _field_data_T_1048 : _GEN_2983; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2985 = 14'h37 == field_data_lo_240 ? _field_data_T_1049 : _GEN_2984; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2986 = 14'h38 == field_data_lo_240 ? _field_data_T_1050 : _GEN_2985; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2987 = 14'h39 == field_data_lo_240 ? _field_data_T_1051 : _GEN_2986; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2988 = 14'h3a == field_data_lo_240 ? _field_data_T_1052 : _GEN_2987; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2989 = 14'h3b == field_data_lo_240 ? _field_data_T_1053 : _GEN_2988; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2990 = 14'h3c == field_data_lo_240 ? _field_data_T_1054 : _GEN_2989; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2991 = 14'h3d == field_data_lo_240 ? _field_data_T_1055 : _GEN_2990; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2992 = 14'h3e == field_data_lo_240 ? _field_data_T_1056 : _GEN_2991; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2993 = 14'h3f == field_data_lo_240 ? _field_data_T_1057 : _GEN_2992; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2994 = 14'h40 == field_data_lo_240 ? _field_data_T_1058 : _GEN_2993; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2995 = 14'h41 == field_data_lo_240 ? _field_data_T_1059 : _GEN_2994; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2996 = 14'h42 == field_data_lo_240 ? _field_data_T_1060 : _GEN_2995; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2997 = 14'h43 == field_data_lo_240 ? _field_data_T_1061 : _GEN_2996; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2998 = 14'h44 == field_data_lo_240 ? _field_data_T_1062 : _GEN_2997; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_2999 = 14'h45 == field_data_lo_240 ? _field_data_T_1063 : _GEN_2998; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_61 = vliw_61[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_261 = vliw_61[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_61 = field_data_lo_261[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_61 = field_data_lo_261[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_124 = {{1'd0}, args_offset_61}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_124 = _total_offset_T_124[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3003 = 3'h1 == total_offset_124 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3004 = 3'h2 == total_offset_124 ? args_2 : _GEN_3003; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3005 = 3'h3 == total_offset_124 ? args_3 : _GEN_3004; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3006 = 3'h4 == total_offset_124 ? args_4 : _GEN_3005; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3007 = 3'h5 == total_offset_124 ? args_5 : _GEN_3006; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3008 = 3'h6 == total_offset_124 ? args_6 : _GEN_3007; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3009 = total_offset_124 < 3'h7 ? _GEN_3008 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_61_3 = 3'h0 < args_length_61 ? _GEN_3009 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_125 = args_offset_61 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3012 = 3'h1 == total_offset_125 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3013 = 3'h2 == total_offset_125 ? args_2 : _GEN_3012; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3014 = 3'h3 == total_offset_125 ? args_3 : _GEN_3013; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3015 = 3'h4 == total_offset_125 ? args_4 : _GEN_3014; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3016 = 3'h5 == total_offset_125 ? args_5 : _GEN_3015; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3017 = 3'h6 == total_offset_125 ? args_6 : _GEN_3016; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3018 = total_offset_125 < 3'h7 ? _GEN_3017 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_61_2 = 3'h1 < args_length_61 ? _GEN_3018 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_126 = args_offset_61 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3021 = 3'h1 == total_offset_126 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3022 = 3'h2 == total_offset_126 ? args_2 : _GEN_3021; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3023 = 3'h3 == total_offset_126 ? args_3 : _GEN_3022; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3024 = 3'h4 == total_offset_126 ? args_4 : _GEN_3023; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3025 = 3'h5 == total_offset_126 ? args_5 : _GEN_3024; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3026 = 3'h6 == total_offset_126 ? args_6 : _GEN_3025; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3027 = total_offset_126 < 3'h7 ? _GEN_3026 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_61_1 = 3'h2 < args_length_61 ? _GEN_3027 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_127 = args_offset_61 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3030 = 3'h1 == total_offset_127 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3031 = 3'h2 == total_offset_127 ? args_2 : _GEN_3030; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3032 = 3'h3 == total_offset_127 ? args_3 : _GEN_3031; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3033 = 3'h4 == total_offset_127 ? args_4 : _GEN_3032; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3034 = 3'h5 == total_offset_127 ? args_5 : _GEN_3033; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3035 = 3'h6 == total_offset_127 ? args_6 : _GEN_3034; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3036 = total_offset_127 < 3'h7 ? _GEN_3035 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_61_0 = 3'h3 < args_length_61 ? _GEN_3036 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1304 = {field_bytes_61_0,field_bytes_61_1,field_bytes_61_2,field_bytes_61_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3038 = opcode_61 == 4'ha ? _field_data_T_1304 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3039 = opcode_61 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2082 = opcode_61 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_285 = field_data_lo_261[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1307 = {field_data_hi_285,field_data_lo_261}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_123 = _T_2082 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3040 = opcode_61 == 4'h8 | opcode_61 == 4'hb ? _field_data_T_1307 : _GEN_3038; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3041 = opcode_61 == 4'h8 | opcode_61 == 4'hb ? _field_tag_T_123 : _GEN_3039; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3042 = 14'h32 == field_data_lo_261 ? _field_data_T_1044 : _GEN_3040; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3043 = 14'h33 == field_data_lo_261 ? _field_data_T_1045 : _GEN_3042; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3044 = 14'h34 == field_data_lo_261 ? _field_data_T_1046 : _GEN_3043; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3045 = 14'h35 == field_data_lo_261 ? _field_data_T_1047 : _GEN_3044; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3046 = 14'h36 == field_data_lo_261 ? _field_data_T_1048 : _GEN_3045; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3047 = 14'h37 == field_data_lo_261 ? _field_data_T_1049 : _GEN_3046; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3048 = 14'h38 == field_data_lo_261 ? _field_data_T_1050 : _GEN_3047; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3049 = 14'h39 == field_data_lo_261 ? _field_data_T_1051 : _GEN_3048; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3050 = 14'h3a == field_data_lo_261 ? _field_data_T_1052 : _GEN_3049; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3051 = 14'h3b == field_data_lo_261 ? _field_data_T_1053 : _GEN_3050; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3052 = 14'h3c == field_data_lo_261 ? _field_data_T_1054 : _GEN_3051; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3053 = 14'h3d == field_data_lo_261 ? _field_data_T_1055 : _GEN_3052; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3054 = 14'h3e == field_data_lo_261 ? _field_data_T_1056 : _GEN_3053; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3055 = 14'h3f == field_data_lo_261 ? _field_data_T_1057 : _GEN_3054; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3056 = 14'h40 == field_data_lo_261 ? _field_data_T_1058 : _GEN_3055; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3057 = 14'h41 == field_data_lo_261 ? _field_data_T_1059 : _GEN_3056; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3058 = 14'h42 == field_data_lo_261 ? _field_data_T_1060 : _GEN_3057; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3059 = 14'h43 == field_data_lo_261 ? _field_data_T_1061 : _GEN_3058; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3060 = 14'h44 == field_data_lo_261 ? _field_data_T_1062 : _GEN_3059; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3061 = 14'h45 == field_data_lo_261 ? _field_data_T_1063 : _GEN_3060; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_62 = vliw_62[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_282 = vliw_62[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_62 = field_data_lo_282[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_62 = field_data_lo_282[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_128 = {{1'd0}, args_offset_62}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_128 = _total_offset_T_128[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3065 = 3'h1 == total_offset_128 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3066 = 3'h2 == total_offset_128 ? args_2 : _GEN_3065; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3067 = 3'h3 == total_offset_128 ? args_3 : _GEN_3066; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3068 = 3'h4 == total_offset_128 ? args_4 : _GEN_3067; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3069 = 3'h5 == total_offset_128 ? args_5 : _GEN_3068; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3070 = 3'h6 == total_offset_128 ? args_6 : _GEN_3069; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3071 = total_offset_128 < 3'h7 ? _GEN_3070 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_62_3 = 3'h0 < args_length_62 ? _GEN_3071 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_129 = args_offset_62 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3074 = 3'h1 == total_offset_129 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3075 = 3'h2 == total_offset_129 ? args_2 : _GEN_3074; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3076 = 3'h3 == total_offset_129 ? args_3 : _GEN_3075; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3077 = 3'h4 == total_offset_129 ? args_4 : _GEN_3076; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3078 = 3'h5 == total_offset_129 ? args_5 : _GEN_3077; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3079 = 3'h6 == total_offset_129 ? args_6 : _GEN_3078; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3080 = total_offset_129 < 3'h7 ? _GEN_3079 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_62_2 = 3'h1 < args_length_62 ? _GEN_3080 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_130 = args_offset_62 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3083 = 3'h1 == total_offset_130 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3084 = 3'h2 == total_offset_130 ? args_2 : _GEN_3083; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3085 = 3'h3 == total_offset_130 ? args_3 : _GEN_3084; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3086 = 3'h4 == total_offset_130 ? args_4 : _GEN_3085; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3087 = 3'h5 == total_offset_130 ? args_5 : _GEN_3086; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3088 = 3'h6 == total_offset_130 ? args_6 : _GEN_3087; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3089 = total_offset_130 < 3'h7 ? _GEN_3088 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_62_1 = 3'h2 < args_length_62 ? _GEN_3089 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_131 = args_offset_62 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3092 = 3'h1 == total_offset_131 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3093 = 3'h2 == total_offset_131 ? args_2 : _GEN_3092; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3094 = 3'h3 == total_offset_131 ? args_3 : _GEN_3093; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3095 = 3'h4 == total_offset_131 ? args_4 : _GEN_3094; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3096 = 3'h5 == total_offset_131 ? args_5 : _GEN_3095; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3097 = 3'h6 == total_offset_131 ? args_6 : _GEN_3096; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3098 = total_offset_131 < 3'h7 ? _GEN_3097 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_62_0 = 3'h3 < args_length_62 ? _GEN_3098 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1328 = {field_bytes_62_0,field_bytes_62_1,field_bytes_62_2,field_bytes_62_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3100 = opcode_62 == 4'ha ? _field_data_T_1328 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3101 = opcode_62 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2115 = opcode_62 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_308 = field_data_lo_282[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1331 = {field_data_hi_308,field_data_lo_282}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_125 = _T_2115 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3102 = opcode_62 == 4'h8 | opcode_62 == 4'hb ? _field_data_T_1331 : _GEN_3100; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3103 = opcode_62 == 4'h8 | opcode_62 == 4'hb ? _field_tag_T_125 : _GEN_3101; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3104 = 14'h32 == field_data_lo_282 ? _field_data_T_1044 : _GEN_3102; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3105 = 14'h33 == field_data_lo_282 ? _field_data_T_1045 : _GEN_3104; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3106 = 14'h34 == field_data_lo_282 ? _field_data_T_1046 : _GEN_3105; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3107 = 14'h35 == field_data_lo_282 ? _field_data_T_1047 : _GEN_3106; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3108 = 14'h36 == field_data_lo_282 ? _field_data_T_1048 : _GEN_3107; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3109 = 14'h37 == field_data_lo_282 ? _field_data_T_1049 : _GEN_3108; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3110 = 14'h38 == field_data_lo_282 ? _field_data_T_1050 : _GEN_3109; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3111 = 14'h39 == field_data_lo_282 ? _field_data_T_1051 : _GEN_3110; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3112 = 14'h3a == field_data_lo_282 ? _field_data_T_1052 : _GEN_3111; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3113 = 14'h3b == field_data_lo_282 ? _field_data_T_1053 : _GEN_3112; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3114 = 14'h3c == field_data_lo_282 ? _field_data_T_1054 : _GEN_3113; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3115 = 14'h3d == field_data_lo_282 ? _field_data_T_1055 : _GEN_3114; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3116 = 14'h3e == field_data_lo_282 ? _field_data_T_1056 : _GEN_3115; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3117 = 14'h3f == field_data_lo_282 ? _field_data_T_1057 : _GEN_3116; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3118 = 14'h40 == field_data_lo_282 ? _field_data_T_1058 : _GEN_3117; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3119 = 14'h41 == field_data_lo_282 ? _field_data_T_1059 : _GEN_3118; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3120 = 14'h42 == field_data_lo_282 ? _field_data_T_1060 : _GEN_3119; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3121 = 14'h43 == field_data_lo_282 ? _field_data_T_1061 : _GEN_3120; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3122 = 14'h44 == field_data_lo_282 ? _field_data_T_1062 : _GEN_3121; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3123 = 14'h45 == field_data_lo_282 ? _field_data_T_1063 : _GEN_3122; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_63 = vliw_63[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_303 = vliw_63[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_63 = field_data_lo_303[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_63 = field_data_lo_303[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_132 = {{1'd0}, args_offset_63}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_132 = _total_offset_T_132[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3127 = 3'h1 == total_offset_132 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3128 = 3'h2 == total_offset_132 ? args_2 : _GEN_3127; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3129 = 3'h3 == total_offset_132 ? args_3 : _GEN_3128; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3130 = 3'h4 == total_offset_132 ? args_4 : _GEN_3129; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3131 = 3'h5 == total_offset_132 ? args_5 : _GEN_3130; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3132 = 3'h6 == total_offset_132 ? args_6 : _GEN_3131; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3133 = total_offset_132 < 3'h7 ? _GEN_3132 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_63_3 = 3'h0 < args_length_63 ? _GEN_3133 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_133 = args_offset_63 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3136 = 3'h1 == total_offset_133 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3137 = 3'h2 == total_offset_133 ? args_2 : _GEN_3136; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3138 = 3'h3 == total_offset_133 ? args_3 : _GEN_3137; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3139 = 3'h4 == total_offset_133 ? args_4 : _GEN_3138; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3140 = 3'h5 == total_offset_133 ? args_5 : _GEN_3139; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3141 = 3'h6 == total_offset_133 ? args_6 : _GEN_3140; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3142 = total_offset_133 < 3'h7 ? _GEN_3141 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_63_2 = 3'h1 < args_length_63 ? _GEN_3142 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_134 = args_offset_63 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3145 = 3'h1 == total_offset_134 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3146 = 3'h2 == total_offset_134 ? args_2 : _GEN_3145; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3147 = 3'h3 == total_offset_134 ? args_3 : _GEN_3146; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3148 = 3'h4 == total_offset_134 ? args_4 : _GEN_3147; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3149 = 3'h5 == total_offset_134 ? args_5 : _GEN_3148; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3150 = 3'h6 == total_offset_134 ? args_6 : _GEN_3149; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3151 = total_offset_134 < 3'h7 ? _GEN_3150 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_63_1 = 3'h2 < args_length_63 ? _GEN_3151 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_135 = args_offset_63 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3154 = 3'h1 == total_offset_135 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3155 = 3'h2 == total_offset_135 ? args_2 : _GEN_3154; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3156 = 3'h3 == total_offset_135 ? args_3 : _GEN_3155; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3157 = 3'h4 == total_offset_135 ? args_4 : _GEN_3156; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3158 = 3'h5 == total_offset_135 ? args_5 : _GEN_3157; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3159 = 3'h6 == total_offset_135 ? args_6 : _GEN_3158; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3160 = total_offset_135 < 3'h7 ? _GEN_3159 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_63_0 = 3'h3 < args_length_63 ? _GEN_3160 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1352 = {field_bytes_63_0,field_bytes_63_1,field_bytes_63_2,field_bytes_63_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3162 = opcode_63 == 4'ha ? _field_data_T_1352 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3163 = opcode_63 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2148 = opcode_63 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_331 = field_data_lo_303[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1355 = {field_data_hi_331,field_data_lo_303}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_127 = _T_2148 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3164 = opcode_63 == 4'h8 | opcode_63 == 4'hb ? _field_data_T_1355 : _GEN_3162; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3165 = opcode_63 == 4'h8 | opcode_63 == 4'hb ? _field_tag_T_127 : _GEN_3163; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3166 = 14'h32 == field_data_lo_303 ? _field_data_T_1044 : _GEN_3164; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3167 = 14'h33 == field_data_lo_303 ? _field_data_T_1045 : _GEN_3166; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3168 = 14'h34 == field_data_lo_303 ? _field_data_T_1046 : _GEN_3167; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3169 = 14'h35 == field_data_lo_303 ? _field_data_T_1047 : _GEN_3168; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3170 = 14'h36 == field_data_lo_303 ? _field_data_T_1048 : _GEN_3169; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3171 = 14'h37 == field_data_lo_303 ? _field_data_T_1049 : _GEN_3170; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3172 = 14'h38 == field_data_lo_303 ? _field_data_T_1050 : _GEN_3171; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3173 = 14'h39 == field_data_lo_303 ? _field_data_T_1051 : _GEN_3172; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3174 = 14'h3a == field_data_lo_303 ? _field_data_T_1052 : _GEN_3173; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3175 = 14'h3b == field_data_lo_303 ? _field_data_T_1053 : _GEN_3174; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3176 = 14'h3c == field_data_lo_303 ? _field_data_T_1054 : _GEN_3175; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3177 = 14'h3d == field_data_lo_303 ? _field_data_T_1055 : _GEN_3176; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3178 = 14'h3e == field_data_lo_303 ? _field_data_T_1056 : _GEN_3177; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3179 = 14'h3f == field_data_lo_303 ? _field_data_T_1057 : _GEN_3178; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3180 = 14'h40 == field_data_lo_303 ? _field_data_T_1058 : _GEN_3179; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3181 = 14'h41 == field_data_lo_303 ? _field_data_T_1059 : _GEN_3180; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3182 = 14'h42 == field_data_lo_303 ? _field_data_T_1060 : _GEN_3181; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3183 = 14'h43 == field_data_lo_303 ? _field_data_T_1061 : _GEN_3182; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3184 = 14'h44 == field_data_lo_303 ? _field_data_T_1062 : _GEN_3183; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3185 = 14'h45 == field_data_lo_303 ? _field_data_T_1063 : _GEN_3184; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_64 = vliw_64[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_324 = vliw_64[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_64 = field_data_lo_324[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_64 = field_data_lo_324[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_136 = {{1'd0}, args_offset_64}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_136 = _total_offset_T_136[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3189 = 3'h1 == total_offset_136 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3190 = 3'h2 == total_offset_136 ? args_2 : _GEN_3189; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3191 = 3'h3 == total_offset_136 ? args_3 : _GEN_3190; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3192 = 3'h4 == total_offset_136 ? args_4 : _GEN_3191; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3193 = 3'h5 == total_offset_136 ? args_5 : _GEN_3192; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3194 = 3'h6 == total_offset_136 ? args_6 : _GEN_3193; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3195 = total_offset_136 < 3'h7 ? _GEN_3194 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_3 = 3'h0 < args_length_64 ? _GEN_3195 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_137 = args_offset_64 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3198 = 3'h1 == total_offset_137 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3199 = 3'h2 == total_offset_137 ? args_2 : _GEN_3198; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3200 = 3'h3 == total_offset_137 ? args_3 : _GEN_3199; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3201 = 3'h4 == total_offset_137 ? args_4 : _GEN_3200; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3202 = 3'h5 == total_offset_137 ? args_5 : _GEN_3201; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3203 = 3'h6 == total_offset_137 ? args_6 : _GEN_3202; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3204 = total_offset_137 < 3'h7 ? _GEN_3203 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_2 = 3'h1 < args_length_64 ? _GEN_3204 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_138 = args_offset_64 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3207 = 3'h1 == total_offset_138 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3208 = 3'h2 == total_offset_138 ? args_2 : _GEN_3207; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3209 = 3'h3 == total_offset_138 ? args_3 : _GEN_3208; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3210 = 3'h4 == total_offset_138 ? args_4 : _GEN_3209; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3211 = 3'h5 == total_offset_138 ? args_5 : _GEN_3210; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3212 = 3'h6 == total_offset_138 ? args_6 : _GEN_3211; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3213 = total_offset_138 < 3'h7 ? _GEN_3212 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_1 = 3'h2 < args_length_64 ? _GEN_3213 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_139 = args_offset_64 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3216 = 3'h1 == total_offset_139 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3217 = 3'h2 == total_offset_139 ? args_2 : _GEN_3216; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3218 = 3'h3 == total_offset_139 ? args_3 : _GEN_3217; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3219 = 3'h4 == total_offset_139 ? args_4 : _GEN_3218; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3220 = 3'h5 == total_offset_139 ? args_5 : _GEN_3219; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3221 = 3'h6 == total_offset_139 ? args_6 : _GEN_3220; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3222 = total_offset_139 < 3'h7 ? _GEN_3221 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_64_0 = 3'h3 < args_length_64 ? _GEN_3222 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1376 = {field_bytes_64_0,field_bytes_64_1,field_bytes_64_2,field_bytes_64_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3224 = opcode_64 == 4'ha ? _field_data_T_1376 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3225 = opcode_64 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2181 = opcode_64 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_354 = field_data_lo_324[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1379 = {field_data_hi_354,field_data_lo_324}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_129 = _T_2181 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3226 = opcode_64 == 4'h8 | opcode_64 == 4'hb ? _field_data_T_1379 : _GEN_3224; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3227 = opcode_64 == 4'h8 | opcode_64 == 4'hb ? _field_tag_T_129 : _GEN_3225; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3228 = 14'h32 == field_data_lo_324 ? _field_data_T_1044 : _GEN_3226; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3229 = 14'h33 == field_data_lo_324 ? _field_data_T_1045 : _GEN_3228; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3230 = 14'h34 == field_data_lo_324 ? _field_data_T_1046 : _GEN_3229; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3231 = 14'h35 == field_data_lo_324 ? _field_data_T_1047 : _GEN_3230; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3232 = 14'h36 == field_data_lo_324 ? _field_data_T_1048 : _GEN_3231; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3233 = 14'h37 == field_data_lo_324 ? _field_data_T_1049 : _GEN_3232; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3234 = 14'h38 == field_data_lo_324 ? _field_data_T_1050 : _GEN_3233; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3235 = 14'h39 == field_data_lo_324 ? _field_data_T_1051 : _GEN_3234; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3236 = 14'h3a == field_data_lo_324 ? _field_data_T_1052 : _GEN_3235; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3237 = 14'h3b == field_data_lo_324 ? _field_data_T_1053 : _GEN_3236; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3238 = 14'h3c == field_data_lo_324 ? _field_data_T_1054 : _GEN_3237; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3239 = 14'h3d == field_data_lo_324 ? _field_data_T_1055 : _GEN_3238; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3240 = 14'h3e == field_data_lo_324 ? _field_data_T_1056 : _GEN_3239; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3241 = 14'h3f == field_data_lo_324 ? _field_data_T_1057 : _GEN_3240; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3242 = 14'h40 == field_data_lo_324 ? _field_data_T_1058 : _GEN_3241; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3243 = 14'h41 == field_data_lo_324 ? _field_data_T_1059 : _GEN_3242; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3244 = 14'h42 == field_data_lo_324 ? _field_data_T_1060 : _GEN_3243; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3245 = 14'h43 == field_data_lo_324 ? _field_data_T_1061 : _GEN_3244; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3246 = 14'h44 == field_data_lo_324 ? _field_data_T_1062 : _GEN_3245; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3247 = 14'h45 == field_data_lo_324 ? _field_data_T_1063 : _GEN_3246; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_65 = vliw_65[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_345 = vliw_65[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_65 = field_data_lo_345[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_65 = field_data_lo_345[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_140 = {{1'd0}, args_offset_65}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_140 = _total_offset_T_140[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3251 = 3'h1 == total_offset_140 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3252 = 3'h2 == total_offset_140 ? args_2 : _GEN_3251; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3253 = 3'h3 == total_offset_140 ? args_3 : _GEN_3252; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3254 = 3'h4 == total_offset_140 ? args_4 : _GEN_3253; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3255 = 3'h5 == total_offset_140 ? args_5 : _GEN_3254; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3256 = 3'h6 == total_offset_140 ? args_6 : _GEN_3255; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3257 = total_offset_140 < 3'h7 ? _GEN_3256 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_3 = 3'h0 < args_length_65 ? _GEN_3257 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_141 = args_offset_65 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3260 = 3'h1 == total_offset_141 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3261 = 3'h2 == total_offset_141 ? args_2 : _GEN_3260; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3262 = 3'h3 == total_offset_141 ? args_3 : _GEN_3261; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3263 = 3'h4 == total_offset_141 ? args_4 : _GEN_3262; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3264 = 3'h5 == total_offset_141 ? args_5 : _GEN_3263; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3265 = 3'h6 == total_offset_141 ? args_6 : _GEN_3264; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3266 = total_offset_141 < 3'h7 ? _GEN_3265 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_2 = 3'h1 < args_length_65 ? _GEN_3266 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_142 = args_offset_65 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3269 = 3'h1 == total_offset_142 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3270 = 3'h2 == total_offset_142 ? args_2 : _GEN_3269; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3271 = 3'h3 == total_offset_142 ? args_3 : _GEN_3270; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3272 = 3'h4 == total_offset_142 ? args_4 : _GEN_3271; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3273 = 3'h5 == total_offset_142 ? args_5 : _GEN_3272; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3274 = 3'h6 == total_offset_142 ? args_6 : _GEN_3273; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3275 = total_offset_142 < 3'h7 ? _GEN_3274 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_1 = 3'h2 < args_length_65 ? _GEN_3275 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_143 = args_offset_65 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3278 = 3'h1 == total_offset_143 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3279 = 3'h2 == total_offset_143 ? args_2 : _GEN_3278; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3280 = 3'h3 == total_offset_143 ? args_3 : _GEN_3279; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3281 = 3'h4 == total_offset_143 ? args_4 : _GEN_3280; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3282 = 3'h5 == total_offset_143 ? args_5 : _GEN_3281; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3283 = 3'h6 == total_offset_143 ? args_6 : _GEN_3282; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3284 = total_offset_143 < 3'h7 ? _GEN_3283 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_65_0 = 3'h3 < args_length_65 ? _GEN_3284 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1400 = {field_bytes_65_0,field_bytes_65_1,field_bytes_65_2,field_bytes_65_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3286 = opcode_65 == 4'ha ? _field_data_T_1400 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3287 = opcode_65 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2214 = opcode_65 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_377 = field_data_lo_345[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1403 = {field_data_hi_377,field_data_lo_345}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_131 = _T_2214 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3288 = opcode_65 == 4'h8 | opcode_65 == 4'hb ? _field_data_T_1403 : _GEN_3286; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3289 = opcode_65 == 4'h8 | opcode_65 == 4'hb ? _field_tag_T_131 : _GEN_3287; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3290 = 14'h32 == field_data_lo_345 ? _field_data_T_1044 : _GEN_3288; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3291 = 14'h33 == field_data_lo_345 ? _field_data_T_1045 : _GEN_3290; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3292 = 14'h34 == field_data_lo_345 ? _field_data_T_1046 : _GEN_3291; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3293 = 14'h35 == field_data_lo_345 ? _field_data_T_1047 : _GEN_3292; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3294 = 14'h36 == field_data_lo_345 ? _field_data_T_1048 : _GEN_3293; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3295 = 14'h37 == field_data_lo_345 ? _field_data_T_1049 : _GEN_3294; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3296 = 14'h38 == field_data_lo_345 ? _field_data_T_1050 : _GEN_3295; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3297 = 14'h39 == field_data_lo_345 ? _field_data_T_1051 : _GEN_3296; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3298 = 14'h3a == field_data_lo_345 ? _field_data_T_1052 : _GEN_3297; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3299 = 14'h3b == field_data_lo_345 ? _field_data_T_1053 : _GEN_3298; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3300 = 14'h3c == field_data_lo_345 ? _field_data_T_1054 : _GEN_3299; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3301 = 14'h3d == field_data_lo_345 ? _field_data_T_1055 : _GEN_3300; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3302 = 14'h3e == field_data_lo_345 ? _field_data_T_1056 : _GEN_3301; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3303 = 14'h3f == field_data_lo_345 ? _field_data_T_1057 : _GEN_3302; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3304 = 14'h40 == field_data_lo_345 ? _field_data_T_1058 : _GEN_3303; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3305 = 14'h41 == field_data_lo_345 ? _field_data_T_1059 : _GEN_3304; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3306 = 14'h42 == field_data_lo_345 ? _field_data_T_1060 : _GEN_3305; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3307 = 14'h43 == field_data_lo_345 ? _field_data_T_1061 : _GEN_3306; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3308 = 14'h44 == field_data_lo_345 ? _field_data_T_1062 : _GEN_3307; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3309 = 14'h45 == field_data_lo_345 ? _field_data_T_1063 : _GEN_3308; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_66 = vliw_66[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_366 = vliw_66[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_66 = field_data_lo_366[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_66 = field_data_lo_366[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_144 = {{1'd0}, args_offset_66}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_144 = _total_offset_T_144[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3313 = 3'h1 == total_offset_144 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3314 = 3'h2 == total_offset_144 ? args_2 : _GEN_3313; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3315 = 3'h3 == total_offset_144 ? args_3 : _GEN_3314; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3316 = 3'h4 == total_offset_144 ? args_4 : _GEN_3315; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3317 = 3'h5 == total_offset_144 ? args_5 : _GEN_3316; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3318 = 3'h6 == total_offset_144 ? args_6 : _GEN_3317; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3319 = total_offset_144 < 3'h7 ? _GEN_3318 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_3 = 3'h0 < args_length_66 ? _GEN_3319 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_145 = args_offset_66 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3322 = 3'h1 == total_offset_145 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3323 = 3'h2 == total_offset_145 ? args_2 : _GEN_3322; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3324 = 3'h3 == total_offset_145 ? args_3 : _GEN_3323; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3325 = 3'h4 == total_offset_145 ? args_4 : _GEN_3324; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3326 = 3'h5 == total_offset_145 ? args_5 : _GEN_3325; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3327 = 3'h6 == total_offset_145 ? args_6 : _GEN_3326; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3328 = total_offset_145 < 3'h7 ? _GEN_3327 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_2 = 3'h1 < args_length_66 ? _GEN_3328 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_146 = args_offset_66 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3331 = 3'h1 == total_offset_146 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3332 = 3'h2 == total_offset_146 ? args_2 : _GEN_3331; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3333 = 3'h3 == total_offset_146 ? args_3 : _GEN_3332; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3334 = 3'h4 == total_offset_146 ? args_4 : _GEN_3333; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3335 = 3'h5 == total_offset_146 ? args_5 : _GEN_3334; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3336 = 3'h6 == total_offset_146 ? args_6 : _GEN_3335; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3337 = total_offset_146 < 3'h7 ? _GEN_3336 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_1 = 3'h2 < args_length_66 ? _GEN_3337 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_147 = args_offset_66 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3340 = 3'h1 == total_offset_147 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3341 = 3'h2 == total_offset_147 ? args_2 : _GEN_3340; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3342 = 3'h3 == total_offset_147 ? args_3 : _GEN_3341; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3343 = 3'h4 == total_offset_147 ? args_4 : _GEN_3342; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3344 = 3'h5 == total_offset_147 ? args_5 : _GEN_3343; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3345 = 3'h6 == total_offset_147 ? args_6 : _GEN_3344; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3346 = total_offset_147 < 3'h7 ? _GEN_3345 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_66_0 = 3'h3 < args_length_66 ? _GEN_3346 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1424 = {field_bytes_66_0,field_bytes_66_1,field_bytes_66_2,field_bytes_66_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3348 = opcode_66 == 4'ha ? _field_data_T_1424 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3349 = opcode_66 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2247 = opcode_66 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_400 = field_data_lo_366[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1427 = {field_data_hi_400,field_data_lo_366}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_133 = _T_2247 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3350 = opcode_66 == 4'h8 | opcode_66 == 4'hb ? _field_data_T_1427 : _GEN_3348; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3351 = opcode_66 == 4'h8 | opcode_66 == 4'hb ? _field_tag_T_133 : _GEN_3349; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3352 = 14'h32 == field_data_lo_366 ? _field_data_T_1044 : _GEN_3350; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3353 = 14'h33 == field_data_lo_366 ? _field_data_T_1045 : _GEN_3352; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3354 = 14'h34 == field_data_lo_366 ? _field_data_T_1046 : _GEN_3353; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3355 = 14'h35 == field_data_lo_366 ? _field_data_T_1047 : _GEN_3354; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3356 = 14'h36 == field_data_lo_366 ? _field_data_T_1048 : _GEN_3355; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3357 = 14'h37 == field_data_lo_366 ? _field_data_T_1049 : _GEN_3356; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3358 = 14'h38 == field_data_lo_366 ? _field_data_T_1050 : _GEN_3357; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3359 = 14'h39 == field_data_lo_366 ? _field_data_T_1051 : _GEN_3358; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3360 = 14'h3a == field_data_lo_366 ? _field_data_T_1052 : _GEN_3359; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3361 = 14'h3b == field_data_lo_366 ? _field_data_T_1053 : _GEN_3360; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3362 = 14'h3c == field_data_lo_366 ? _field_data_T_1054 : _GEN_3361; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3363 = 14'h3d == field_data_lo_366 ? _field_data_T_1055 : _GEN_3362; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3364 = 14'h3e == field_data_lo_366 ? _field_data_T_1056 : _GEN_3363; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3365 = 14'h3f == field_data_lo_366 ? _field_data_T_1057 : _GEN_3364; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3366 = 14'h40 == field_data_lo_366 ? _field_data_T_1058 : _GEN_3365; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3367 = 14'h41 == field_data_lo_366 ? _field_data_T_1059 : _GEN_3366; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3368 = 14'h42 == field_data_lo_366 ? _field_data_T_1060 : _GEN_3367; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3369 = 14'h43 == field_data_lo_366 ? _field_data_T_1061 : _GEN_3368; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3370 = 14'h44 == field_data_lo_366 ? _field_data_T_1062 : _GEN_3369; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3371 = 14'h45 == field_data_lo_366 ? _field_data_T_1063 : _GEN_3370; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_67 = vliw_67[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_387 = vliw_67[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_67 = field_data_lo_387[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_67 = field_data_lo_387[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_148 = {{1'd0}, args_offset_67}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_148 = _total_offset_T_148[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3375 = 3'h1 == total_offset_148 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3376 = 3'h2 == total_offset_148 ? args_2 : _GEN_3375; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3377 = 3'h3 == total_offset_148 ? args_3 : _GEN_3376; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3378 = 3'h4 == total_offset_148 ? args_4 : _GEN_3377; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3379 = 3'h5 == total_offset_148 ? args_5 : _GEN_3378; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3380 = 3'h6 == total_offset_148 ? args_6 : _GEN_3379; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3381 = total_offset_148 < 3'h7 ? _GEN_3380 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_3 = 3'h0 < args_length_67 ? _GEN_3381 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_149 = args_offset_67 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3384 = 3'h1 == total_offset_149 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3385 = 3'h2 == total_offset_149 ? args_2 : _GEN_3384; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3386 = 3'h3 == total_offset_149 ? args_3 : _GEN_3385; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3387 = 3'h4 == total_offset_149 ? args_4 : _GEN_3386; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3388 = 3'h5 == total_offset_149 ? args_5 : _GEN_3387; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3389 = 3'h6 == total_offset_149 ? args_6 : _GEN_3388; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3390 = total_offset_149 < 3'h7 ? _GEN_3389 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_2 = 3'h1 < args_length_67 ? _GEN_3390 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_150 = args_offset_67 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3393 = 3'h1 == total_offset_150 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3394 = 3'h2 == total_offset_150 ? args_2 : _GEN_3393; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3395 = 3'h3 == total_offset_150 ? args_3 : _GEN_3394; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3396 = 3'h4 == total_offset_150 ? args_4 : _GEN_3395; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3397 = 3'h5 == total_offset_150 ? args_5 : _GEN_3396; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3398 = 3'h6 == total_offset_150 ? args_6 : _GEN_3397; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3399 = total_offset_150 < 3'h7 ? _GEN_3398 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_1 = 3'h2 < args_length_67 ? _GEN_3399 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_151 = args_offset_67 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3402 = 3'h1 == total_offset_151 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3403 = 3'h2 == total_offset_151 ? args_2 : _GEN_3402; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3404 = 3'h3 == total_offset_151 ? args_3 : _GEN_3403; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3405 = 3'h4 == total_offset_151 ? args_4 : _GEN_3404; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3406 = 3'h5 == total_offset_151 ? args_5 : _GEN_3405; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3407 = 3'h6 == total_offset_151 ? args_6 : _GEN_3406; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3408 = total_offset_151 < 3'h7 ? _GEN_3407 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_67_0 = 3'h3 < args_length_67 ? _GEN_3408 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1448 = {field_bytes_67_0,field_bytes_67_1,field_bytes_67_2,field_bytes_67_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3410 = opcode_67 == 4'ha ? _field_data_T_1448 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3411 = opcode_67 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2280 = opcode_67 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_423 = field_data_lo_387[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1451 = {field_data_hi_423,field_data_lo_387}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_135 = _T_2280 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3412 = opcode_67 == 4'h8 | opcode_67 == 4'hb ? _field_data_T_1451 : _GEN_3410; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3413 = opcode_67 == 4'h8 | opcode_67 == 4'hb ? _field_tag_T_135 : _GEN_3411; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3414 = 14'h32 == field_data_lo_387 ? _field_data_T_1044 : _GEN_3412; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3415 = 14'h33 == field_data_lo_387 ? _field_data_T_1045 : _GEN_3414; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3416 = 14'h34 == field_data_lo_387 ? _field_data_T_1046 : _GEN_3415; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3417 = 14'h35 == field_data_lo_387 ? _field_data_T_1047 : _GEN_3416; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3418 = 14'h36 == field_data_lo_387 ? _field_data_T_1048 : _GEN_3417; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3419 = 14'h37 == field_data_lo_387 ? _field_data_T_1049 : _GEN_3418; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3420 = 14'h38 == field_data_lo_387 ? _field_data_T_1050 : _GEN_3419; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3421 = 14'h39 == field_data_lo_387 ? _field_data_T_1051 : _GEN_3420; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3422 = 14'h3a == field_data_lo_387 ? _field_data_T_1052 : _GEN_3421; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3423 = 14'h3b == field_data_lo_387 ? _field_data_T_1053 : _GEN_3422; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3424 = 14'h3c == field_data_lo_387 ? _field_data_T_1054 : _GEN_3423; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3425 = 14'h3d == field_data_lo_387 ? _field_data_T_1055 : _GEN_3424; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3426 = 14'h3e == field_data_lo_387 ? _field_data_T_1056 : _GEN_3425; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3427 = 14'h3f == field_data_lo_387 ? _field_data_T_1057 : _GEN_3426; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3428 = 14'h40 == field_data_lo_387 ? _field_data_T_1058 : _GEN_3427; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3429 = 14'h41 == field_data_lo_387 ? _field_data_T_1059 : _GEN_3428; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3430 = 14'h42 == field_data_lo_387 ? _field_data_T_1060 : _GEN_3429; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3431 = 14'h43 == field_data_lo_387 ? _field_data_T_1061 : _GEN_3430; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3432 = 14'h44 == field_data_lo_387 ? _field_data_T_1062 : _GEN_3431; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3433 = 14'h45 == field_data_lo_387 ? _field_data_T_1063 : _GEN_3432; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_68 = vliw_68[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_408 = vliw_68[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_68 = field_data_lo_408[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_68 = field_data_lo_408[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_152 = {{1'd0}, args_offset_68}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_152 = _total_offset_T_152[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3437 = 3'h1 == total_offset_152 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3438 = 3'h2 == total_offset_152 ? args_2 : _GEN_3437; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3439 = 3'h3 == total_offset_152 ? args_3 : _GEN_3438; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3440 = 3'h4 == total_offset_152 ? args_4 : _GEN_3439; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3441 = 3'h5 == total_offset_152 ? args_5 : _GEN_3440; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3442 = 3'h6 == total_offset_152 ? args_6 : _GEN_3441; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3443 = total_offset_152 < 3'h7 ? _GEN_3442 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_3 = 3'h0 < args_length_68 ? _GEN_3443 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_153 = args_offset_68 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3446 = 3'h1 == total_offset_153 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3447 = 3'h2 == total_offset_153 ? args_2 : _GEN_3446; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3448 = 3'h3 == total_offset_153 ? args_3 : _GEN_3447; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3449 = 3'h4 == total_offset_153 ? args_4 : _GEN_3448; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3450 = 3'h5 == total_offset_153 ? args_5 : _GEN_3449; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3451 = 3'h6 == total_offset_153 ? args_6 : _GEN_3450; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3452 = total_offset_153 < 3'h7 ? _GEN_3451 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_2 = 3'h1 < args_length_68 ? _GEN_3452 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_154 = args_offset_68 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3455 = 3'h1 == total_offset_154 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3456 = 3'h2 == total_offset_154 ? args_2 : _GEN_3455; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3457 = 3'h3 == total_offset_154 ? args_3 : _GEN_3456; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3458 = 3'h4 == total_offset_154 ? args_4 : _GEN_3457; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3459 = 3'h5 == total_offset_154 ? args_5 : _GEN_3458; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3460 = 3'h6 == total_offset_154 ? args_6 : _GEN_3459; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3461 = total_offset_154 < 3'h7 ? _GEN_3460 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_1 = 3'h2 < args_length_68 ? _GEN_3461 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_155 = args_offset_68 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3464 = 3'h1 == total_offset_155 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3465 = 3'h2 == total_offset_155 ? args_2 : _GEN_3464; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3466 = 3'h3 == total_offset_155 ? args_3 : _GEN_3465; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3467 = 3'h4 == total_offset_155 ? args_4 : _GEN_3466; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3468 = 3'h5 == total_offset_155 ? args_5 : _GEN_3467; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3469 = 3'h6 == total_offset_155 ? args_6 : _GEN_3468; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3470 = total_offset_155 < 3'h7 ? _GEN_3469 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_68_0 = 3'h3 < args_length_68 ? _GEN_3470 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1472 = {field_bytes_68_0,field_bytes_68_1,field_bytes_68_2,field_bytes_68_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3472 = opcode_68 == 4'ha ? _field_data_T_1472 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3473 = opcode_68 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2313 = opcode_68 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_446 = field_data_lo_408[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1475 = {field_data_hi_446,field_data_lo_408}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_137 = _T_2313 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3474 = opcode_68 == 4'h8 | opcode_68 == 4'hb ? _field_data_T_1475 : _GEN_3472; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3475 = opcode_68 == 4'h8 | opcode_68 == 4'hb ? _field_tag_T_137 : _GEN_3473; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3476 = 14'h32 == field_data_lo_408 ? _field_data_T_1044 : _GEN_3474; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3477 = 14'h33 == field_data_lo_408 ? _field_data_T_1045 : _GEN_3476; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3478 = 14'h34 == field_data_lo_408 ? _field_data_T_1046 : _GEN_3477; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3479 = 14'h35 == field_data_lo_408 ? _field_data_T_1047 : _GEN_3478; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3480 = 14'h36 == field_data_lo_408 ? _field_data_T_1048 : _GEN_3479; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3481 = 14'h37 == field_data_lo_408 ? _field_data_T_1049 : _GEN_3480; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3482 = 14'h38 == field_data_lo_408 ? _field_data_T_1050 : _GEN_3481; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3483 = 14'h39 == field_data_lo_408 ? _field_data_T_1051 : _GEN_3482; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3484 = 14'h3a == field_data_lo_408 ? _field_data_T_1052 : _GEN_3483; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3485 = 14'h3b == field_data_lo_408 ? _field_data_T_1053 : _GEN_3484; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3486 = 14'h3c == field_data_lo_408 ? _field_data_T_1054 : _GEN_3485; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3487 = 14'h3d == field_data_lo_408 ? _field_data_T_1055 : _GEN_3486; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3488 = 14'h3e == field_data_lo_408 ? _field_data_T_1056 : _GEN_3487; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3489 = 14'h3f == field_data_lo_408 ? _field_data_T_1057 : _GEN_3488; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3490 = 14'h40 == field_data_lo_408 ? _field_data_T_1058 : _GEN_3489; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3491 = 14'h41 == field_data_lo_408 ? _field_data_T_1059 : _GEN_3490; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3492 = 14'h42 == field_data_lo_408 ? _field_data_T_1060 : _GEN_3491; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3493 = 14'h43 == field_data_lo_408 ? _field_data_T_1061 : _GEN_3492; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3494 = 14'h44 == field_data_lo_408 ? _field_data_T_1062 : _GEN_3493; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3495 = 14'h45 == field_data_lo_408 ? _field_data_T_1063 : _GEN_3494; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [3:0] opcode_69 = vliw_69[17:14]; // @[executor_pisa.scala 182:38]
  wire [13:0] field_data_lo_429 = vliw_69[13:0]; // @[executor_pisa.scala 183:38]
  wire [2:0] args_offset_69 = field_data_lo_429[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_69 = field_data_lo_429[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _total_offset_T_156 = {{1'd0}, args_offset_69}; // @[executor_pisa.scala 194:49]
  wire [2:0] total_offset_156 = _total_offset_T_156[2:0]; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3499 = 3'h1 == total_offset_156 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3500 = 3'h2 == total_offset_156 ? args_2 : _GEN_3499; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3501 = 3'h3 == total_offset_156 ? args_3 : _GEN_3500; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3502 = 3'h4 == total_offset_156 ? args_4 : _GEN_3501; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3503 = 3'h5 == total_offset_156 ? args_5 : _GEN_3502; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3504 = 3'h6 == total_offset_156 ? args_6 : _GEN_3503; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3505 = total_offset_156 < 3'h7 ? _GEN_3504 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_3 = 3'h0 < args_length_69 ? _GEN_3505 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_157 = args_offset_69 + 3'h1; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3508 = 3'h1 == total_offset_157 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3509 = 3'h2 == total_offset_157 ? args_2 : _GEN_3508; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3510 = 3'h3 == total_offset_157 ? args_3 : _GEN_3509; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3511 = 3'h4 == total_offset_157 ? args_4 : _GEN_3510; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3512 = 3'h5 == total_offset_157 ? args_5 : _GEN_3511; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3513 = 3'h6 == total_offset_157 ? args_6 : _GEN_3512; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3514 = total_offset_157 < 3'h7 ? _GEN_3513 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_2 = 3'h1 < args_length_69 ? _GEN_3514 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_158 = args_offset_69 + 3'h2; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3517 = 3'h1 == total_offset_158 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3518 = 3'h2 == total_offset_158 ? args_2 : _GEN_3517; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3519 = 3'h3 == total_offset_158 ? args_3 : _GEN_3518; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3520 = 3'h4 == total_offset_158 ? args_4 : _GEN_3519; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3521 = 3'h5 == total_offset_158 ? args_5 : _GEN_3520; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3522 = 3'h6 == total_offset_158 ? args_6 : _GEN_3521; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3523 = total_offset_158 < 3'h7 ? _GEN_3522 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_1 = 3'h2 < args_length_69 ? _GEN_3523 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [2:0] total_offset_159 = args_offset_69 + 3'h3; // @[executor_pisa.scala 194:49]
  wire [7:0] _GEN_3526 = 3'h1 == total_offset_159 ? args_1 : args_0; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3527 = 3'h2 == total_offset_159 ? args_2 : _GEN_3526; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3528 = 3'h3 == total_offset_159 ? args_3 : _GEN_3527; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3529 = 3'h4 == total_offset_159 ? args_4 : _GEN_3528; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3530 = 3'h5 == total_offset_159 ? args_5 : _GEN_3529; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3531 = 3'h6 == total_offset_159 ? args_6 : _GEN_3530; // @[executor_pisa.scala 196:59 executor_pisa.scala 196:59]
  wire [7:0] _GEN_3532 = total_offset_159 < 3'h7 ? _GEN_3531 : 8'h0; // @[executor_pisa.scala 195:72 executor_pisa.scala 196:59 executor_pisa.scala 191:51]
  wire [7:0] field_bytes_69_0 = 3'h3 < args_length_69 ? _GEN_3532 : 8'h0; // @[executor_pisa.scala 193:55 executor_pisa.scala 191:51]
  wire [31:0] _field_data_T_1496 = {field_bytes_69_0,field_bytes_69_1,field_bytes_69_2,field_bytes_69_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3534 = opcode_69 == 4'ha ? _field_data_T_1496 : 32'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 200:28 executor_pisa.scala 179:24]
  wire [1:0] _GEN_3535 = opcode_69 == 4'ha ? 2'h2 : 2'h0; // @[executor_pisa.scala 185:47 executor_pisa.scala 201:28 executor_pisa.scala 180:24]
  wire  _T_2346 = opcode_69 == 4'h8; // @[executor_pisa.scala 203:26]
  wire [17:0] field_data_hi_469 = field_data_lo_429[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _field_data_T_1499 = {field_data_hi_469,field_data_lo_429}; // @[Cat.scala 30:58]
  wire [1:0] _field_tag_T_139 = _T_2346 ? 2'h1 : 2'h2; // @[executor_pisa.scala 210:35]
  wire [31:0] _GEN_3536 = opcode_69 == 4'h8 | opcode_69 == 4'hb ? _field_data_T_1499 : _GEN_3534; // @[executor_pisa.scala 203:79 executor_pisa.scala 208:32]
  wire [1:0] _GEN_3537 = opcode_69 == 4'h8 | opcode_69 == 4'hb ? _field_tag_T_139 : _GEN_3535; // @[executor_pisa.scala 203:79 executor_pisa.scala 210:29]
  wire [31:0] _GEN_3538 = 14'h32 == field_data_lo_429 ? _field_data_T_1044 : _GEN_3536; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3539 = 14'h33 == field_data_lo_429 ? _field_data_T_1045 : _GEN_3538; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3540 = 14'h34 == field_data_lo_429 ? _field_data_T_1046 : _GEN_3539; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3541 = 14'h35 == field_data_lo_429 ? _field_data_T_1047 : _GEN_3540; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3542 = 14'h36 == field_data_lo_429 ? _field_data_T_1048 : _GEN_3541; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3543 = 14'h37 == field_data_lo_429 ? _field_data_T_1049 : _GEN_3542; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3544 = 14'h38 == field_data_lo_429 ? _field_data_T_1050 : _GEN_3543; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3545 = 14'h39 == field_data_lo_429 ? _field_data_T_1051 : _GEN_3544; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3546 = 14'h3a == field_data_lo_429 ? _field_data_T_1052 : _GEN_3545; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3547 = 14'h3b == field_data_lo_429 ? _field_data_T_1053 : _GEN_3546; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3548 = 14'h3c == field_data_lo_429 ? _field_data_T_1054 : _GEN_3547; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3549 = 14'h3d == field_data_lo_429 ? _field_data_T_1055 : _GEN_3548; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3550 = 14'h3e == field_data_lo_429 ? _field_data_T_1056 : _GEN_3549; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3551 = 14'h3f == field_data_lo_429 ? _field_data_T_1057 : _GEN_3550; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3552 = 14'h40 == field_data_lo_429 ? _field_data_T_1058 : _GEN_3551; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3553 = 14'h41 == field_data_lo_429 ? _field_data_T_1059 : _GEN_3552; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3554 = 14'h42 == field_data_lo_429 ? _field_data_T_1060 : _GEN_3553; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3555 = 14'h43 == field_data_lo_429 ? _field_data_T_1061 : _GEN_3554; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3556 = 14'h44 == field_data_lo_429 ? _field_data_T_1062 : _GEN_3555; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  wire [31:0] _GEN_3557 = 14'h45 == field_data_lo_429 ? _field_data_T_1063 : _GEN_3556; // @[executor_pisa.scala 216:52 executor_pisa.scala 217:40]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor_pisa.scala 163:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[executor_pisa.scala 163:25]
  assign io_nid_out = nid; // @[executor_pisa.scala 173:20]
  assign io_tag_out_0 = opcode == 4'h9 ? 2'h2 : _GEN_12; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_1 = opcode_1 == 4'h9 ? 2'h2 : _GEN_47; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_2 = opcode_2 == 4'h9 ? 2'h2 : _GEN_82; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_3 = opcode_3 == 4'h9 ? 2'h2 : _GEN_117; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_4 = opcode_4 == 4'h9 ? 2'h2 : _GEN_152; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_5 = opcode_5 == 4'h9 ? 2'h2 : _GEN_187; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_6 = opcode_6 == 4'h9 ? 2'h2 : _GEN_222; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_7 = opcode_7 == 4'h9 ? 2'h2 : _GEN_257; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_8 = opcode_8 == 4'h9 ? 2'h2 : _GEN_292; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_9 = opcode_9 == 4'h9 ? 2'h2 : _GEN_327; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_10 = opcode_10 == 4'h9 ? 2'h2 : _GEN_362; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_11 = opcode_11 == 4'h9 ? 2'h2 : _GEN_397; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_12 = opcode_12 == 4'h9 ? 2'h2 : _GEN_432; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_13 = opcode_13 == 4'h9 ? 2'h2 : _GEN_467; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_14 = opcode_14 == 4'h9 ? 2'h2 : _GEN_502; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_15 = opcode_15 == 4'h9 ? 2'h2 : _GEN_537; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_16 = opcode_16 == 4'h9 ? 2'h2 : _GEN_572; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_17 = opcode_17 == 4'h9 ? 2'h2 : _GEN_607; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_18 = opcode_18 == 4'h9 ? 2'h2 : _GEN_642; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_19 = opcode_19 == 4'h9 ? 2'h2 : _GEN_677; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_20 = opcode_20 == 4'h9 ? 2'h2 : _GEN_721; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_21 = opcode_21 == 4'h9 ? 2'h2 : _GEN_775; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_22 = opcode_22 == 4'h9 ? 2'h2 : _GEN_829; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_23 = opcode_23 == 4'h9 ? 2'h2 : _GEN_883; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_24 = opcode_24 == 4'h9 ? 2'h2 : _GEN_937; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_25 = opcode_25 == 4'h9 ? 2'h2 : _GEN_991; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_26 = opcode_26 == 4'h9 ? 2'h2 : _GEN_1045; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_27 = opcode_27 == 4'h9 ? 2'h2 : _GEN_1099; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_28 = opcode_28 == 4'h9 ? 2'h2 : _GEN_1153; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_29 = opcode_29 == 4'h9 ? 2'h2 : _GEN_1207; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_30 = opcode_30 == 4'h9 ? 2'h2 : _GEN_1261; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_31 = opcode_31 == 4'h9 ? 2'h2 : _GEN_1315; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_32 = opcode_32 == 4'h9 ? 2'h2 : _GEN_1369; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_33 = opcode_33 == 4'h9 ? 2'h2 : _GEN_1423; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_34 = opcode_34 == 4'h9 ? 2'h2 : _GEN_1477; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_35 = opcode_35 == 4'h9 ? 2'h2 : _GEN_1531; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_36 = opcode_36 == 4'h9 ? 2'h2 : _GEN_1585; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_37 = opcode_37 == 4'h9 ? 2'h2 : _GEN_1639; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_38 = opcode_38 == 4'h9 ? 2'h2 : _GEN_1693; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_39 = opcode_39 == 4'h9 ? 2'h2 : _GEN_1747; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_40 = opcode_40 == 4'h9 ? 2'h2 : _GEN_1801; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_41 = opcode_41 == 4'h9 ? 2'h2 : _GEN_1855; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_42 = opcode_42 == 4'h9 ? 2'h2 : _GEN_1909; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_43 = opcode_43 == 4'h9 ? 2'h2 : _GEN_1963; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_44 = opcode_44 == 4'h9 ? 2'h2 : _GEN_2017; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_45 = opcode_45 == 4'h9 ? 2'h2 : _GEN_2071; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_46 = opcode_46 == 4'h9 ? 2'h2 : _GEN_2125; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_47 = opcode_47 == 4'h9 ? 2'h2 : _GEN_2179; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_48 = opcode_48 == 4'h9 ? 2'h2 : _GEN_2233; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_49 = opcode_49 == 4'h9 ? 2'h2 : _GEN_2287; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_50 = opcode_50 == 4'h9 ? 2'h2 : _GEN_2359; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_51 = opcode_51 == 4'h9 ? 2'h2 : _GEN_2421; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_52 = opcode_52 == 4'h9 ? 2'h2 : _GEN_2483; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_53 = opcode_53 == 4'h9 ? 2'h2 : _GEN_2545; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_54 = opcode_54 == 4'h9 ? 2'h2 : _GEN_2607; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_55 = opcode_55 == 4'h9 ? 2'h2 : _GEN_2669; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_56 = opcode_56 == 4'h9 ? 2'h2 : _GEN_2731; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_57 = opcode_57 == 4'h9 ? 2'h2 : _GEN_2793; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_58 = opcode_58 == 4'h9 ? 2'h2 : _GEN_2855; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_59 = opcode_59 == 4'h9 ? 2'h2 : _GEN_2917; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_60 = opcode_60 == 4'h9 ? 2'h2 : _GEN_2979; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_61 = opcode_61 == 4'h9 ? 2'h2 : _GEN_3041; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_62 = opcode_62 == 4'h9 ? 2'h2 : _GEN_3103; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_63 = opcode_63 == 4'h9 ? 2'h2 : _GEN_3165; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_64 = opcode_64 == 4'h9 ? 2'h2 : _GEN_3227; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_65 = opcode_65 == 4'h9 ? 2'h2 : _GEN_3289; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_66 = opcode_66 == 4'h9 ? 2'h2 : _GEN_3351; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_67 = opcode_67 == 4'h9 ? 2'h2 : _GEN_3413; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_68 = opcode_68 == 4'h9 ? 2'h2 : _GEN_3475; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_tag_out_69 = opcode_69 == 4'h9 ? 2'h2 : _GEN_3537; // @[executor_pisa.scala 212:48 executor_pisa.scala 221:29]
  assign io_field_set_field8_0 = opcode == 4'h9 ? _GEN_32 : _GEN_11; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_1 = opcode_1 == 4'h9 ? _GEN_67 : _GEN_46; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_2 = opcode_2 == 4'h9 ? _GEN_102 : _GEN_81; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_3 = opcode_3 == 4'h9 ? _GEN_137 : _GEN_116; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_4 = opcode_4 == 4'h9 ? _GEN_172 : _GEN_151; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_5 = opcode_5 == 4'h9 ? _GEN_207 : _GEN_186; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_6 = opcode_6 == 4'h9 ? _GEN_242 : _GEN_221; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_7 = opcode_7 == 4'h9 ? _GEN_277 : _GEN_256; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_8 = opcode_8 == 4'h9 ? _GEN_312 : _GEN_291; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_9 = opcode_9 == 4'h9 ? _GEN_347 : _GEN_326; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_10 = opcode_10 == 4'h9 ? _GEN_382 : _GEN_361; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_11 = opcode_11 == 4'h9 ? _GEN_417 : _GEN_396; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_12 = opcode_12 == 4'h9 ? _GEN_452 : _GEN_431; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_13 = opcode_13 == 4'h9 ? _GEN_487 : _GEN_466; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_14 = opcode_14 == 4'h9 ? _GEN_522 : _GEN_501; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_15 = opcode_15 == 4'h9 ? _GEN_557 : _GEN_536; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_16 = opcode_16 == 4'h9 ? _GEN_592 : _GEN_571; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_17 = opcode_17 == 4'h9 ? _GEN_627 : _GEN_606; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_18 = opcode_18 == 4'h9 ? _GEN_662 : _GEN_641; // @[executor_pisa.scala 212:48]
  assign io_field_set_field8_19 = opcode_19 == 4'h9 ? _GEN_697 : _GEN_676; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_0 = opcode_20 == 4'h9 ? _GEN_751 : _GEN_720; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_1 = opcode_21 == 4'h9 ? _GEN_805 : _GEN_774; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_2 = opcode_22 == 4'h9 ? _GEN_859 : _GEN_828; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_3 = opcode_23 == 4'h9 ? _GEN_913 : _GEN_882; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_4 = opcode_24 == 4'h9 ? _GEN_967 : _GEN_936; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_5 = opcode_25 == 4'h9 ? _GEN_1021 : _GEN_990; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_6 = opcode_26 == 4'h9 ? _GEN_1075 : _GEN_1044; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_7 = opcode_27 == 4'h9 ? _GEN_1129 : _GEN_1098; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_8 = opcode_28 == 4'h9 ? _GEN_1183 : _GEN_1152; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_9 = opcode_29 == 4'h9 ? _GEN_1237 : _GEN_1206; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_10 = opcode_30 == 4'h9 ? _GEN_1291 : _GEN_1260; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_11 = opcode_31 == 4'h9 ? _GEN_1345 : _GEN_1314; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_12 = opcode_32 == 4'h9 ? _GEN_1399 : _GEN_1368; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_13 = opcode_33 == 4'h9 ? _GEN_1453 : _GEN_1422; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_14 = opcode_34 == 4'h9 ? _GEN_1507 : _GEN_1476; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_15 = opcode_35 == 4'h9 ? _GEN_1561 : _GEN_1530; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_16 = opcode_36 == 4'h9 ? _GEN_1615 : _GEN_1584; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_17 = opcode_37 == 4'h9 ? _GEN_1669 : _GEN_1638; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_18 = opcode_38 == 4'h9 ? _GEN_1723 : _GEN_1692; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_19 = opcode_39 == 4'h9 ? _GEN_1777 : _GEN_1746; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_20 = opcode_40 == 4'h9 ? _GEN_1831 : _GEN_1800; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_21 = opcode_41 == 4'h9 ? _GEN_1885 : _GEN_1854; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_22 = opcode_42 == 4'h9 ? _GEN_1939 : _GEN_1908; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_23 = opcode_43 == 4'h9 ? _GEN_1993 : _GEN_1962; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_24 = opcode_44 == 4'h9 ? _GEN_2047 : _GEN_2016; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_25 = opcode_45 == 4'h9 ? _GEN_2101 : _GEN_2070; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_26 = opcode_46 == 4'h9 ? _GEN_2155 : _GEN_2124; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_27 = opcode_47 == 4'h9 ? _GEN_2209 : _GEN_2178; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_28 = opcode_48 == 4'h9 ? _GEN_2263 : _GEN_2232; // @[executor_pisa.scala 212:48]
  assign io_field_set_field16_29 = opcode_49 == 4'h9 ? _GEN_2317 : _GEN_2286; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_0 = opcode_50 == 4'h9 ? _GEN_2379 : _GEN_2358; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_1 = opcode_51 == 4'h9 ? _GEN_2441 : _GEN_2420; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_2 = opcode_52 == 4'h9 ? _GEN_2503 : _GEN_2482; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_3 = opcode_53 == 4'h9 ? _GEN_2565 : _GEN_2544; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_4 = opcode_54 == 4'h9 ? _GEN_2627 : _GEN_2606; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_5 = opcode_55 == 4'h9 ? _GEN_2689 : _GEN_2668; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_6 = opcode_56 == 4'h9 ? _GEN_2751 : _GEN_2730; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_7 = opcode_57 == 4'h9 ? _GEN_2813 : _GEN_2792; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_8 = opcode_58 == 4'h9 ? _GEN_2875 : _GEN_2854; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_9 = opcode_59 == 4'h9 ? _GEN_2937 : _GEN_2916; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_10 = opcode_60 == 4'h9 ? _GEN_2999 : _GEN_2978; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_11 = opcode_61 == 4'h9 ? _GEN_3061 : _GEN_3040; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_12 = opcode_62 == 4'h9 ? _GEN_3123 : _GEN_3102; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_13 = opcode_63 == 4'h9 ? _GEN_3185 : _GEN_3164; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_14 = opcode_64 == 4'h9 ? _GEN_3247 : _GEN_3226; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_15 = opcode_65 == 4'h9 ? _GEN_3309 : _GEN_3288; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_16 = opcode_66 == 4'h9 ? _GEN_3371 : _GEN_3350; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_17 = opcode_67 == 4'h9 ? _GEN_3433 : _GEN_3412; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_18 = opcode_68 == 4'h9 ? _GEN_3495 : _GEN_3474; // @[executor_pisa.scala 212:48]
  assign io_field_set_field32_19 = opcode_69 == 4'h9 ? _GEN_3557 : _GEN_3536; // @[executor_pisa.scala 212:48]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor_pisa.scala 162:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor_pisa.scala 162:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor_pisa.scala 162:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor_pisa.scala 162:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor_pisa.scala 162:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor_pisa.scala 162:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor_pisa.scala 162:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor_pisa.scala 162:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor_pisa.scala 162:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor_pisa.scala 162:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor_pisa.scala 162:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor_pisa.scala 162:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor_pisa.scala 162:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor_pisa.scala 162:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor_pisa.scala 162:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor_pisa.scala 162:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor_pisa.scala 162:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor_pisa.scala 162:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor_pisa.scala 162:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor_pisa.scala 162:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor_pisa.scala 162:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor_pisa.scala 162:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor_pisa.scala 162:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor_pisa.scala 162:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor_pisa.scala 162:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor_pisa.scala 162:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor_pisa.scala 162:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor_pisa.scala 162:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor_pisa.scala 162:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor_pisa.scala 162:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor_pisa.scala 162:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor_pisa.scala 162:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor_pisa.scala 162:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor_pisa.scala 162:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor_pisa.scala 162:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor_pisa.scala 162:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor_pisa.scala 162:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor_pisa.scala 162:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor_pisa.scala 162:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor_pisa.scala 162:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor_pisa.scala 162:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor_pisa.scala 162:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor_pisa.scala 162:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor_pisa.scala 162:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor_pisa.scala 162:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor_pisa.scala 162:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor_pisa.scala 162:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor_pisa.scala 162:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor_pisa.scala 162:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor_pisa.scala 162:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor_pisa.scala 162:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor_pisa.scala 162:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor_pisa.scala 162:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor_pisa.scala 162:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor_pisa.scala 162:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor_pisa.scala 162:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor_pisa.scala 162:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor_pisa.scala 162:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor_pisa.scala 162:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor_pisa.scala 162:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor_pisa.scala 162:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor_pisa.scala 162:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor_pisa.scala 162:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor_pisa.scala 162:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor_pisa.scala 162:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor_pisa.scala 162:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor_pisa.scala 162:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor_pisa.scala 162:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor_pisa.scala 162:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor_pisa.scala 162:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor_pisa.scala 162:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor_pisa.scala 162:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor_pisa.scala 162:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor_pisa.scala 162:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor_pisa.scala 162:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor_pisa.scala 162:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor_pisa.scala 162:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor_pisa.scala 162:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor_pisa.scala 162:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor_pisa.scala 162:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor_pisa.scala 162:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor_pisa.scala 162:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor_pisa.scala 162:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor_pisa.scala 162:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor_pisa.scala 162:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor_pisa.scala 162:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor_pisa.scala 162:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor_pisa.scala 162:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor_pisa.scala 162:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor_pisa.scala 162:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor_pisa.scala 162:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor_pisa.scala 162:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor_pisa.scala 162:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor_pisa.scala 162:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor_pisa.scala 162:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor_pisa.scala 162:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor_pisa.scala 162:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor_pisa.scala 162:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor_pisa.scala 162:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor_pisa.scala 162:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor_pisa.scala 162:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor_pisa.scala 162:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor_pisa.scala 162:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor_pisa.scala 162:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor_pisa.scala 162:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor_pisa.scala 162:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor_pisa.scala 162:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor_pisa.scala 162:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor_pisa.scala 162:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor_pisa.scala 162:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor_pisa.scala 162:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor_pisa.scala 162:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor_pisa.scala 162:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor_pisa.scala 162:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor_pisa.scala 162:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor_pisa.scala 162:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor_pisa.scala 162:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor_pisa.scala 162:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor_pisa.scala 162:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor_pisa.scala 162:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor_pisa.scala 162:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor_pisa.scala 162:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor_pisa.scala 162:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor_pisa.scala 162:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor_pisa.scala 162:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor_pisa.scala 162:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor_pisa.scala 162:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor_pisa.scala 162:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor_pisa.scala 162:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor_pisa.scala 162:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor_pisa.scala 162:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor_pisa.scala 162:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor_pisa.scala 162:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor_pisa.scala 162:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor_pisa.scala 162:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor_pisa.scala 162:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor_pisa.scala 162:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor_pisa.scala 162:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor_pisa.scala 162:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor_pisa.scala 162:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor_pisa.scala 162:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor_pisa.scala 162:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor_pisa.scala 162:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor_pisa.scala 162:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor_pisa.scala 162:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor_pisa.scala 162:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor_pisa.scala 162:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor_pisa.scala 162:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor_pisa.scala 162:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor_pisa.scala 162:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor_pisa.scala 162:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor_pisa.scala 162:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor_pisa.scala 162:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor_pisa.scala 162:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor_pisa.scala 162:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor_pisa.scala 162:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor_pisa.scala 162:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor_pisa.scala 162:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor_pisa.scala 162:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor_pisa.scala 162:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor_pisa.scala 162:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 162:13]
    args_0 <= io_args_in_0; // @[executor_pisa.scala 166:14]
    args_1 <= io_args_in_1; // @[executor_pisa.scala 166:14]
    args_2 <= io_args_in_2; // @[executor_pisa.scala 166:14]
    args_3 <= io_args_in_3; // @[executor_pisa.scala 166:14]
    args_4 <= io_args_in_4; // @[executor_pisa.scala 166:14]
    args_5 <= io_args_in_5; // @[executor_pisa.scala 166:14]
    args_6 <= io_args_in_6; // @[executor_pisa.scala 166:14]
    vliw_0 <= io_vliw_in_0; // @[executor_pisa.scala 169:14]
    vliw_1 <= io_vliw_in_1; // @[executor_pisa.scala 169:14]
    vliw_2 <= io_vliw_in_2; // @[executor_pisa.scala 169:14]
    vliw_3 <= io_vliw_in_3; // @[executor_pisa.scala 169:14]
    vliw_4 <= io_vliw_in_4; // @[executor_pisa.scala 169:14]
    vliw_5 <= io_vliw_in_5; // @[executor_pisa.scala 169:14]
    vliw_6 <= io_vliw_in_6; // @[executor_pisa.scala 169:14]
    vliw_7 <= io_vliw_in_7; // @[executor_pisa.scala 169:14]
    vliw_8 <= io_vliw_in_8; // @[executor_pisa.scala 169:14]
    vliw_9 <= io_vliw_in_9; // @[executor_pisa.scala 169:14]
    vliw_10 <= io_vliw_in_10; // @[executor_pisa.scala 169:14]
    vliw_11 <= io_vliw_in_11; // @[executor_pisa.scala 169:14]
    vliw_12 <= io_vliw_in_12; // @[executor_pisa.scala 169:14]
    vliw_13 <= io_vliw_in_13; // @[executor_pisa.scala 169:14]
    vliw_14 <= io_vliw_in_14; // @[executor_pisa.scala 169:14]
    vliw_15 <= io_vliw_in_15; // @[executor_pisa.scala 169:14]
    vliw_16 <= io_vliw_in_16; // @[executor_pisa.scala 169:14]
    vliw_17 <= io_vliw_in_17; // @[executor_pisa.scala 169:14]
    vliw_18 <= io_vliw_in_18; // @[executor_pisa.scala 169:14]
    vliw_19 <= io_vliw_in_19; // @[executor_pisa.scala 169:14]
    vliw_20 <= io_vliw_in_20; // @[executor_pisa.scala 169:14]
    vliw_21 <= io_vliw_in_21; // @[executor_pisa.scala 169:14]
    vliw_22 <= io_vliw_in_22; // @[executor_pisa.scala 169:14]
    vliw_23 <= io_vliw_in_23; // @[executor_pisa.scala 169:14]
    vliw_24 <= io_vliw_in_24; // @[executor_pisa.scala 169:14]
    vliw_25 <= io_vliw_in_25; // @[executor_pisa.scala 169:14]
    vliw_26 <= io_vliw_in_26; // @[executor_pisa.scala 169:14]
    vliw_27 <= io_vliw_in_27; // @[executor_pisa.scala 169:14]
    vliw_28 <= io_vliw_in_28; // @[executor_pisa.scala 169:14]
    vliw_29 <= io_vliw_in_29; // @[executor_pisa.scala 169:14]
    vliw_30 <= io_vliw_in_30; // @[executor_pisa.scala 169:14]
    vliw_31 <= io_vliw_in_31; // @[executor_pisa.scala 169:14]
    vliw_32 <= io_vliw_in_32; // @[executor_pisa.scala 169:14]
    vliw_33 <= io_vliw_in_33; // @[executor_pisa.scala 169:14]
    vliw_34 <= io_vliw_in_34; // @[executor_pisa.scala 169:14]
    vliw_35 <= io_vliw_in_35; // @[executor_pisa.scala 169:14]
    vliw_36 <= io_vliw_in_36; // @[executor_pisa.scala 169:14]
    vliw_37 <= io_vliw_in_37; // @[executor_pisa.scala 169:14]
    vliw_38 <= io_vliw_in_38; // @[executor_pisa.scala 169:14]
    vliw_39 <= io_vliw_in_39; // @[executor_pisa.scala 169:14]
    vliw_40 <= io_vliw_in_40; // @[executor_pisa.scala 169:14]
    vliw_41 <= io_vliw_in_41; // @[executor_pisa.scala 169:14]
    vliw_42 <= io_vliw_in_42; // @[executor_pisa.scala 169:14]
    vliw_43 <= io_vliw_in_43; // @[executor_pisa.scala 169:14]
    vliw_44 <= io_vliw_in_44; // @[executor_pisa.scala 169:14]
    vliw_45 <= io_vliw_in_45; // @[executor_pisa.scala 169:14]
    vliw_46 <= io_vliw_in_46; // @[executor_pisa.scala 169:14]
    vliw_47 <= io_vliw_in_47; // @[executor_pisa.scala 169:14]
    vliw_48 <= io_vliw_in_48; // @[executor_pisa.scala 169:14]
    vliw_49 <= io_vliw_in_49; // @[executor_pisa.scala 169:14]
    vliw_50 <= io_vliw_in_50; // @[executor_pisa.scala 169:14]
    vliw_51 <= io_vliw_in_51; // @[executor_pisa.scala 169:14]
    vliw_52 <= io_vliw_in_52; // @[executor_pisa.scala 169:14]
    vliw_53 <= io_vliw_in_53; // @[executor_pisa.scala 169:14]
    vliw_54 <= io_vliw_in_54; // @[executor_pisa.scala 169:14]
    vliw_55 <= io_vliw_in_55; // @[executor_pisa.scala 169:14]
    vliw_56 <= io_vliw_in_56; // @[executor_pisa.scala 169:14]
    vliw_57 <= io_vliw_in_57; // @[executor_pisa.scala 169:14]
    vliw_58 <= io_vliw_in_58; // @[executor_pisa.scala 169:14]
    vliw_59 <= io_vliw_in_59; // @[executor_pisa.scala 169:14]
    vliw_60 <= io_vliw_in_60; // @[executor_pisa.scala 169:14]
    vliw_61 <= io_vliw_in_61; // @[executor_pisa.scala 169:14]
    vliw_62 <= io_vliw_in_62; // @[executor_pisa.scala 169:14]
    vliw_63 <= io_vliw_in_63; // @[executor_pisa.scala 169:14]
    vliw_64 <= io_vliw_in_64; // @[executor_pisa.scala 169:14]
    vliw_65 <= io_vliw_in_65; // @[executor_pisa.scala 169:14]
    vliw_66 <= io_vliw_in_66; // @[executor_pisa.scala 169:14]
    vliw_67 <= io_vliw_in_67; // @[executor_pisa.scala 169:14]
    vliw_68 <= io_vliw_in_68; // @[executor_pisa.scala 169:14]
    vliw_69 <= io_vliw_in_69; // @[executor_pisa.scala 169:14]
    nid <= io_nid_in; // @[executor_pisa.scala 172:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  phv_next_config_id = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  args_0 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  args_1 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  args_2 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  args_3 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  args_4 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  args_5 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  args_6 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  vliw_0 = _RAND_169[17:0];
  _RAND_170 = {1{`RANDOM}};
  vliw_1 = _RAND_170[17:0];
  _RAND_171 = {1{`RANDOM}};
  vliw_2 = _RAND_171[17:0];
  _RAND_172 = {1{`RANDOM}};
  vliw_3 = _RAND_172[17:0];
  _RAND_173 = {1{`RANDOM}};
  vliw_4 = _RAND_173[17:0];
  _RAND_174 = {1{`RANDOM}};
  vliw_5 = _RAND_174[17:0];
  _RAND_175 = {1{`RANDOM}};
  vliw_6 = _RAND_175[17:0];
  _RAND_176 = {1{`RANDOM}};
  vliw_7 = _RAND_176[17:0];
  _RAND_177 = {1{`RANDOM}};
  vliw_8 = _RAND_177[17:0];
  _RAND_178 = {1{`RANDOM}};
  vliw_9 = _RAND_178[17:0];
  _RAND_179 = {1{`RANDOM}};
  vliw_10 = _RAND_179[17:0];
  _RAND_180 = {1{`RANDOM}};
  vliw_11 = _RAND_180[17:0];
  _RAND_181 = {1{`RANDOM}};
  vliw_12 = _RAND_181[17:0];
  _RAND_182 = {1{`RANDOM}};
  vliw_13 = _RAND_182[17:0];
  _RAND_183 = {1{`RANDOM}};
  vliw_14 = _RAND_183[17:0];
  _RAND_184 = {1{`RANDOM}};
  vliw_15 = _RAND_184[17:0];
  _RAND_185 = {1{`RANDOM}};
  vliw_16 = _RAND_185[17:0];
  _RAND_186 = {1{`RANDOM}};
  vliw_17 = _RAND_186[17:0];
  _RAND_187 = {1{`RANDOM}};
  vliw_18 = _RAND_187[17:0];
  _RAND_188 = {1{`RANDOM}};
  vliw_19 = _RAND_188[17:0];
  _RAND_189 = {1{`RANDOM}};
  vliw_20 = _RAND_189[17:0];
  _RAND_190 = {1{`RANDOM}};
  vliw_21 = _RAND_190[17:0];
  _RAND_191 = {1{`RANDOM}};
  vliw_22 = _RAND_191[17:0];
  _RAND_192 = {1{`RANDOM}};
  vliw_23 = _RAND_192[17:0];
  _RAND_193 = {1{`RANDOM}};
  vliw_24 = _RAND_193[17:0];
  _RAND_194 = {1{`RANDOM}};
  vliw_25 = _RAND_194[17:0];
  _RAND_195 = {1{`RANDOM}};
  vliw_26 = _RAND_195[17:0];
  _RAND_196 = {1{`RANDOM}};
  vliw_27 = _RAND_196[17:0];
  _RAND_197 = {1{`RANDOM}};
  vliw_28 = _RAND_197[17:0];
  _RAND_198 = {1{`RANDOM}};
  vliw_29 = _RAND_198[17:0];
  _RAND_199 = {1{`RANDOM}};
  vliw_30 = _RAND_199[17:0];
  _RAND_200 = {1{`RANDOM}};
  vliw_31 = _RAND_200[17:0];
  _RAND_201 = {1{`RANDOM}};
  vliw_32 = _RAND_201[17:0];
  _RAND_202 = {1{`RANDOM}};
  vliw_33 = _RAND_202[17:0];
  _RAND_203 = {1{`RANDOM}};
  vliw_34 = _RAND_203[17:0];
  _RAND_204 = {1{`RANDOM}};
  vliw_35 = _RAND_204[17:0];
  _RAND_205 = {1{`RANDOM}};
  vliw_36 = _RAND_205[17:0];
  _RAND_206 = {1{`RANDOM}};
  vliw_37 = _RAND_206[17:0];
  _RAND_207 = {1{`RANDOM}};
  vliw_38 = _RAND_207[17:0];
  _RAND_208 = {1{`RANDOM}};
  vliw_39 = _RAND_208[17:0];
  _RAND_209 = {1{`RANDOM}};
  vliw_40 = _RAND_209[17:0];
  _RAND_210 = {1{`RANDOM}};
  vliw_41 = _RAND_210[17:0];
  _RAND_211 = {1{`RANDOM}};
  vliw_42 = _RAND_211[17:0];
  _RAND_212 = {1{`RANDOM}};
  vliw_43 = _RAND_212[17:0];
  _RAND_213 = {1{`RANDOM}};
  vliw_44 = _RAND_213[17:0];
  _RAND_214 = {1{`RANDOM}};
  vliw_45 = _RAND_214[17:0];
  _RAND_215 = {1{`RANDOM}};
  vliw_46 = _RAND_215[17:0];
  _RAND_216 = {1{`RANDOM}};
  vliw_47 = _RAND_216[17:0];
  _RAND_217 = {1{`RANDOM}};
  vliw_48 = _RAND_217[17:0];
  _RAND_218 = {1{`RANDOM}};
  vliw_49 = _RAND_218[17:0];
  _RAND_219 = {1{`RANDOM}};
  vliw_50 = _RAND_219[17:0];
  _RAND_220 = {1{`RANDOM}};
  vliw_51 = _RAND_220[17:0];
  _RAND_221 = {1{`RANDOM}};
  vliw_52 = _RAND_221[17:0];
  _RAND_222 = {1{`RANDOM}};
  vliw_53 = _RAND_222[17:0];
  _RAND_223 = {1{`RANDOM}};
  vliw_54 = _RAND_223[17:0];
  _RAND_224 = {1{`RANDOM}};
  vliw_55 = _RAND_224[17:0];
  _RAND_225 = {1{`RANDOM}};
  vliw_56 = _RAND_225[17:0];
  _RAND_226 = {1{`RANDOM}};
  vliw_57 = _RAND_226[17:0];
  _RAND_227 = {1{`RANDOM}};
  vliw_58 = _RAND_227[17:0];
  _RAND_228 = {1{`RANDOM}};
  vliw_59 = _RAND_228[17:0];
  _RAND_229 = {1{`RANDOM}};
  vliw_60 = _RAND_229[17:0];
  _RAND_230 = {1{`RANDOM}};
  vliw_61 = _RAND_230[17:0];
  _RAND_231 = {1{`RANDOM}};
  vliw_62 = _RAND_231[17:0];
  _RAND_232 = {1{`RANDOM}};
  vliw_63 = _RAND_232[17:0];
  _RAND_233 = {1{`RANDOM}};
  vliw_64 = _RAND_233[17:0];
  _RAND_234 = {1{`RANDOM}};
  vliw_65 = _RAND_234[17:0];
  _RAND_235 = {1{`RANDOM}};
  vliw_66 = _RAND_235[17:0];
  _RAND_236 = {1{`RANDOM}};
  vliw_67 = _RAND_236[17:0];
  _RAND_237 = {1{`RANDOM}};
  vliw_68 = _RAND_237[17:0];
  _RAND_238 = {1{`RANDOM}};
  vliw_69 = _RAND_238[17:0];
  _RAND_239 = {1{`RANDOM}};
  nid = _RAND_239[14:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
