module IPSAPCIE(
  input         clock,
  input         reset,
  input         io_pcie_r_en,
  input  [19:0] io_pcie_r_addr,
  output [63:0] io_pcie_r_data,
  input         io_pcie_w_en,
  input  [19:0] io_pcie_w_addr,
  input  [63:0] io_pcie_w_data
);
  wire  ipsa_clock; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_0; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_1; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_2; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_3; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_4; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_5; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_6; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_7; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_8; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_9; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_10; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_11; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_12; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_13; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_14; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_15; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_16; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_17; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_18; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_19; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_20; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_21; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_22; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_23; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_24; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_25; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_26; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_27; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_28; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_29; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_30; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_31; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_32; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_33; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_34; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_35; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_36; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_37; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_38; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_39; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_40; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_41; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_42; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_43; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_44; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_45; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_46; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_47; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_48; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_49; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_50; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_51; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_52; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_53; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_54; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_55; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_56; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_57; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_58; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_59; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_60; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_61; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_62; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_63; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_64; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_65; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_66; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_67; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_68; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_69; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_70; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_71; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_72; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_73; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_74; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_75; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_76; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_77; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_78; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_79; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_80; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_81; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_82; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_83; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_84; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_85; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_86; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_87; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_88; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_89; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_90; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_91; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_92; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_93; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_94; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_95; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_96; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_97; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_98; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_99; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_100; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_101; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_102; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_103; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_104; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_105; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_106; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_107; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_108; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_109; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_110; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_111; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_112; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_113; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_114; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_115; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_116; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_117; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_118; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_119; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_120; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_121; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_122; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_123; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_124; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_125; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_126; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_127; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_128; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_129; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_130; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_131; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_132; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_133; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_134; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_135; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_136; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_137; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_138; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_139; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_140; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_141; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_142; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_143; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_144; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_145; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_146; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_147; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_148; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_149; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_150; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_151; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_152; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_153; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_154; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_155; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_156; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_157; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_158; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_159; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_160; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_161; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_162; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_163; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_164; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_165; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_166; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_167; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_168; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_169; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_170; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_171; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_172; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_173; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_174; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_175; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_176; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_177; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_178; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_179; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_180; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_181; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_182; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_183; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_184; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_185; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_186; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_187; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_188; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_189; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_190; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_in_data_191; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_0; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_1; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_2; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_3; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_4; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_5; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_6; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_7; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_8; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_9; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_10; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_11; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_12; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_13; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_14; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_15; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_16; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_17; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_18; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_19; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_20; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_21; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_22; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_23; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_24; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_25; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_26; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_27; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_28; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_29; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_30; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_31; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_32; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_33; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_34; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_35; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_36; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_37; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_38; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_39; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_40; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_41; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_42; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_43; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_44; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_45; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_46; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_47; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_48; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_49; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_50; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_51; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_52; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_53; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_54; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_55; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_56; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_57; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_58; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_59; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_60; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_61; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_62; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_63; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_64; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_65; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_66; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_67; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_68; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_69; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_70; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_71; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_72; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_73; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_74; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_75; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_76; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_77; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_78; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_79; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_80; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_81; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_82; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_83; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_84; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_85; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_86; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_87; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_88; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_89; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_90; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_91; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_92; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_93; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_94; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_95; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_96; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_97; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_98; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_99; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_100; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_101; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_102; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_103; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_104; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_105; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_106; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_107; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_108; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_109; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_110; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_111; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_112; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_113; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_114; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_115; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_116; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_117; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_118; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_119; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_120; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_121; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_122; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_123; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_124; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_125; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_126; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_127; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_128; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_129; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_130; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_131; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_132; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_133; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_134; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_135; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_136; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_137; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_138; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_139; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_140; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_141; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_142; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_143; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_144; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_145; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_146; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_147; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_148; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_149; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_150; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_151; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_152; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_153; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_154; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_155; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_156; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_157; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_158; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_159; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_160; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_161; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_162; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_163; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_164; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_165; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_166; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_167; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_168; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_169; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_170; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_171; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_172; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_173; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_174; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_175; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_176; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_177; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_178; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_179; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_180; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_181; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_182; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_183; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_184; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_185; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_186; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_187; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_188; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_189; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_190; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_191; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_192; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_193; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_194; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_195; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_196; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_197; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_198; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_199; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_200; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_201; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_202; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_203; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_204; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_205; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_206; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_207; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_208; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_209; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_210; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_211; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_212; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_213; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_214; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_215; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_216; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_217; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_218; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_219; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_220; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_221; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_222; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_223; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_224; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_225; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_226; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_227; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_228; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_229; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_230; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_231; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_232; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_233; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_234; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_235; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_236; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_237; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_238; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_239; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_240; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_241; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_242; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_243; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_244; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_245; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_246; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_247; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_248; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_249; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_250; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_251; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_252; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_253; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_254; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_pipe_phv_out_data_255; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_par_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_0_par_mod_last_mau_id; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_0_par_mod_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_0_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_mat_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_mat_mod_config_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_0_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_0_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_0_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_0_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_act_mod_en_0; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_0_act_mod_en_1; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_0_act_mod_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_0_act_mod_data_0; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_0_act_mod_data_1; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_par_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_1_par_mod_last_mau_id; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_1_par_mod_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_1_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_mat_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_mat_mod_config_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_1_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_1_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_1_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_1_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_act_mod_en_0; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_1_act_mod_en_1; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_1_act_mod_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_1_act_mod_data_0; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_1_act_mod_data_1; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_par_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_2_par_mod_last_mau_id; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_2_par_mod_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_2_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_mat_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_mat_mod_config_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_2_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_2_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_2_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_2_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_act_mod_en_0; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_2_act_mod_en_1; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_2_act_mod_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_2_act_mod_data_0; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_2_act_mod_data_1; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_par_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_3_par_mod_last_mau_id; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_proc_mod_3_par_mod_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_3_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_mat_mod_en; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_mat_mod_config_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_3_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_3_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_3_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 13:22]
  wire [6:0] ipsa_io_mod_proc_mod_3_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_act_mod_en_0; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_proc_mod_3_act_mod_en_1; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_mod_proc_mod_3_act_mod_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_3_act_mod_data_0; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_mod_proc_mod_3_act_mod_data_1; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_mod_xbar_mod_en; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_xbar_mod_first_proc_id; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_xbar_mod_last_proc_id; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_xbar_mod_next_proc_id_0; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_xbar_mod_next_proc_id_1; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_xbar_mod_next_proc_id_2; // @[ipsa_pcie.scala 13:22]
  wire [1:0] ipsa_io_mod_xbar_mod_next_proc_id_3; // @[ipsa_pcie.scala 13:22]
  wire [5:0] ipsa_io_w_0_wcs; // @[ipsa_pcie.scala 13:22]
  wire  ipsa_io_w_0_w_en; // @[ipsa_pcie.scala 13:22]
  wire [7:0] ipsa_io_w_0_w_addr; // @[ipsa_pcie.scala 13:22]
  wire [63:0] ipsa_io_w_0_w_data; // @[ipsa_pcie.scala 13:22]
  wire  pcie_clock; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_pcie_r_en; // @[ipsa_pcie.scala 14:22]
  wire [19:0] pcie_io_pcie_r_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_pcie_r_data; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_pcie_w_en; // @[ipsa_pcie.scala 14:22]
  wire [19:0] pcie_io_pcie_w_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_pcie_w_data; // @[ipsa_pcie.scala 14:22]
  wire [4:0] pcie_io_pcie_o_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_pcie_o_r_en; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_pcie_o_r_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_pcie_o_r_data; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_par_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_0_par_mod_last_mau_id; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_0_par_mod_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_0_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_mat_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_mat_mod_config_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_0_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_0_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_0_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_0_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_act_mod_en_0; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_0_act_mod_en_1; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_0_act_mod_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_0_act_mod_data_0; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_0_act_mod_data_1; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_par_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_1_par_mod_last_mau_id; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_1_par_mod_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_1_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_mat_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_mat_mod_config_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_1_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_1_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_1_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_1_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_act_mod_en_0; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_1_act_mod_en_1; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_1_act_mod_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_1_act_mod_data_0; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_1_act_mod_data_1; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_par_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_2_par_mod_last_mau_id; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_2_par_mod_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_2_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_mat_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_mat_mod_config_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_2_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_2_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_2_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_2_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_act_mod_en_0; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_2_act_mod_en_1; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_2_act_mod_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_2_act_mod_data_0; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_2_act_mod_data_1; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_par_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_3_par_mod_last_mau_id; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_proc_mod_3_par_mod_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_par_mod_module_mod_state_id_mod; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_3_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_mat_mod_en; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_mat_mod_config_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_3_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_3_mat_mod_key_mod_internal_offset; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_3_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 14:22]
  wire [6:0] pcie_io_mod_proc_mod_3_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_act_mod_en_0; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_proc_mod_3_act_mod_en_1; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_mod_proc_mod_3_act_mod_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_3_act_mod_data_0; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_mod_proc_mod_3_act_mod_data_1; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_mod_xbar_mod_en; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_xbar_mod_first_proc_id; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_xbar_mod_last_proc_id; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_xbar_mod_next_proc_id_0; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_xbar_mod_next_proc_id_1; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_xbar_mod_next_proc_id_2; // @[ipsa_pcie.scala 14:22]
  wire [1:0] pcie_io_mod_xbar_mod_next_proc_id_3; // @[ipsa_pcie.scala 14:22]
  wire [5:0] pcie_io_w_0_wcs; // @[ipsa_pcie.scala 14:22]
  wire  pcie_io_w_0_w_en; // @[ipsa_pcie.scala 14:22]
  wire [7:0] pcie_io_w_0_w_addr; // @[ipsa_pcie.scala 14:22]
  wire [63:0] pcie_io_w_0_w_data; // @[ipsa_pcie.scala 14:22]
  wire  outp_clock; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_0; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_1; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_2; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_3; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_4; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_5; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_6; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_7; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_8; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_9; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_10; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_11; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_12; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_13; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_14; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_15; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_16; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_17; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_18; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_19; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_20; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_21; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_22; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_23; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_24; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_25; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_26; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_27; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_28; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_29; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_30; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_31; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_32; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_33; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_34; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_35; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_36; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_37; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_38; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_39; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_40; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_41; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_42; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_43; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_44; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_45; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_46; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_47; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_48; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_49; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_50; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_51; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_52; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_53; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_54; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_55; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_56; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_57; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_58; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_59; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_60; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_61; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_62; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_63; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_64; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_65; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_66; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_67; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_68; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_69; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_70; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_71; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_72; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_73; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_74; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_75; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_76; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_77; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_78; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_79; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_80; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_81; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_82; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_83; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_84; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_85; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_86; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_87; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_88; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_89; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_90; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_91; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_92; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_93; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_94; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_95; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_96; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_97; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_98; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_99; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_100; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_101; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_102; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_103; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_104; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_105; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_106; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_107; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_108; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_109; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_110; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_111; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_112; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_113; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_114; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_115; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_116; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_117; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_118; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_119; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_120; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_121; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_122; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_123; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_124; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_125; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_126; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_127; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_128; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_129; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_130; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_131; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_132; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_133; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_134; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_135; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_136; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_137; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_138; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_139; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_140; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_141; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_142; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_143; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_144; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_145; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_146; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_147; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_148; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_149; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_150; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_151; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_152; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_153; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_154; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_155; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_156; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_157; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_158; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_159; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_160; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_161; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_162; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_163; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_164; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_165; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_166; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_167; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_168; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_169; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_170; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_171; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_172; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_173; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_174; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_175; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_176; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_177; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_178; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_179; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_180; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_181; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_182; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_183; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_184; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_185; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_186; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_187; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_188; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_189; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_190; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_191; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_192; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_193; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_194; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_195; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_196; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_197; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_198; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_199; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_200; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_201; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_202; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_203; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_204; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_205; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_206; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_207; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_208; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_209; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_210; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_211; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_212; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_213; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_214; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_215; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_216; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_217; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_218; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_219; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_220; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_221; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_222; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_223; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_224; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_225; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_226; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_227; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_228; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_229; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_230; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_231; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_232; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_233; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_234; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_235; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_236; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_237; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_238; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_239; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_240; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_241; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_242; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_243; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_244; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_245; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_246; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_247; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_248; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_249; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_250; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_251; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_252; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_253; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_254; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_phv_in_data_255; // @[ipsa_pcie.scala 15:22]
  wire [4:0] outp_io_pcie_o_cs; // @[ipsa_pcie.scala 15:22]
  wire  outp_io_pcie_o_r_en; // @[ipsa_pcie.scala 15:22]
  wire [7:0] outp_io_pcie_o_r_addr; // @[ipsa_pcie.scala 15:22]
  wire [63:0] outp_io_pcie_o_r_data; // @[ipsa_pcie.scala 15:22]
  wire  inp_clock; // @[ipsa_pcie.scala 16:22]
  wire  inp_reset; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_0; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_1; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_2; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_3; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_4; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_5; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_6; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_7; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_8; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_9; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_10; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_11; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_12; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_13; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_14; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_15; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_16; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_17; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_18; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_19; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_20; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_21; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_22; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_23; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_24; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_25; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_26; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_27; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_28; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_29; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_30; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_31; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_32; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_33; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_34; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_35; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_36; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_37; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_38; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_39; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_40; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_41; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_42; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_43; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_44; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_45; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_46; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_47; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_48; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_49; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_50; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_51; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_52; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_53; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_54; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_55; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_56; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_57; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_58; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_59; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_60; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_61; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_62; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_63; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_64; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_65; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_66; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_67; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_68; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_69; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_70; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_71; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_72; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_73; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_74; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_75; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_76; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_77; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_78; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_79; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_80; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_81; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_82; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_83; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_84; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_85; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_86; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_87; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_88; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_89; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_90; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_91; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_92; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_93; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_94; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_95; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_96; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_97; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_98; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_99; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_100; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_101; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_102; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_103; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_104; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_105; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_106; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_107; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_108; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_109; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_110; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_111; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_112; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_113; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_114; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_115; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_116; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_117; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_118; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_119; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_120; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_121; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_122; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_123; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_124; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_125; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_126; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_127; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_128; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_129; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_130; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_131; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_132; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_133; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_134; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_135; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_136; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_137; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_138; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_139; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_140; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_141; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_142; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_143; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_144; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_145; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_146; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_147; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_148; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_149; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_150; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_151; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_152; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_153; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_154; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_155; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_156; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_157; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_158; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_159; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_160; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_161; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_162; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_163; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_164; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_165; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_166; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_167; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_168; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_169; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_170; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_171; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_172; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_173; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_174; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_175; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_176; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_177; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_178; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_179; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_180; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_181; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_182; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_183; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_184; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_185; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_186; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_187; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_188; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_189; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_190; // @[ipsa_pcie.scala 16:22]
  wire [7:0] inp_io_phv_out_data_191; // @[ipsa_pcie.scala 16:22]
  IPSA ipsa ( // @[ipsa_pcie.scala 13:22]
    .clock(ipsa_clock),
    .io_pipe_phv_in_data_0(ipsa_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(ipsa_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(ipsa_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(ipsa_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(ipsa_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(ipsa_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(ipsa_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(ipsa_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(ipsa_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(ipsa_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(ipsa_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(ipsa_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(ipsa_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(ipsa_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(ipsa_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(ipsa_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(ipsa_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(ipsa_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(ipsa_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(ipsa_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(ipsa_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(ipsa_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(ipsa_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(ipsa_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(ipsa_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(ipsa_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(ipsa_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(ipsa_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(ipsa_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(ipsa_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(ipsa_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(ipsa_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(ipsa_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(ipsa_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(ipsa_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(ipsa_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(ipsa_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(ipsa_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(ipsa_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(ipsa_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(ipsa_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(ipsa_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(ipsa_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(ipsa_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(ipsa_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(ipsa_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(ipsa_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(ipsa_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(ipsa_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(ipsa_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(ipsa_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(ipsa_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(ipsa_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(ipsa_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(ipsa_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(ipsa_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(ipsa_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(ipsa_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(ipsa_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(ipsa_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(ipsa_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(ipsa_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(ipsa_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(ipsa_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(ipsa_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(ipsa_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(ipsa_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(ipsa_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(ipsa_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(ipsa_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(ipsa_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(ipsa_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(ipsa_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(ipsa_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(ipsa_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(ipsa_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(ipsa_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(ipsa_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(ipsa_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(ipsa_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(ipsa_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(ipsa_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(ipsa_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(ipsa_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(ipsa_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(ipsa_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(ipsa_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(ipsa_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(ipsa_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(ipsa_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(ipsa_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(ipsa_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(ipsa_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(ipsa_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(ipsa_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(ipsa_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(ipsa_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(ipsa_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(ipsa_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(ipsa_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(ipsa_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(ipsa_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(ipsa_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(ipsa_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(ipsa_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(ipsa_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(ipsa_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(ipsa_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(ipsa_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(ipsa_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(ipsa_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(ipsa_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(ipsa_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(ipsa_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(ipsa_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(ipsa_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(ipsa_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(ipsa_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(ipsa_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(ipsa_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(ipsa_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(ipsa_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(ipsa_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(ipsa_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(ipsa_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(ipsa_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(ipsa_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(ipsa_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(ipsa_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(ipsa_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(ipsa_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(ipsa_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(ipsa_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(ipsa_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(ipsa_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(ipsa_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(ipsa_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(ipsa_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(ipsa_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(ipsa_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(ipsa_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(ipsa_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(ipsa_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(ipsa_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(ipsa_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(ipsa_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(ipsa_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(ipsa_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(ipsa_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(ipsa_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(ipsa_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(ipsa_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(ipsa_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(ipsa_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(ipsa_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(ipsa_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(ipsa_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(ipsa_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(ipsa_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(ipsa_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(ipsa_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(ipsa_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(ipsa_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(ipsa_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(ipsa_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(ipsa_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(ipsa_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(ipsa_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(ipsa_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(ipsa_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(ipsa_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(ipsa_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(ipsa_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(ipsa_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(ipsa_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(ipsa_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(ipsa_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(ipsa_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(ipsa_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(ipsa_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(ipsa_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(ipsa_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(ipsa_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(ipsa_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(ipsa_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(ipsa_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(ipsa_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(ipsa_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(ipsa_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(ipsa_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(ipsa_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(ipsa_io_pipe_phv_in_data_191),
    .io_pipe_phv_out_data_0(ipsa_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(ipsa_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(ipsa_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(ipsa_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(ipsa_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(ipsa_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(ipsa_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(ipsa_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(ipsa_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(ipsa_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(ipsa_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(ipsa_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(ipsa_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(ipsa_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(ipsa_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(ipsa_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(ipsa_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(ipsa_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(ipsa_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(ipsa_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(ipsa_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(ipsa_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(ipsa_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(ipsa_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(ipsa_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(ipsa_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(ipsa_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(ipsa_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(ipsa_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(ipsa_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(ipsa_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(ipsa_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(ipsa_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(ipsa_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(ipsa_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(ipsa_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(ipsa_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(ipsa_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(ipsa_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(ipsa_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(ipsa_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(ipsa_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(ipsa_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(ipsa_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(ipsa_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(ipsa_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(ipsa_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(ipsa_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(ipsa_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(ipsa_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(ipsa_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(ipsa_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(ipsa_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(ipsa_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(ipsa_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(ipsa_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(ipsa_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(ipsa_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(ipsa_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(ipsa_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(ipsa_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(ipsa_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(ipsa_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(ipsa_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(ipsa_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(ipsa_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(ipsa_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(ipsa_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(ipsa_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(ipsa_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(ipsa_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(ipsa_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(ipsa_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(ipsa_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(ipsa_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(ipsa_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(ipsa_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(ipsa_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(ipsa_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(ipsa_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(ipsa_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(ipsa_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(ipsa_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(ipsa_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(ipsa_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(ipsa_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(ipsa_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(ipsa_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(ipsa_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(ipsa_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(ipsa_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(ipsa_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(ipsa_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(ipsa_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(ipsa_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(ipsa_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(ipsa_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(ipsa_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(ipsa_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(ipsa_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(ipsa_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(ipsa_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(ipsa_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(ipsa_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(ipsa_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(ipsa_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(ipsa_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(ipsa_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(ipsa_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(ipsa_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(ipsa_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(ipsa_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(ipsa_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(ipsa_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(ipsa_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(ipsa_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(ipsa_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(ipsa_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(ipsa_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(ipsa_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(ipsa_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(ipsa_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(ipsa_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(ipsa_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(ipsa_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(ipsa_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(ipsa_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(ipsa_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(ipsa_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(ipsa_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(ipsa_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(ipsa_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(ipsa_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(ipsa_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(ipsa_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(ipsa_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(ipsa_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(ipsa_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(ipsa_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(ipsa_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(ipsa_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(ipsa_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(ipsa_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(ipsa_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(ipsa_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(ipsa_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(ipsa_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(ipsa_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(ipsa_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(ipsa_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(ipsa_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(ipsa_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(ipsa_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(ipsa_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(ipsa_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(ipsa_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(ipsa_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(ipsa_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(ipsa_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(ipsa_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(ipsa_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(ipsa_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(ipsa_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(ipsa_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(ipsa_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(ipsa_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(ipsa_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(ipsa_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(ipsa_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(ipsa_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(ipsa_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(ipsa_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(ipsa_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(ipsa_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(ipsa_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(ipsa_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(ipsa_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(ipsa_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(ipsa_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(ipsa_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(ipsa_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(ipsa_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(ipsa_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(ipsa_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(ipsa_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(ipsa_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(ipsa_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(ipsa_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(ipsa_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(ipsa_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(ipsa_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(ipsa_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(ipsa_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(ipsa_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(ipsa_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(ipsa_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(ipsa_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(ipsa_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(ipsa_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(ipsa_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(ipsa_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(ipsa_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(ipsa_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(ipsa_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(ipsa_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(ipsa_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(ipsa_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(ipsa_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(ipsa_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(ipsa_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(ipsa_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(ipsa_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(ipsa_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(ipsa_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(ipsa_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(ipsa_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(ipsa_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(ipsa_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(ipsa_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(ipsa_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(ipsa_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(ipsa_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(ipsa_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(ipsa_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(ipsa_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(ipsa_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(ipsa_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(ipsa_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(ipsa_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(ipsa_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(ipsa_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(ipsa_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(ipsa_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(ipsa_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(ipsa_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(ipsa_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(ipsa_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(ipsa_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(ipsa_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(ipsa_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(ipsa_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(ipsa_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(ipsa_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(ipsa_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(ipsa_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(ipsa_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(ipsa_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(ipsa_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(ipsa_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(ipsa_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(ipsa_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(ipsa_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(ipsa_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(ipsa_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(ipsa_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(ipsa_io_pipe_phv_out_data_255),
    .io_mod_proc_mod_0_par_mod_en(ipsa_io_mod_proc_mod_0_par_mod_en),
    .io_mod_proc_mod_0_par_mod_last_mau_id_mod(ipsa_io_mod_proc_mod_0_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_0_par_mod_last_mau_id(ipsa_io_mod_proc_mod_0_par_mod_last_mau_id),
    .io_mod_proc_mod_0_par_mod_cs(ipsa_io_mod_proc_mod_0_par_mod_cs),
    .io_mod_proc_mod_0_par_mod_module_mod_state_id_mod(ipsa_io_mod_proc_mod_0_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_0_par_mod_module_mod_state_id(ipsa_io_mod_proc_mod_0_par_mod_module_mod_state_id),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs(ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_en(ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr(ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_data(ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_0_mat_mod_en(ipsa_io_mod_proc_mod_0_mat_mod_en),
    .io_mod_proc_mod_0_mat_mod_config_id(ipsa_io_mod_proc_mod_0_mat_mod_config_id),
    .io_mod_proc_mod_0_mat_mod_key_mod_header_id(ipsa_io_mod_proc_mod_0_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_0_mat_mod_key_mod_internal_offset(ipsa_io_mod_proc_mod_0_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_0_mat_mod_key_mod_key_length(ipsa_io_mod_proc_mod_0_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_0_mat_mod_table_mod_table_width(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_0_mat_mod_table_mod_table_depth(ipsa_io_mod_proc_mod_0_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_0_act_mod_en_0(ipsa_io_mod_proc_mod_0_act_mod_en_0),
    .io_mod_proc_mod_0_act_mod_en_1(ipsa_io_mod_proc_mod_0_act_mod_en_1),
    .io_mod_proc_mod_0_act_mod_addr(ipsa_io_mod_proc_mod_0_act_mod_addr),
    .io_mod_proc_mod_0_act_mod_data_0(ipsa_io_mod_proc_mod_0_act_mod_data_0),
    .io_mod_proc_mod_0_act_mod_data_1(ipsa_io_mod_proc_mod_0_act_mod_data_1),
    .io_mod_proc_mod_1_par_mod_en(ipsa_io_mod_proc_mod_1_par_mod_en),
    .io_mod_proc_mod_1_par_mod_last_mau_id_mod(ipsa_io_mod_proc_mod_1_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_1_par_mod_last_mau_id(ipsa_io_mod_proc_mod_1_par_mod_last_mau_id),
    .io_mod_proc_mod_1_par_mod_cs(ipsa_io_mod_proc_mod_1_par_mod_cs),
    .io_mod_proc_mod_1_par_mod_module_mod_state_id_mod(ipsa_io_mod_proc_mod_1_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_1_par_mod_module_mod_state_id(ipsa_io_mod_proc_mod_1_par_mod_module_mod_state_id),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs(ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_en(ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr(ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_data(ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_1_mat_mod_en(ipsa_io_mod_proc_mod_1_mat_mod_en),
    .io_mod_proc_mod_1_mat_mod_config_id(ipsa_io_mod_proc_mod_1_mat_mod_config_id),
    .io_mod_proc_mod_1_mat_mod_key_mod_header_id(ipsa_io_mod_proc_mod_1_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_1_mat_mod_key_mod_internal_offset(ipsa_io_mod_proc_mod_1_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_1_mat_mod_key_mod_key_length(ipsa_io_mod_proc_mod_1_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_1_mat_mod_table_mod_table_width(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_1_mat_mod_table_mod_table_depth(ipsa_io_mod_proc_mod_1_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_1_act_mod_en_0(ipsa_io_mod_proc_mod_1_act_mod_en_0),
    .io_mod_proc_mod_1_act_mod_en_1(ipsa_io_mod_proc_mod_1_act_mod_en_1),
    .io_mod_proc_mod_1_act_mod_addr(ipsa_io_mod_proc_mod_1_act_mod_addr),
    .io_mod_proc_mod_1_act_mod_data_0(ipsa_io_mod_proc_mod_1_act_mod_data_0),
    .io_mod_proc_mod_1_act_mod_data_1(ipsa_io_mod_proc_mod_1_act_mod_data_1),
    .io_mod_proc_mod_2_par_mod_en(ipsa_io_mod_proc_mod_2_par_mod_en),
    .io_mod_proc_mod_2_par_mod_last_mau_id_mod(ipsa_io_mod_proc_mod_2_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_2_par_mod_last_mau_id(ipsa_io_mod_proc_mod_2_par_mod_last_mau_id),
    .io_mod_proc_mod_2_par_mod_cs(ipsa_io_mod_proc_mod_2_par_mod_cs),
    .io_mod_proc_mod_2_par_mod_module_mod_state_id_mod(ipsa_io_mod_proc_mod_2_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_2_par_mod_module_mod_state_id(ipsa_io_mod_proc_mod_2_par_mod_module_mod_state_id),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs(ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_en(ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr(ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_data(ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_2_mat_mod_en(ipsa_io_mod_proc_mod_2_mat_mod_en),
    .io_mod_proc_mod_2_mat_mod_config_id(ipsa_io_mod_proc_mod_2_mat_mod_config_id),
    .io_mod_proc_mod_2_mat_mod_key_mod_header_id(ipsa_io_mod_proc_mod_2_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_2_mat_mod_key_mod_internal_offset(ipsa_io_mod_proc_mod_2_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_2_mat_mod_key_mod_key_length(ipsa_io_mod_proc_mod_2_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_2_mat_mod_table_mod_table_width(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_2_mat_mod_table_mod_table_depth(ipsa_io_mod_proc_mod_2_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_2_act_mod_en_0(ipsa_io_mod_proc_mod_2_act_mod_en_0),
    .io_mod_proc_mod_2_act_mod_en_1(ipsa_io_mod_proc_mod_2_act_mod_en_1),
    .io_mod_proc_mod_2_act_mod_addr(ipsa_io_mod_proc_mod_2_act_mod_addr),
    .io_mod_proc_mod_2_act_mod_data_0(ipsa_io_mod_proc_mod_2_act_mod_data_0),
    .io_mod_proc_mod_2_act_mod_data_1(ipsa_io_mod_proc_mod_2_act_mod_data_1),
    .io_mod_proc_mod_3_par_mod_en(ipsa_io_mod_proc_mod_3_par_mod_en),
    .io_mod_proc_mod_3_par_mod_last_mau_id_mod(ipsa_io_mod_proc_mod_3_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_3_par_mod_last_mau_id(ipsa_io_mod_proc_mod_3_par_mod_last_mau_id),
    .io_mod_proc_mod_3_par_mod_cs(ipsa_io_mod_proc_mod_3_par_mod_cs),
    .io_mod_proc_mod_3_par_mod_module_mod_state_id_mod(ipsa_io_mod_proc_mod_3_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_3_par_mod_module_mod_state_id(ipsa_io_mod_proc_mod_3_par_mod_module_mod_state_id),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs(ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_en(ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr(ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_data(ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_3_mat_mod_en(ipsa_io_mod_proc_mod_3_mat_mod_en),
    .io_mod_proc_mod_3_mat_mod_config_id(ipsa_io_mod_proc_mod_3_mat_mod_config_id),
    .io_mod_proc_mod_3_mat_mod_key_mod_header_id(ipsa_io_mod_proc_mod_3_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_3_mat_mod_key_mod_internal_offset(ipsa_io_mod_proc_mod_3_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_3_mat_mod_key_mod_key_length(ipsa_io_mod_proc_mod_3_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_3_mat_mod_table_mod_table_width(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_3_mat_mod_table_mod_table_depth(ipsa_io_mod_proc_mod_3_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_3_act_mod_en_0(ipsa_io_mod_proc_mod_3_act_mod_en_0),
    .io_mod_proc_mod_3_act_mod_en_1(ipsa_io_mod_proc_mod_3_act_mod_en_1),
    .io_mod_proc_mod_3_act_mod_addr(ipsa_io_mod_proc_mod_3_act_mod_addr),
    .io_mod_proc_mod_3_act_mod_data_0(ipsa_io_mod_proc_mod_3_act_mod_data_0),
    .io_mod_proc_mod_3_act_mod_data_1(ipsa_io_mod_proc_mod_3_act_mod_data_1),
    .io_mod_xbar_mod_en(ipsa_io_mod_xbar_mod_en),
    .io_mod_xbar_mod_first_proc_id(ipsa_io_mod_xbar_mod_first_proc_id),
    .io_mod_xbar_mod_last_proc_id(ipsa_io_mod_xbar_mod_last_proc_id),
    .io_mod_xbar_mod_next_proc_id_0(ipsa_io_mod_xbar_mod_next_proc_id_0),
    .io_mod_xbar_mod_next_proc_id_1(ipsa_io_mod_xbar_mod_next_proc_id_1),
    .io_mod_xbar_mod_next_proc_id_2(ipsa_io_mod_xbar_mod_next_proc_id_2),
    .io_mod_xbar_mod_next_proc_id_3(ipsa_io_mod_xbar_mod_next_proc_id_3),
    .io_w_0_wcs(ipsa_io_w_0_wcs),
    .io_w_0_w_en(ipsa_io_w_0_w_en),
    .io_w_0_w_addr(ipsa_io_w_0_w_addr),
    .io_w_0_w_data(ipsa_io_w_0_w_data)
  );
  PCIEInterface pcie ( // @[ipsa_pcie.scala 14:22]
    .clock(pcie_clock),
    .io_pcie_r_en(pcie_io_pcie_r_en),
    .io_pcie_r_addr(pcie_io_pcie_r_addr),
    .io_pcie_r_data(pcie_io_pcie_r_data),
    .io_pcie_w_en(pcie_io_pcie_w_en),
    .io_pcie_w_addr(pcie_io_pcie_w_addr),
    .io_pcie_w_data(pcie_io_pcie_w_data),
    .io_pcie_o_cs(pcie_io_pcie_o_cs),
    .io_pcie_o_r_en(pcie_io_pcie_o_r_en),
    .io_pcie_o_r_addr(pcie_io_pcie_o_r_addr),
    .io_pcie_o_r_data(pcie_io_pcie_o_r_data),
    .io_mod_proc_mod_0_par_mod_en(pcie_io_mod_proc_mod_0_par_mod_en),
    .io_mod_proc_mod_0_par_mod_last_mau_id_mod(pcie_io_mod_proc_mod_0_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_0_par_mod_last_mau_id(pcie_io_mod_proc_mod_0_par_mod_last_mau_id),
    .io_mod_proc_mod_0_par_mod_cs(pcie_io_mod_proc_mod_0_par_mod_cs),
    .io_mod_proc_mod_0_par_mod_module_mod_state_id_mod(pcie_io_mod_proc_mod_0_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_0_par_mod_module_mod_state_id(pcie_io_mod_proc_mod_0_par_mod_module_mod_state_id),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs(pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_en(pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr(pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_0_par_mod_module_mod_sram_w_data(pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_0_mat_mod_en(pcie_io_mod_proc_mod_0_mat_mod_en),
    .io_mod_proc_mod_0_mat_mod_config_id(pcie_io_mod_proc_mod_0_mat_mod_config_id),
    .io_mod_proc_mod_0_mat_mod_key_mod_header_id(pcie_io_mod_proc_mod_0_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_0_mat_mod_key_mod_internal_offset(pcie_io_mod_proc_mod_0_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_0_mat_mod_key_mod_key_length(pcie_io_mod_proc_mod_0_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63(pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_0_mat_mod_table_mod_table_width(pcie_io_mod_proc_mod_0_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_0_mat_mod_table_mod_table_depth(pcie_io_mod_proc_mod_0_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_0_act_mod_en_0(pcie_io_mod_proc_mod_0_act_mod_en_0),
    .io_mod_proc_mod_0_act_mod_en_1(pcie_io_mod_proc_mod_0_act_mod_en_1),
    .io_mod_proc_mod_0_act_mod_addr(pcie_io_mod_proc_mod_0_act_mod_addr),
    .io_mod_proc_mod_0_act_mod_data_0(pcie_io_mod_proc_mod_0_act_mod_data_0),
    .io_mod_proc_mod_0_act_mod_data_1(pcie_io_mod_proc_mod_0_act_mod_data_1),
    .io_mod_proc_mod_1_par_mod_en(pcie_io_mod_proc_mod_1_par_mod_en),
    .io_mod_proc_mod_1_par_mod_last_mau_id_mod(pcie_io_mod_proc_mod_1_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_1_par_mod_last_mau_id(pcie_io_mod_proc_mod_1_par_mod_last_mau_id),
    .io_mod_proc_mod_1_par_mod_cs(pcie_io_mod_proc_mod_1_par_mod_cs),
    .io_mod_proc_mod_1_par_mod_module_mod_state_id_mod(pcie_io_mod_proc_mod_1_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_1_par_mod_module_mod_state_id(pcie_io_mod_proc_mod_1_par_mod_module_mod_state_id),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs(pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_en(pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr(pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_1_par_mod_module_mod_sram_w_data(pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_1_mat_mod_en(pcie_io_mod_proc_mod_1_mat_mod_en),
    .io_mod_proc_mod_1_mat_mod_config_id(pcie_io_mod_proc_mod_1_mat_mod_config_id),
    .io_mod_proc_mod_1_mat_mod_key_mod_header_id(pcie_io_mod_proc_mod_1_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_1_mat_mod_key_mod_internal_offset(pcie_io_mod_proc_mod_1_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_1_mat_mod_key_mod_key_length(pcie_io_mod_proc_mod_1_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63(pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_1_mat_mod_table_mod_table_width(pcie_io_mod_proc_mod_1_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_1_mat_mod_table_mod_table_depth(pcie_io_mod_proc_mod_1_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_1_act_mod_en_0(pcie_io_mod_proc_mod_1_act_mod_en_0),
    .io_mod_proc_mod_1_act_mod_en_1(pcie_io_mod_proc_mod_1_act_mod_en_1),
    .io_mod_proc_mod_1_act_mod_addr(pcie_io_mod_proc_mod_1_act_mod_addr),
    .io_mod_proc_mod_1_act_mod_data_0(pcie_io_mod_proc_mod_1_act_mod_data_0),
    .io_mod_proc_mod_1_act_mod_data_1(pcie_io_mod_proc_mod_1_act_mod_data_1),
    .io_mod_proc_mod_2_par_mod_en(pcie_io_mod_proc_mod_2_par_mod_en),
    .io_mod_proc_mod_2_par_mod_last_mau_id_mod(pcie_io_mod_proc_mod_2_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_2_par_mod_last_mau_id(pcie_io_mod_proc_mod_2_par_mod_last_mau_id),
    .io_mod_proc_mod_2_par_mod_cs(pcie_io_mod_proc_mod_2_par_mod_cs),
    .io_mod_proc_mod_2_par_mod_module_mod_state_id_mod(pcie_io_mod_proc_mod_2_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_2_par_mod_module_mod_state_id(pcie_io_mod_proc_mod_2_par_mod_module_mod_state_id),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs(pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_en(pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr(pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_2_par_mod_module_mod_sram_w_data(pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_2_mat_mod_en(pcie_io_mod_proc_mod_2_mat_mod_en),
    .io_mod_proc_mod_2_mat_mod_config_id(pcie_io_mod_proc_mod_2_mat_mod_config_id),
    .io_mod_proc_mod_2_mat_mod_key_mod_header_id(pcie_io_mod_proc_mod_2_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_2_mat_mod_key_mod_internal_offset(pcie_io_mod_proc_mod_2_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_2_mat_mod_key_mod_key_length(pcie_io_mod_proc_mod_2_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63(pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_2_mat_mod_table_mod_table_width(pcie_io_mod_proc_mod_2_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_2_mat_mod_table_mod_table_depth(pcie_io_mod_proc_mod_2_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_2_act_mod_en_0(pcie_io_mod_proc_mod_2_act_mod_en_0),
    .io_mod_proc_mod_2_act_mod_en_1(pcie_io_mod_proc_mod_2_act_mod_en_1),
    .io_mod_proc_mod_2_act_mod_addr(pcie_io_mod_proc_mod_2_act_mod_addr),
    .io_mod_proc_mod_2_act_mod_data_0(pcie_io_mod_proc_mod_2_act_mod_data_0),
    .io_mod_proc_mod_2_act_mod_data_1(pcie_io_mod_proc_mod_2_act_mod_data_1),
    .io_mod_proc_mod_3_par_mod_en(pcie_io_mod_proc_mod_3_par_mod_en),
    .io_mod_proc_mod_3_par_mod_last_mau_id_mod(pcie_io_mod_proc_mod_3_par_mod_last_mau_id_mod),
    .io_mod_proc_mod_3_par_mod_last_mau_id(pcie_io_mod_proc_mod_3_par_mod_last_mau_id),
    .io_mod_proc_mod_3_par_mod_cs(pcie_io_mod_proc_mod_3_par_mod_cs),
    .io_mod_proc_mod_3_par_mod_module_mod_state_id_mod(pcie_io_mod_proc_mod_3_par_mod_module_mod_state_id_mod),
    .io_mod_proc_mod_3_par_mod_module_mod_state_id(pcie_io_mod_proc_mod_3_par_mod_module_mod_state_id),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs(pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_en(pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_en),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr(pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr),
    .io_mod_proc_mod_3_par_mod_module_mod_sram_w_data(pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_data),
    .io_mod_proc_mod_3_mat_mod_en(pcie_io_mod_proc_mod_3_mat_mod_en),
    .io_mod_proc_mod_3_mat_mod_config_id(pcie_io_mod_proc_mod_3_mat_mod_config_id),
    .io_mod_proc_mod_3_mat_mod_key_mod_header_id(pcie_io_mod_proc_mod_3_mat_mod_key_mod_header_id),
    .io_mod_proc_mod_3_mat_mod_key_mod_internal_offset(pcie_io_mod_proc_mod_3_mat_mod_key_mod_internal_offset),
    .io_mod_proc_mod_3_mat_mod_key_mod_key_length(pcie_io_mod_proc_mod_3_mat_mod_key_mod_key_length),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62),
    .io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63(pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63),
    .io_mod_proc_mod_3_mat_mod_table_mod_table_width(pcie_io_mod_proc_mod_3_mat_mod_table_mod_table_width),
    .io_mod_proc_mod_3_mat_mod_table_mod_table_depth(pcie_io_mod_proc_mod_3_mat_mod_table_mod_table_depth),
    .io_mod_proc_mod_3_act_mod_en_0(pcie_io_mod_proc_mod_3_act_mod_en_0),
    .io_mod_proc_mod_3_act_mod_en_1(pcie_io_mod_proc_mod_3_act_mod_en_1),
    .io_mod_proc_mod_3_act_mod_addr(pcie_io_mod_proc_mod_3_act_mod_addr),
    .io_mod_proc_mod_3_act_mod_data_0(pcie_io_mod_proc_mod_3_act_mod_data_0),
    .io_mod_proc_mod_3_act_mod_data_1(pcie_io_mod_proc_mod_3_act_mod_data_1),
    .io_mod_xbar_mod_en(pcie_io_mod_xbar_mod_en),
    .io_mod_xbar_mod_first_proc_id(pcie_io_mod_xbar_mod_first_proc_id),
    .io_mod_xbar_mod_last_proc_id(pcie_io_mod_xbar_mod_last_proc_id),
    .io_mod_xbar_mod_next_proc_id_0(pcie_io_mod_xbar_mod_next_proc_id_0),
    .io_mod_xbar_mod_next_proc_id_1(pcie_io_mod_xbar_mod_next_proc_id_1),
    .io_mod_xbar_mod_next_proc_id_2(pcie_io_mod_xbar_mod_next_proc_id_2),
    .io_mod_xbar_mod_next_proc_id_3(pcie_io_mod_xbar_mod_next_proc_id_3),
    .io_w_0_wcs(pcie_io_w_0_wcs),
    .io_w_0_w_en(pcie_io_w_0_w_en),
    .io_w_0_w_addr(pcie_io_w_0_w_addr),
    .io_w_0_w_data(pcie_io_w_0_w_data)
  );
  OutPort outp ( // @[ipsa_pcie.scala 15:22]
    .clock(outp_clock),
    .io_phv_in_data_0(outp_io_phv_in_data_0),
    .io_phv_in_data_1(outp_io_phv_in_data_1),
    .io_phv_in_data_2(outp_io_phv_in_data_2),
    .io_phv_in_data_3(outp_io_phv_in_data_3),
    .io_phv_in_data_4(outp_io_phv_in_data_4),
    .io_phv_in_data_5(outp_io_phv_in_data_5),
    .io_phv_in_data_6(outp_io_phv_in_data_6),
    .io_phv_in_data_7(outp_io_phv_in_data_7),
    .io_phv_in_data_8(outp_io_phv_in_data_8),
    .io_phv_in_data_9(outp_io_phv_in_data_9),
    .io_phv_in_data_10(outp_io_phv_in_data_10),
    .io_phv_in_data_11(outp_io_phv_in_data_11),
    .io_phv_in_data_12(outp_io_phv_in_data_12),
    .io_phv_in_data_13(outp_io_phv_in_data_13),
    .io_phv_in_data_14(outp_io_phv_in_data_14),
    .io_phv_in_data_15(outp_io_phv_in_data_15),
    .io_phv_in_data_16(outp_io_phv_in_data_16),
    .io_phv_in_data_17(outp_io_phv_in_data_17),
    .io_phv_in_data_18(outp_io_phv_in_data_18),
    .io_phv_in_data_19(outp_io_phv_in_data_19),
    .io_phv_in_data_20(outp_io_phv_in_data_20),
    .io_phv_in_data_21(outp_io_phv_in_data_21),
    .io_phv_in_data_22(outp_io_phv_in_data_22),
    .io_phv_in_data_23(outp_io_phv_in_data_23),
    .io_phv_in_data_24(outp_io_phv_in_data_24),
    .io_phv_in_data_25(outp_io_phv_in_data_25),
    .io_phv_in_data_26(outp_io_phv_in_data_26),
    .io_phv_in_data_27(outp_io_phv_in_data_27),
    .io_phv_in_data_28(outp_io_phv_in_data_28),
    .io_phv_in_data_29(outp_io_phv_in_data_29),
    .io_phv_in_data_30(outp_io_phv_in_data_30),
    .io_phv_in_data_31(outp_io_phv_in_data_31),
    .io_phv_in_data_32(outp_io_phv_in_data_32),
    .io_phv_in_data_33(outp_io_phv_in_data_33),
    .io_phv_in_data_34(outp_io_phv_in_data_34),
    .io_phv_in_data_35(outp_io_phv_in_data_35),
    .io_phv_in_data_36(outp_io_phv_in_data_36),
    .io_phv_in_data_37(outp_io_phv_in_data_37),
    .io_phv_in_data_38(outp_io_phv_in_data_38),
    .io_phv_in_data_39(outp_io_phv_in_data_39),
    .io_phv_in_data_40(outp_io_phv_in_data_40),
    .io_phv_in_data_41(outp_io_phv_in_data_41),
    .io_phv_in_data_42(outp_io_phv_in_data_42),
    .io_phv_in_data_43(outp_io_phv_in_data_43),
    .io_phv_in_data_44(outp_io_phv_in_data_44),
    .io_phv_in_data_45(outp_io_phv_in_data_45),
    .io_phv_in_data_46(outp_io_phv_in_data_46),
    .io_phv_in_data_47(outp_io_phv_in_data_47),
    .io_phv_in_data_48(outp_io_phv_in_data_48),
    .io_phv_in_data_49(outp_io_phv_in_data_49),
    .io_phv_in_data_50(outp_io_phv_in_data_50),
    .io_phv_in_data_51(outp_io_phv_in_data_51),
    .io_phv_in_data_52(outp_io_phv_in_data_52),
    .io_phv_in_data_53(outp_io_phv_in_data_53),
    .io_phv_in_data_54(outp_io_phv_in_data_54),
    .io_phv_in_data_55(outp_io_phv_in_data_55),
    .io_phv_in_data_56(outp_io_phv_in_data_56),
    .io_phv_in_data_57(outp_io_phv_in_data_57),
    .io_phv_in_data_58(outp_io_phv_in_data_58),
    .io_phv_in_data_59(outp_io_phv_in_data_59),
    .io_phv_in_data_60(outp_io_phv_in_data_60),
    .io_phv_in_data_61(outp_io_phv_in_data_61),
    .io_phv_in_data_62(outp_io_phv_in_data_62),
    .io_phv_in_data_63(outp_io_phv_in_data_63),
    .io_phv_in_data_64(outp_io_phv_in_data_64),
    .io_phv_in_data_65(outp_io_phv_in_data_65),
    .io_phv_in_data_66(outp_io_phv_in_data_66),
    .io_phv_in_data_67(outp_io_phv_in_data_67),
    .io_phv_in_data_68(outp_io_phv_in_data_68),
    .io_phv_in_data_69(outp_io_phv_in_data_69),
    .io_phv_in_data_70(outp_io_phv_in_data_70),
    .io_phv_in_data_71(outp_io_phv_in_data_71),
    .io_phv_in_data_72(outp_io_phv_in_data_72),
    .io_phv_in_data_73(outp_io_phv_in_data_73),
    .io_phv_in_data_74(outp_io_phv_in_data_74),
    .io_phv_in_data_75(outp_io_phv_in_data_75),
    .io_phv_in_data_76(outp_io_phv_in_data_76),
    .io_phv_in_data_77(outp_io_phv_in_data_77),
    .io_phv_in_data_78(outp_io_phv_in_data_78),
    .io_phv_in_data_79(outp_io_phv_in_data_79),
    .io_phv_in_data_80(outp_io_phv_in_data_80),
    .io_phv_in_data_81(outp_io_phv_in_data_81),
    .io_phv_in_data_82(outp_io_phv_in_data_82),
    .io_phv_in_data_83(outp_io_phv_in_data_83),
    .io_phv_in_data_84(outp_io_phv_in_data_84),
    .io_phv_in_data_85(outp_io_phv_in_data_85),
    .io_phv_in_data_86(outp_io_phv_in_data_86),
    .io_phv_in_data_87(outp_io_phv_in_data_87),
    .io_phv_in_data_88(outp_io_phv_in_data_88),
    .io_phv_in_data_89(outp_io_phv_in_data_89),
    .io_phv_in_data_90(outp_io_phv_in_data_90),
    .io_phv_in_data_91(outp_io_phv_in_data_91),
    .io_phv_in_data_92(outp_io_phv_in_data_92),
    .io_phv_in_data_93(outp_io_phv_in_data_93),
    .io_phv_in_data_94(outp_io_phv_in_data_94),
    .io_phv_in_data_95(outp_io_phv_in_data_95),
    .io_phv_in_data_96(outp_io_phv_in_data_96),
    .io_phv_in_data_97(outp_io_phv_in_data_97),
    .io_phv_in_data_98(outp_io_phv_in_data_98),
    .io_phv_in_data_99(outp_io_phv_in_data_99),
    .io_phv_in_data_100(outp_io_phv_in_data_100),
    .io_phv_in_data_101(outp_io_phv_in_data_101),
    .io_phv_in_data_102(outp_io_phv_in_data_102),
    .io_phv_in_data_103(outp_io_phv_in_data_103),
    .io_phv_in_data_104(outp_io_phv_in_data_104),
    .io_phv_in_data_105(outp_io_phv_in_data_105),
    .io_phv_in_data_106(outp_io_phv_in_data_106),
    .io_phv_in_data_107(outp_io_phv_in_data_107),
    .io_phv_in_data_108(outp_io_phv_in_data_108),
    .io_phv_in_data_109(outp_io_phv_in_data_109),
    .io_phv_in_data_110(outp_io_phv_in_data_110),
    .io_phv_in_data_111(outp_io_phv_in_data_111),
    .io_phv_in_data_112(outp_io_phv_in_data_112),
    .io_phv_in_data_113(outp_io_phv_in_data_113),
    .io_phv_in_data_114(outp_io_phv_in_data_114),
    .io_phv_in_data_115(outp_io_phv_in_data_115),
    .io_phv_in_data_116(outp_io_phv_in_data_116),
    .io_phv_in_data_117(outp_io_phv_in_data_117),
    .io_phv_in_data_118(outp_io_phv_in_data_118),
    .io_phv_in_data_119(outp_io_phv_in_data_119),
    .io_phv_in_data_120(outp_io_phv_in_data_120),
    .io_phv_in_data_121(outp_io_phv_in_data_121),
    .io_phv_in_data_122(outp_io_phv_in_data_122),
    .io_phv_in_data_123(outp_io_phv_in_data_123),
    .io_phv_in_data_124(outp_io_phv_in_data_124),
    .io_phv_in_data_125(outp_io_phv_in_data_125),
    .io_phv_in_data_126(outp_io_phv_in_data_126),
    .io_phv_in_data_127(outp_io_phv_in_data_127),
    .io_phv_in_data_128(outp_io_phv_in_data_128),
    .io_phv_in_data_129(outp_io_phv_in_data_129),
    .io_phv_in_data_130(outp_io_phv_in_data_130),
    .io_phv_in_data_131(outp_io_phv_in_data_131),
    .io_phv_in_data_132(outp_io_phv_in_data_132),
    .io_phv_in_data_133(outp_io_phv_in_data_133),
    .io_phv_in_data_134(outp_io_phv_in_data_134),
    .io_phv_in_data_135(outp_io_phv_in_data_135),
    .io_phv_in_data_136(outp_io_phv_in_data_136),
    .io_phv_in_data_137(outp_io_phv_in_data_137),
    .io_phv_in_data_138(outp_io_phv_in_data_138),
    .io_phv_in_data_139(outp_io_phv_in_data_139),
    .io_phv_in_data_140(outp_io_phv_in_data_140),
    .io_phv_in_data_141(outp_io_phv_in_data_141),
    .io_phv_in_data_142(outp_io_phv_in_data_142),
    .io_phv_in_data_143(outp_io_phv_in_data_143),
    .io_phv_in_data_144(outp_io_phv_in_data_144),
    .io_phv_in_data_145(outp_io_phv_in_data_145),
    .io_phv_in_data_146(outp_io_phv_in_data_146),
    .io_phv_in_data_147(outp_io_phv_in_data_147),
    .io_phv_in_data_148(outp_io_phv_in_data_148),
    .io_phv_in_data_149(outp_io_phv_in_data_149),
    .io_phv_in_data_150(outp_io_phv_in_data_150),
    .io_phv_in_data_151(outp_io_phv_in_data_151),
    .io_phv_in_data_152(outp_io_phv_in_data_152),
    .io_phv_in_data_153(outp_io_phv_in_data_153),
    .io_phv_in_data_154(outp_io_phv_in_data_154),
    .io_phv_in_data_155(outp_io_phv_in_data_155),
    .io_phv_in_data_156(outp_io_phv_in_data_156),
    .io_phv_in_data_157(outp_io_phv_in_data_157),
    .io_phv_in_data_158(outp_io_phv_in_data_158),
    .io_phv_in_data_159(outp_io_phv_in_data_159),
    .io_phv_in_data_160(outp_io_phv_in_data_160),
    .io_phv_in_data_161(outp_io_phv_in_data_161),
    .io_phv_in_data_162(outp_io_phv_in_data_162),
    .io_phv_in_data_163(outp_io_phv_in_data_163),
    .io_phv_in_data_164(outp_io_phv_in_data_164),
    .io_phv_in_data_165(outp_io_phv_in_data_165),
    .io_phv_in_data_166(outp_io_phv_in_data_166),
    .io_phv_in_data_167(outp_io_phv_in_data_167),
    .io_phv_in_data_168(outp_io_phv_in_data_168),
    .io_phv_in_data_169(outp_io_phv_in_data_169),
    .io_phv_in_data_170(outp_io_phv_in_data_170),
    .io_phv_in_data_171(outp_io_phv_in_data_171),
    .io_phv_in_data_172(outp_io_phv_in_data_172),
    .io_phv_in_data_173(outp_io_phv_in_data_173),
    .io_phv_in_data_174(outp_io_phv_in_data_174),
    .io_phv_in_data_175(outp_io_phv_in_data_175),
    .io_phv_in_data_176(outp_io_phv_in_data_176),
    .io_phv_in_data_177(outp_io_phv_in_data_177),
    .io_phv_in_data_178(outp_io_phv_in_data_178),
    .io_phv_in_data_179(outp_io_phv_in_data_179),
    .io_phv_in_data_180(outp_io_phv_in_data_180),
    .io_phv_in_data_181(outp_io_phv_in_data_181),
    .io_phv_in_data_182(outp_io_phv_in_data_182),
    .io_phv_in_data_183(outp_io_phv_in_data_183),
    .io_phv_in_data_184(outp_io_phv_in_data_184),
    .io_phv_in_data_185(outp_io_phv_in_data_185),
    .io_phv_in_data_186(outp_io_phv_in_data_186),
    .io_phv_in_data_187(outp_io_phv_in_data_187),
    .io_phv_in_data_188(outp_io_phv_in_data_188),
    .io_phv_in_data_189(outp_io_phv_in_data_189),
    .io_phv_in_data_190(outp_io_phv_in_data_190),
    .io_phv_in_data_191(outp_io_phv_in_data_191),
    .io_phv_in_data_192(outp_io_phv_in_data_192),
    .io_phv_in_data_193(outp_io_phv_in_data_193),
    .io_phv_in_data_194(outp_io_phv_in_data_194),
    .io_phv_in_data_195(outp_io_phv_in_data_195),
    .io_phv_in_data_196(outp_io_phv_in_data_196),
    .io_phv_in_data_197(outp_io_phv_in_data_197),
    .io_phv_in_data_198(outp_io_phv_in_data_198),
    .io_phv_in_data_199(outp_io_phv_in_data_199),
    .io_phv_in_data_200(outp_io_phv_in_data_200),
    .io_phv_in_data_201(outp_io_phv_in_data_201),
    .io_phv_in_data_202(outp_io_phv_in_data_202),
    .io_phv_in_data_203(outp_io_phv_in_data_203),
    .io_phv_in_data_204(outp_io_phv_in_data_204),
    .io_phv_in_data_205(outp_io_phv_in_data_205),
    .io_phv_in_data_206(outp_io_phv_in_data_206),
    .io_phv_in_data_207(outp_io_phv_in_data_207),
    .io_phv_in_data_208(outp_io_phv_in_data_208),
    .io_phv_in_data_209(outp_io_phv_in_data_209),
    .io_phv_in_data_210(outp_io_phv_in_data_210),
    .io_phv_in_data_211(outp_io_phv_in_data_211),
    .io_phv_in_data_212(outp_io_phv_in_data_212),
    .io_phv_in_data_213(outp_io_phv_in_data_213),
    .io_phv_in_data_214(outp_io_phv_in_data_214),
    .io_phv_in_data_215(outp_io_phv_in_data_215),
    .io_phv_in_data_216(outp_io_phv_in_data_216),
    .io_phv_in_data_217(outp_io_phv_in_data_217),
    .io_phv_in_data_218(outp_io_phv_in_data_218),
    .io_phv_in_data_219(outp_io_phv_in_data_219),
    .io_phv_in_data_220(outp_io_phv_in_data_220),
    .io_phv_in_data_221(outp_io_phv_in_data_221),
    .io_phv_in_data_222(outp_io_phv_in_data_222),
    .io_phv_in_data_223(outp_io_phv_in_data_223),
    .io_phv_in_data_224(outp_io_phv_in_data_224),
    .io_phv_in_data_225(outp_io_phv_in_data_225),
    .io_phv_in_data_226(outp_io_phv_in_data_226),
    .io_phv_in_data_227(outp_io_phv_in_data_227),
    .io_phv_in_data_228(outp_io_phv_in_data_228),
    .io_phv_in_data_229(outp_io_phv_in_data_229),
    .io_phv_in_data_230(outp_io_phv_in_data_230),
    .io_phv_in_data_231(outp_io_phv_in_data_231),
    .io_phv_in_data_232(outp_io_phv_in_data_232),
    .io_phv_in_data_233(outp_io_phv_in_data_233),
    .io_phv_in_data_234(outp_io_phv_in_data_234),
    .io_phv_in_data_235(outp_io_phv_in_data_235),
    .io_phv_in_data_236(outp_io_phv_in_data_236),
    .io_phv_in_data_237(outp_io_phv_in_data_237),
    .io_phv_in_data_238(outp_io_phv_in_data_238),
    .io_phv_in_data_239(outp_io_phv_in_data_239),
    .io_phv_in_data_240(outp_io_phv_in_data_240),
    .io_phv_in_data_241(outp_io_phv_in_data_241),
    .io_phv_in_data_242(outp_io_phv_in_data_242),
    .io_phv_in_data_243(outp_io_phv_in_data_243),
    .io_phv_in_data_244(outp_io_phv_in_data_244),
    .io_phv_in_data_245(outp_io_phv_in_data_245),
    .io_phv_in_data_246(outp_io_phv_in_data_246),
    .io_phv_in_data_247(outp_io_phv_in_data_247),
    .io_phv_in_data_248(outp_io_phv_in_data_248),
    .io_phv_in_data_249(outp_io_phv_in_data_249),
    .io_phv_in_data_250(outp_io_phv_in_data_250),
    .io_phv_in_data_251(outp_io_phv_in_data_251),
    .io_phv_in_data_252(outp_io_phv_in_data_252),
    .io_phv_in_data_253(outp_io_phv_in_data_253),
    .io_phv_in_data_254(outp_io_phv_in_data_254),
    .io_phv_in_data_255(outp_io_phv_in_data_255),
    .io_pcie_o_cs(outp_io_pcie_o_cs),
    .io_pcie_o_r_en(outp_io_pcie_o_r_en),
    .io_pcie_o_r_addr(outp_io_pcie_o_r_addr),
    .io_pcie_o_r_data(outp_io_pcie_o_r_data)
  );
  InPort inp ( // @[ipsa_pcie.scala 16:22]
    .clock(inp_clock),
    .reset(inp_reset),
    .io_phv_out_data_0(inp_io_phv_out_data_0),
    .io_phv_out_data_1(inp_io_phv_out_data_1),
    .io_phv_out_data_2(inp_io_phv_out_data_2),
    .io_phv_out_data_3(inp_io_phv_out_data_3),
    .io_phv_out_data_4(inp_io_phv_out_data_4),
    .io_phv_out_data_5(inp_io_phv_out_data_5),
    .io_phv_out_data_6(inp_io_phv_out_data_6),
    .io_phv_out_data_7(inp_io_phv_out_data_7),
    .io_phv_out_data_8(inp_io_phv_out_data_8),
    .io_phv_out_data_9(inp_io_phv_out_data_9),
    .io_phv_out_data_10(inp_io_phv_out_data_10),
    .io_phv_out_data_11(inp_io_phv_out_data_11),
    .io_phv_out_data_12(inp_io_phv_out_data_12),
    .io_phv_out_data_13(inp_io_phv_out_data_13),
    .io_phv_out_data_14(inp_io_phv_out_data_14),
    .io_phv_out_data_15(inp_io_phv_out_data_15),
    .io_phv_out_data_16(inp_io_phv_out_data_16),
    .io_phv_out_data_17(inp_io_phv_out_data_17),
    .io_phv_out_data_18(inp_io_phv_out_data_18),
    .io_phv_out_data_19(inp_io_phv_out_data_19),
    .io_phv_out_data_20(inp_io_phv_out_data_20),
    .io_phv_out_data_21(inp_io_phv_out_data_21),
    .io_phv_out_data_22(inp_io_phv_out_data_22),
    .io_phv_out_data_23(inp_io_phv_out_data_23),
    .io_phv_out_data_24(inp_io_phv_out_data_24),
    .io_phv_out_data_25(inp_io_phv_out_data_25),
    .io_phv_out_data_26(inp_io_phv_out_data_26),
    .io_phv_out_data_27(inp_io_phv_out_data_27),
    .io_phv_out_data_28(inp_io_phv_out_data_28),
    .io_phv_out_data_29(inp_io_phv_out_data_29),
    .io_phv_out_data_30(inp_io_phv_out_data_30),
    .io_phv_out_data_31(inp_io_phv_out_data_31),
    .io_phv_out_data_32(inp_io_phv_out_data_32),
    .io_phv_out_data_33(inp_io_phv_out_data_33),
    .io_phv_out_data_34(inp_io_phv_out_data_34),
    .io_phv_out_data_35(inp_io_phv_out_data_35),
    .io_phv_out_data_36(inp_io_phv_out_data_36),
    .io_phv_out_data_37(inp_io_phv_out_data_37),
    .io_phv_out_data_38(inp_io_phv_out_data_38),
    .io_phv_out_data_39(inp_io_phv_out_data_39),
    .io_phv_out_data_40(inp_io_phv_out_data_40),
    .io_phv_out_data_41(inp_io_phv_out_data_41),
    .io_phv_out_data_42(inp_io_phv_out_data_42),
    .io_phv_out_data_43(inp_io_phv_out_data_43),
    .io_phv_out_data_44(inp_io_phv_out_data_44),
    .io_phv_out_data_45(inp_io_phv_out_data_45),
    .io_phv_out_data_46(inp_io_phv_out_data_46),
    .io_phv_out_data_47(inp_io_phv_out_data_47),
    .io_phv_out_data_48(inp_io_phv_out_data_48),
    .io_phv_out_data_49(inp_io_phv_out_data_49),
    .io_phv_out_data_50(inp_io_phv_out_data_50),
    .io_phv_out_data_51(inp_io_phv_out_data_51),
    .io_phv_out_data_52(inp_io_phv_out_data_52),
    .io_phv_out_data_53(inp_io_phv_out_data_53),
    .io_phv_out_data_54(inp_io_phv_out_data_54),
    .io_phv_out_data_55(inp_io_phv_out_data_55),
    .io_phv_out_data_56(inp_io_phv_out_data_56),
    .io_phv_out_data_57(inp_io_phv_out_data_57),
    .io_phv_out_data_58(inp_io_phv_out_data_58),
    .io_phv_out_data_59(inp_io_phv_out_data_59),
    .io_phv_out_data_60(inp_io_phv_out_data_60),
    .io_phv_out_data_61(inp_io_phv_out_data_61),
    .io_phv_out_data_62(inp_io_phv_out_data_62),
    .io_phv_out_data_63(inp_io_phv_out_data_63),
    .io_phv_out_data_64(inp_io_phv_out_data_64),
    .io_phv_out_data_65(inp_io_phv_out_data_65),
    .io_phv_out_data_66(inp_io_phv_out_data_66),
    .io_phv_out_data_67(inp_io_phv_out_data_67),
    .io_phv_out_data_68(inp_io_phv_out_data_68),
    .io_phv_out_data_69(inp_io_phv_out_data_69),
    .io_phv_out_data_70(inp_io_phv_out_data_70),
    .io_phv_out_data_71(inp_io_phv_out_data_71),
    .io_phv_out_data_72(inp_io_phv_out_data_72),
    .io_phv_out_data_73(inp_io_phv_out_data_73),
    .io_phv_out_data_74(inp_io_phv_out_data_74),
    .io_phv_out_data_75(inp_io_phv_out_data_75),
    .io_phv_out_data_76(inp_io_phv_out_data_76),
    .io_phv_out_data_77(inp_io_phv_out_data_77),
    .io_phv_out_data_78(inp_io_phv_out_data_78),
    .io_phv_out_data_79(inp_io_phv_out_data_79),
    .io_phv_out_data_80(inp_io_phv_out_data_80),
    .io_phv_out_data_81(inp_io_phv_out_data_81),
    .io_phv_out_data_82(inp_io_phv_out_data_82),
    .io_phv_out_data_83(inp_io_phv_out_data_83),
    .io_phv_out_data_84(inp_io_phv_out_data_84),
    .io_phv_out_data_85(inp_io_phv_out_data_85),
    .io_phv_out_data_86(inp_io_phv_out_data_86),
    .io_phv_out_data_87(inp_io_phv_out_data_87),
    .io_phv_out_data_88(inp_io_phv_out_data_88),
    .io_phv_out_data_89(inp_io_phv_out_data_89),
    .io_phv_out_data_90(inp_io_phv_out_data_90),
    .io_phv_out_data_91(inp_io_phv_out_data_91),
    .io_phv_out_data_92(inp_io_phv_out_data_92),
    .io_phv_out_data_93(inp_io_phv_out_data_93),
    .io_phv_out_data_94(inp_io_phv_out_data_94),
    .io_phv_out_data_95(inp_io_phv_out_data_95),
    .io_phv_out_data_96(inp_io_phv_out_data_96),
    .io_phv_out_data_97(inp_io_phv_out_data_97),
    .io_phv_out_data_98(inp_io_phv_out_data_98),
    .io_phv_out_data_99(inp_io_phv_out_data_99),
    .io_phv_out_data_100(inp_io_phv_out_data_100),
    .io_phv_out_data_101(inp_io_phv_out_data_101),
    .io_phv_out_data_102(inp_io_phv_out_data_102),
    .io_phv_out_data_103(inp_io_phv_out_data_103),
    .io_phv_out_data_104(inp_io_phv_out_data_104),
    .io_phv_out_data_105(inp_io_phv_out_data_105),
    .io_phv_out_data_106(inp_io_phv_out_data_106),
    .io_phv_out_data_107(inp_io_phv_out_data_107),
    .io_phv_out_data_108(inp_io_phv_out_data_108),
    .io_phv_out_data_109(inp_io_phv_out_data_109),
    .io_phv_out_data_110(inp_io_phv_out_data_110),
    .io_phv_out_data_111(inp_io_phv_out_data_111),
    .io_phv_out_data_112(inp_io_phv_out_data_112),
    .io_phv_out_data_113(inp_io_phv_out_data_113),
    .io_phv_out_data_114(inp_io_phv_out_data_114),
    .io_phv_out_data_115(inp_io_phv_out_data_115),
    .io_phv_out_data_116(inp_io_phv_out_data_116),
    .io_phv_out_data_117(inp_io_phv_out_data_117),
    .io_phv_out_data_118(inp_io_phv_out_data_118),
    .io_phv_out_data_119(inp_io_phv_out_data_119),
    .io_phv_out_data_120(inp_io_phv_out_data_120),
    .io_phv_out_data_121(inp_io_phv_out_data_121),
    .io_phv_out_data_122(inp_io_phv_out_data_122),
    .io_phv_out_data_123(inp_io_phv_out_data_123),
    .io_phv_out_data_124(inp_io_phv_out_data_124),
    .io_phv_out_data_125(inp_io_phv_out_data_125),
    .io_phv_out_data_126(inp_io_phv_out_data_126),
    .io_phv_out_data_127(inp_io_phv_out_data_127),
    .io_phv_out_data_128(inp_io_phv_out_data_128),
    .io_phv_out_data_129(inp_io_phv_out_data_129),
    .io_phv_out_data_130(inp_io_phv_out_data_130),
    .io_phv_out_data_131(inp_io_phv_out_data_131),
    .io_phv_out_data_132(inp_io_phv_out_data_132),
    .io_phv_out_data_133(inp_io_phv_out_data_133),
    .io_phv_out_data_134(inp_io_phv_out_data_134),
    .io_phv_out_data_135(inp_io_phv_out_data_135),
    .io_phv_out_data_136(inp_io_phv_out_data_136),
    .io_phv_out_data_137(inp_io_phv_out_data_137),
    .io_phv_out_data_138(inp_io_phv_out_data_138),
    .io_phv_out_data_139(inp_io_phv_out_data_139),
    .io_phv_out_data_140(inp_io_phv_out_data_140),
    .io_phv_out_data_141(inp_io_phv_out_data_141),
    .io_phv_out_data_142(inp_io_phv_out_data_142),
    .io_phv_out_data_143(inp_io_phv_out_data_143),
    .io_phv_out_data_144(inp_io_phv_out_data_144),
    .io_phv_out_data_145(inp_io_phv_out_data_145),
    .io_phv_out_data_146(inp_io_phv_out_data_146),
    .io_phv_out_data_147(inp_io_phv_out_data_147),
    .io_phv_out_data_148(inp_io_phv_out_data_148),
    .io_phv_out_data_149(inp_io_phv_out_data_149),
    .io_phv_out_data_150(inp_io_phv_out_data_150),
    .io_phv_out_data_151(inp_io_phv_out_data_151),
    .io_phv_out_data_152(inp_io_phv_out_data_152),
    .io_phv_out_data_153(inp_io_phv_out_data_153),
    .io_phv_out_data_154(inp_io_phv_out_data_154),
    .io_phv_out_data_155(inp_io_phv_out_data_155),
    .io_phv_out_data_156(inp_io_phv_out_data_156),
    .io_phv_out_data_157(inp_io_phv_out_data_157),
    .io_phv_out_data_158(inp_io_phv_out_data_158),
    .io_phv_out_data_159(inp_io_phv_out_data_159),
    .io_phv_out_data_160(inp_io_phv_out_data_160),
    .io_phv_out_data_161(inp_io_phv_out_data_161),
    .io_phv_out_data_162(inp_io_phv_out_data_162),
    .io_phv_out_data_163(inp_io_phv_out_data_163),
    .io_phv_out_data_164(inp_io_phv_out_data_164),
    .io_phv_out_data_165(inp_io_phv_out_data_165),
    .io_phv_out_data_166(inp_io_phv_out_data_166),
    .io_phv_out_data_167(inp_io_phv_out_data_167),
    .io_phv_out_data_168(inp_io_phv_out_data_168),
    .io_phv_out_data_169(inp_io_phv_out_data_169),
    .io_phv_out_data_170(inp_io_phv_out_data_170),
    .io_phv_out_data_171(inp_io_phv_out_data_171),
    .io_phv_out_data_172(inp_io_phv_out_data_172),
    .io_phv_out_data_173(inp_io_phv_out_data_173),
    .io_phv_out_data_174(inp_io_phv_out_data_174),
    .io_phv_out_data_175(inp_io_phv_out_data_175),
    .io_phv_out_data_176(inp_io_phv_out_data_176),
    .io_phv_out_data_177(inp_io_phv_out_data_177),
    .io_phv_out_data_178(inp_io_phv_out_data_178),
    .io_phv_out_data_179(inp_io_phv_out_data_179),
    .io_phv_out_data_180(inp_io_phv_out_data_180),
    .io_phv_out_data_181(inp_io_phv_out_data_181),
    .io_phv_out_data_182(inp_io_phv_out_data_182),
    .io_phv_out_data_183(inp_io_phv_out_data_183),
    .io_phv_out_data_184(inp_io_phv_out_data_184),
    .io_phv_out_data_185(inp_io_phv_out_data_185),
    .io_phv_out_data_186(inp_io_phv_out_data_186),
    .io_phv_out_data_187(inp_io_phv_out_data_187),
    .io_phv_out_data_188(inp_io_phv_out_data_188),
    .io_phv_out_data_189(inp_io_phv_out_data_189),
    .io_phv_out_data_190(inp_io_phv_out_data_190),
    .io_phv_out_data_191(inp_io_phv_out_data_191)
  );
  assign io_pcie_r_data = pcie_io_pcie_r_data; // @[ipsa_pcie.scala 20:20]
  assign ipsa_clock = clock;
  assign ipsa_io_pipe_phv_in_data_0 = inp_io_phv_out_data_0; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_1 = inp_io_phv_out_data_1; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_2 = inp_io_phv_out_data_2; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_3 = inp_io_phv_out_data_3; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_4 = inp_io_phv_out_data_4; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_5 = inp_io_phv_out_data_5; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_6 = inp_io_phv_out_data_6; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_7 = inp_io_phv_out_data_7; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_8 = inp_io_phv_out_data_8; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_9 = inp_io_phv_out_data_9; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_10 = inp_io_phv_out_data_10; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_11 = inp_io_phv_out_data_11; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_12 = inp_io_phv_out_data_12; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_13 = inp_io_phv_out_data_13; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_14 = inp_io_phv_out_data_14; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_15 = inp_io_phv_out_data_15; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_16 = inp_io_phv_out_data_16; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_17 = inp_io_phv_out_data_17; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_18 = inp_io_phv_out_data_18; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_19 = inp_io_phv_out_data_19; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_20 = inp_io_phv_out_data_20; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_21 = inp_io_phv_out_data_21; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_22 = inp_io_phv_out_data_22; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_23 = inp_io_phv_out_data_23; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_24 = inp_io_phv_out_data_24; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_25 = inp_io_phv_out_data_25; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_26 = inp_io_phv_out_data_26; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_27 = inp_io_phv_out_data_27; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_28 = inp_io_phv_out_data_28; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_29 = inp_io_phv_out_data_29; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_30 = inp_io_phv_out_data_30; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_31 = inp_io_phv_out_data_31; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_32 = inp_io_phv_out_data_32; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_33 = inp_io_phv_out_data_33; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_34 = inp_io_phv_out_data_34; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_35 = inp_io_phv_out_data_35; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_36 = inp_io_phv_out_data_36; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_37 = inp_io_phv_out_data_37; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_38 = inp_io_phv_out_data_38; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_39 = inp_io_phv_out_data_39; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_40 = inp_io_phv_out_data_40; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_41 = inp_io_phv_out_data_41; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_42 = inp_io_phv_out_data_42; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_43 = inp_io_phv_out_data_43; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_44 = inp_io_phv_out_data_44; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_45 = inp_io_phv_out_data_45; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_46 = inp_io_phv_out_data_46; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_47 = inp_io_phv_out_data_47; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_48 = inp_io_phv_out_data_48; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_49 = inp_io_phv_out_data_49; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_50 = inp_io_phv_out_data_50; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_51 = inp_io_phv_out_data_51; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_52 = inp_io_phv_out_data_52; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_53 = inp_io_phv_out_data_53; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_54 = inp_io_phv_out_data_54; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_55 = inp_io_phv_out_data_55; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_56 = inp_io_phv_out_data_56; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_57 = inp_io_phv_out_data_57; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_58 = inp_io_phv_out_data_58; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_59 = inp_io_phv_out_data_59; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_60 = inp_io_phv_out_data_60; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_61 = inp_io_phv_out_data_61; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_62 = inp_io_phv_out_data_62; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_63 = inp_io_phv_out_data_63; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_64 = inp_io_phv_out_data_64; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_65 = inp_io_phv_out_data_65; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_66 = inp_io_phv_out_data_66; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_67 = inp_io_phv_out_data_67; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_68 = inp_io_phv_out_data_68; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_69 = inp_io_phv_out_data_69; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_70 = inp_io_phv_out_data_70; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_71 = inp_io_phv_out_data_71; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_72 = inp_io_phv_out_data_72; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_73 = inp_io_phv_out_data_73; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_74 = inp_io_phv_out_data_74; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_75 = inp_io_phv_out_data_75; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_76 = inp_io_phv_out_data_76; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_77 = inp_io_phv_out_data_77; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_78 = inp_io_phv_out_data_78; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_79 = inp_io_phv_out_data_79; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_80 = inp_io_phv_out_data_80; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_81 = inp_io_phv_out_data_81; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_82 = inp_io_phv_out_data_82; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_83 = inp_io_phv_out_data_83; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_84 = inp_io_phv_out_data_84; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_85 = inp_io_phv_out_data_85; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_86 = inp_io_phv_out_data_86; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_87 = inp_io_phv_out_data_87; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_88 = inp_io_phv_out_data_88; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_89 = inp_io_phv_out_data_89; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_90 = inp_io_phv_out_data_90; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_91 = inp_io_phv_out_data_91; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_92 = inp_io_phv_out_data_92; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_93 = inp_io_phv_out_data_93; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_94 = inp_io_phv_out_data_94; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_95 = inp_io_phv_out_data_95; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_96 = inp_io_phv_out_data_96; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_97 = inp_io_phv_out_data_97; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_98 = inp_io_phv_out_data_98; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_99 = inp_io_phv_out_data_99; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_100 = inp_io_phv_out_data_100; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_101 = inp_io_phv_out_data_101; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_102 = inp_io_phv_out_data_102; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_103 = inp_io_phv_out_data_103; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_104 = inp_io_phv_out_data_104; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_105 = inp_io_phv_out_data_105; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_106 = inp_io_phv_out_data_106; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_107 = inp_io_phv_out_data_107; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_108 = inp_io_phv_out_data_108; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_109 = inp_io_phv_out_data_109; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_110 = inp_io_phv_out_data_110; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_111 = inp_io_phv_out_data_111; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_112 = inp_io_phv_out_data_112; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_113 = inp_io_phv_out_data_113; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_114 = inp_io_phv_out_data_114; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_115 = inp_io_phv_out_data_115; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_116 = inp_io_phv_out_data_116; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_117 = inp_io_phv_out_data_117; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_118 = inp_io_phv_out_data_118; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_119 = inp_io_phv_out_data_119; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_120 = inp_io_phv_out_data_120; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_121 = inp_io_phv_out_data_121; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_122 = inp_io_phv_out_data_122; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_123 = inp_io_phv_out_data_123; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_124 = inp_io_phv_out_data_124; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_125 = inp_io_phv_out_data_125; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_126 = inp_io_phv_out_data_126; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_127 = inp_io_phv_out_data_127; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_128 = inp_io_phv_out_data_128; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_129 = inp_io_phv_out_data_129; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_130 = inp_io_phv_out_data_130; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_131 = inp_io_phv_out_data_131; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_132 = inp_io_phv_out_data_132; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_133 = inp_io_phv_out_data_133; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_134 = inp_io_phv_out_data_134; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_135 = inp_io_phv_out_data_135; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_136 = inp_io_phv_out_data_136; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_137 = inp_io_phv_out_data_137; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_138 = inp_io_phv_out_data_138; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_139 = inp_io_phv_out_data_139; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_140 = inp_io_phv_out_data_140; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_141 = inp_io_phv_out_data_141; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_142 = inp_io_phv_out_data_142; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_143 = inp_io_phv_out_data_143; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_144 = inp_io_phv_out_data_144; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_145 = inp_io_phv_out_data_145; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_146 = inp_io_phv_out_data_146; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_147 = inp_io_phv_out_data_147; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_148 = inp_io_phv_out_data_148; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_149 = inp_io_phv_out_data_149; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_150 = inp_io_phv_out_data_150; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_151 = inp_io_phv_out_data_151; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_152 = inp_io_phv_out_data_152; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_153 = inp_io_phv_out_data_153; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_154 = inp_io_phv_out_data_154; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_155 = inp_io_phv_out_data_155; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_156 = inp_io_phv_out_data_156; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_157 = inp_io_phv_out_data_157; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_158 = inp_io_phv_out_data_158; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_159 = inp_io_phv_out_data_159; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_160 = inp_io_phv_out_data_160; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_161 = inp_io_phv_out_data_161; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_162 = inp_io_phv_out_data_162; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_163 = inp_io_phv_out_data_163; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_164 = inp_io_phv_out_data_164; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_165 = inp_io_phv_out_data_165; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_166 = inp_io_phv_out_data_166; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_167 = inp_io_phv_out_data_167; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_168 = inp_io_phv_out_data_168; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_169 = inp_io_phv_out_data_169; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_170 = inp_io_phv_out_data_170; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_171 = inp_io_phv_out_data_171; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_172 = inp_io_phv_out_data_172; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_173 = inp_io_phv_out_data_173; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_174 = inp_io_phv_out_data_174; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_175 = inp_io_phv_out_data_175; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_176 = inp_io_phv_out_data_176; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_177 = inp_io_phv_out_data_177; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_178 = inp_io_phv_out_data_178; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_179 = inp_io_phv_out_data_179; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_180 = inp_io_phv_out_data_180; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_181 = inp_io_phv_out_data_181; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_182 = inp_io_phv_out_data_182; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_183 = inp_io_phv_out_data_183; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_184 = inp_io_phv_out_data_184; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_185 = inp_io_phv_out_data_185; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_186 = inp_io_phv_out_data_186; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_187 = inp_io_phv_out_data_187; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_188 = inp_io_phv_out_data_188; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_189 = inp_io_phv_out_data_189; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_190 = inp_io_phv_out_data_190; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_pipe_phv_in_data_191 = inp_io_phv_out_data_191; // @[ipsa_pcie.scala 18:26]
  assign ipsa_io_mod_proc_mod_0_par_mod_en = pcie_io_mod_proc_mod_0_par_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_last_mau_id_mod = pcie_io_mod_proc_mod_0_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_last_mau_id = pcie_io_mod_proc_mod_0_par_mod_last_mau_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_cs = pcie_io_mod_proc_mod_0_par_mod_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_module_mod_state_id_mod = pcie_io_mod_proc_mod_0_par_mod_module_mod_state_id_mod
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_module_mod_state_id = pcie_io_mod_proc_mod_0_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs = pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_en = pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr = pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_par_mod_module_mod_sram_w_data = pcie_io_mod_proc_mod_0_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_en = pcie_io_mod_proc_mod_0_mat_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_config_id = pcie_io_mod_proc_mod_0_mat_mod_config_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_key_mod_header_id = pcie_io_mod_proc_mod_0_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_key_mod_internal_offset = pcie_io_mod_proc_mod_0_mat_mod_key_mod_internal_offset
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_key_mod_key_length = pcie_io_mod_proc_mod_0_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63 =
    pcie_io_mod_proc_mod_0_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_table_width = pcie_io_mod_proc_mod_0_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_mat_mod_table_mod_table_depth = pcie_io_mod_proc_mod_0_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_act_mod_en_0 = pcie_io_mod_proc_mod_0_act_mod_en_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_act_mod_en_1 = pcie_io_mod_proc_mod_0_act_mod_en_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_act_mod_addr = pcie_io_mod_proc_mod_0_act_mod_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_act_mod_data_0 = pcie_io_mod_proc_mod_0_act_mod_data_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_0_act_mod_data_1 = pcie_io_mod_proc_mod_0_act_mod_data_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_en = pcie_io_mod_proc_mod_1_par_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_last_mau_id_mod = pcie_io_mod_proc_mod_1_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_last_mau_id = pcie_io_mod_proc_mod_1_par_mod_last_mau_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_cs = pcie_io_mod_proc_mod_1_par_mod_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_module_mod_state_id_mod = pcie_io_mod_proc_mod_1_par_mod_module_mod_state_id_mod
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_module_mod_state_id = pcie_io_mod_proc_mod_1_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs = pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_en = pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr = pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_par_mod_module_mod_sram_w_data = pcie_io_mod_proc_mod_1_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_en = pcie_io_mod_proc_mod_1_mat_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_config_id = pcie_io_mod_proc_mod_1_mat_mod_config_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_key_mod_header_id = pcie_io_mod_proc_mod_1_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_key_mod_internal_offset = pcie_io_mod_proc_mod_1_mat_mod_key_mod_internal_offset
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_key_mod_key_length = pcie_io_mod_proc_mod_1_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63 =
    pcie_io_mod_proc_mod_1_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_table_width = pcie_io_mod_proc_mod_1_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_mat_mod_table_mod_table_depth = pcie_io_mod_proc_mod_1_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_act_mod_en_0 = pcie_io_mod_proc_mod_1_act_mod_en_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_act_mod_en_1 = pcie_io_mod_proc_mod_1_act_mod_en_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_act_mod_addr = pcie_io_mod_proc_mod_1_act_mod_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_act_mod_data_0 = pcie_io_mod_proc_mod_1_act_mod_data_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_1_act_mod_data_1 = pcie_io_mod_proc_mod_1_act_mod_data_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_en = pcie_io_mod_proc_mod_2_par_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_last_mau_id_mod = pcie_io_mod_proc_mod_2_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_last_mau_id = pcie_io_mod_proc_mod_2_par_mod_last_mau_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_cs = pcie_io_mod_proc_mod_2_par_mod_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_module_mod_state_id_mod = pcie_io_mod_proc_mod_2_par_mod_module_mod_state_id_mod
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_module_mod_state_id = pcie_io_mod_proc_mod_2_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs = pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_en = pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr = pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_par_mod_module_mod_sram_w_data = pcie_io_mod_proc_mod_2_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_en = pcie_io_mod_proc_mod_2_mat_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_config_id = pcie_io_mod_proc_mod_2_mat_mod_config_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_key_mod_header_id = pcie_io_mod_proc_mod_2_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_key_mod_internal_offset = pcie_io_mod_proc_mod_2_mat_mod_key_mod_internal_offset
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_key_mod_key_length = pcie_io_mod_proc_mod_2_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63 =
    pcie_io_mod_proc_mod_2_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_table_width = pcie_io_mod_proc_mod_2_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_mat_mod_table_mod_table_depth = pcie_io_mod_proc_mod_2_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_act_mod_en_0 = pcie_io_mod_proc_mod_2_act_mod_en_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_act_mod_en_1 = pcie_io_mod_proc_mod_2_act_mod_en_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_act_mod_addr = pcie_io_mod_proc_mod_2_act_mod_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_act_mod_data_0 = pcie_io_mod_proc_mod_2_act_mod_data_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_2_act_mod_data_1 = pcie_io_mod_proc_mod_2_act_mod_data_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_en = pcie_io_mod_proc_mod_3_par_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_last_mau_id_mod = pcie_io_mod_proc_mod_3_par_mod_last_mau_id_mod; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_last_mau_id = pcie_io_mod_proc_mod_3_par_mod_last_mau_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_cs = pcie_io_mod_proc_mod_3_par_mod_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_module_mod_state_id_mod = pcie_io_mod_proc_mod_3_par_mod_module_mod_state_id_mod
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_module_mod_state_id = pcie_io_mod_proc_mod_3_par_mod_module_mod_state_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs = pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_cs; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_en = pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr = pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_par_mod_module_mod_sram_w_data = pcie_io_mod_proc_mod_3_par_mod_module_mod_sram_w_data; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_en = pcie_io_mod_proc_mod_3_mat_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_config_id = pcie_io_mod_proc_mod_3_mat_mod_config_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_key_mod_header_id = pcie_io_mod_proc_mod_3_mat_mod_key_mod_header_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_key_mod_internal_offset = pcie_io_mod_proc_mod_3_mat_mod_key_mod_internal_offset
    ; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_key_mod_key_length = pcie_io_mod_proc_mod_3_mat_mod_key_mod_key_length; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_2; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_3; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_4; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_5; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_6; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_7; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_8; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_9; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_10; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_11; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_12; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_13; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_14; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_15; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_16; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_17; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_18; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_19; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_20; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_21; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_22; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_23; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_24; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_25; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_26; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_27; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_28; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_29; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_30; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_31; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_32; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_33; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_34; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_35; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_36; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_37; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_38; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_39; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_40; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_41; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_42; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_43; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_44; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_45; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_46; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_47; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_48; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_49; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_50; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_51; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_52; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_53; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_54; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_55; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_56; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_57; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_58; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_59; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_60; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_61; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_62; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63 =
    pcie_io_mod_proc_mod_3_mat_mod_table_mod_sram_id_table_63; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_table_width = pcie_io_mod_proc_mod_3_mat_mod_table_mod_table_width; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_mat_mod_table_mod_table_depth = pcie_io_mod_proc_mod_3_mat_mod_table_mod_table_depth; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_act_mod_en_0 = pcie_io_mod_proc_mod_3_act_mod_en_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_act_mod_en_1 = pcie_io_mod_proc_mod_3_act_mod_en_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_act_mod_addr = pcie_io_mod_proc_mod_3_act_mod_addr; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_act_mod_data_0 = pcie_io_mod_proc_mod_3_act_mod_data_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_proc_mod_3_act_mod_data_1 = pcie_io_mod_proc_mod_3_act_mod_data_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_xbar_mod_en = pcie_io_mod_xbar_mod_en; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_xbar_mod_first_proc_id = pcie_io_mod_xbar_mod_first_proc_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_xbar_mod_last_proc_id = pcie_io_mod_xbar_mod_last_proc_id; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_xbar_mod_next_proc_id_0 = pcie_io_mod_xbar_mod_next_proc_id_0; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_xbar_mod_next_proc_id_1 = pcie_io_mod_xbar_mod_next_proc_id_1; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_xbar_mod_next_proc_id_2 = pcie_io_mod_xbar_mod_next_proc_id_2; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_mod_xbar_mod_next_proc_id_3 = pcie_io_mod_xbar_mod_next_proc_id_3; // @[ipsa_pcie.scala 22:20]
  assign ipsa_io_w_0_wcs = pcie_io_w_0_wcs; // @[ipsa_pcie.scala 23:20]
  assign ipsa_io_w_0_w_en = pcie_io_w_0_w_en; // @[ipsa_pcie.scala 23:20]
  assign ipsa_io_w_0_w_addr = pcie_io_w_0_w_addr; // @[ipsa_pcie.scala 23:20]
  assign ipsa_io_w_0_w_data = pcie_io_w_0_w_data; // @[ipsa_pcie.scala 23:20]
  assign pcie_clock = clock;
  assign pcie_io_pcie_r_en = io_pcie_r_en; // @[ipsa_pcie.scala 20:20]
  assign pcie_io_pcie_r_addr = io_pcie_r_addr; // @[ipsa_pcie.scala 20:20]
  assign pcie_io_pcie_w_en = io_pcie_w_en; // @[ipsa_pcie.scala 21:20]
  assign pcie_io_pcie_w_addr = io_pcie_w_addr; // @[ipsa_pcie.scala 21:20]
  assign pcie_io_pcie_w_data = io_pcie_w_data; // @[ipsa_pcie.scala 21:20]
  assign pcie_io_pcie_o_r_data = outp_io_pcie_o_r_data; // @[ipsa_pcie.scala 26:26]
  assign outp_clock = clock;
  assign outp_io_phv_in_data_0 = ipsa_io_pipe_phv_out_data_0; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_1 = ipsa_io_pipe_phv_out_data_1; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_2 = ipsa_io_pipe_phv_out_data_2; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_3 = ipsa_io_pipe_phv_out_data_3; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_4 = ipsa_io_pipe_phv_out_data_4; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_5 = ipsa_io_pipe_phv_out_data_5; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_6 = ipsa_io_pipe_phv_out_data_6; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_7 = ipsa_io_pipe_phv_out_data_7; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_8 = ipsa_io_pipe_phv_out_data_8; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_9 = ipsa_io_pipe_phv_out_data_9; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_10 = ipsa_io_pipe_phv_out_data_10; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_11 = ipsa_io_pipe_phv_out_data_11; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_12 = ipsa_io_pipe_phv_out_data_12; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_13 = ipsa_io_pipe_phv_out_data_13; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_14 = ipsa_io_pipe_phv_out_data_14; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_15 = ipsa_io_pipe_phv_out_data_15; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_16 = ipsa_io_pipe_phv_out_data_16; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_17 = ipsa_io_pipe_phv_out_data_17; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_18 = ipsa_io_pipe_phv_out_data_18; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_19 = ipsa_io_pipe_phv_out_data_19; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_20 = ipsa_io_pipe_phv_out_data_20; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_21 = ipsa_io_pipe_phv_out_data_21; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_22 = ipsa_io_pipe_phv_out_data_22; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_23 = ipsa_io_pipe_phv_out_data_23; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_24 = ipsa_io_pipe_phv_out_data_24; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_25 = ipsa_io_pipe_phv_out_data_25; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_26 = ipsa_io_pipe_phv_out_data_26; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_27 = ipsa_io_pipe_phv_out_data_27; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_28 = ipsa_io_pipe_phv_out_data_28; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_29 = ipsa_io_pipe_phv_out_data_29; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_30 = ipsa_io_pipe_phv_out_data_30; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_31 = ipsa_io_pipe_phv_out_data_31; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_32 = ipsa_io_pipe_phv_out_data_32; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_33 = ipsa_io_pipe_phv_out_data_33; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_34 = ipsa_io_pipe_phv_out_data_34; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_35 = ipsa_io_pipe_phv_out_data_35; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_36 = ipsa_io_pipe_phv_out_data_36; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_37 = ipsa_io_pipe_phv_out_data_37; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_38 = ipsa_io_pipe_phv_out_data_38; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_39 = ipsa_io_pipe_phv_out_data_39; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_40 = ipsa_io_pipe_phv_out_data_40; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_41 = ipsa_io_pipe_phv_out_data_41; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_42 = ipsa_io_pipe_phv_out_data_42; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_43 = ipsa_io_pipe_phv_out_data_43; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_44 = ipsa_io_pipe_phv_out_data_44; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_45 = ipsa_io_pipe_phv_out_data_45; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_46 = ipsa_io_pipe_phv_out_data_46; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_47 = ipsa_io_pipe_phv_out_data_47; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_48 = ipsa_io_pipe_phv_out_data_48; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_49 = ipsa_io_pipe_phv_out_data_49; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_50 = ipsa_io_pipe_phv_out_data_50; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_51 = ipsa_io_pipe_phv_out_data_51; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_52 = ipsa_io_pipe_phv_out_data_52; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_53 = ipsa_io_pipe_phv_out_data_53; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_54 = ipsa_io_pipe_phv_out_data_54; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_55 = ipsa_io_pipe_phv_out_data_55; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_56 = ipsa_io_pipe_phv_out_data_56; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_57 = ipsa_io_pipe_phv_out_data_57; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_58 = ipsa_io_pipe_phv_out_data_58; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_59 = ipsa_io_pipe_phv_out_data_59; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_60 = ipsa_io_pipe_phv_out_data_60; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_61 = ipsa_io_pipe_phv_out_data_61; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_62 = ipsa_io_pipe_phv_out_data_62; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_63 = ipsa_io_pipe_phv_out_data_63; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_64 = ipsa_io_pipe_phv_out_data_64; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_65 = ipsa_io_pipe_phv_out_data_65; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_66 = ipsa_io_pipe_phv_out_data_66; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_67 = ipsa_io_pipe_phv_out_data_67; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_68 = ipsa_io_pipe_phv_out_data_68; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_69 = ipsa_io_pipe_phv_out_data_69; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_70 = ipsa_io_pipe_phv_out_data_70; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_71 = ipsa_io_pipe_phv_out_data_71; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_72 = ipsa_io_pipe_phv_out_data_72; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_73 = ipsa_io_pipe_phv_out_data_73; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_74 = ipsa_io_pipe_phv_out_data_74; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_75 = ipsa_io_pipe_phv_out_data_75; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_76 = ipsa_io_pipe_phv_out_data_76; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_77 = ipsa_io_pipe_phv_out_data_77; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_78 = ipsa_io_pipe_phv_out_data_78; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_79 = ipsa_io_pipe_phv_out_data_79; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_80 = ipsa_io_pipe_phv_out_data_80; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_81 = ipsa_io_pipe_phv_out_data_81; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_82 = ipsa_io_pipe_phv_out_data_82; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_83 = ipsa_io_pipe_phv_out_data_83; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_84 = ipsa_io_pipe_phv_out_data_84; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_85 = ipsa_io_pipe_phv_out_data_85; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_86 = ipsa_io_pipe_phv_out_data_86; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_87 = ipsa_io_pipe_phv_out_data_87; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_88 = ipsa_io_pipe_phv_out_data_88; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_89 = ipsa_io_pipe_phv_out_data_89; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_90 = ipsa_io_pipe_phv_out_data_90; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_91 = ipsa_io_pipe_phv_out_data_91; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_92 = ipsa_io_pipe_phv_out_data_92; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_93 = ipsa_io_pipe_phv_out_data_93; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_94 = ipsa_io_pipe_phv_out_data_94; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_95 = ipsa_io_pipe_phv_out_data_95; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_96 = ipsa_io_pipe_phv_out_data_96; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_97 = ipsa_io_pipe_phv_out_data_97; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_98 = ipsa_io_pipe_phv_out_data_98; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_99 = ipsa_io_pipe_phv_out_data_99; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_100 = ipsa_io_pipe_phv_out_data_100; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_101 = ipsa_io_pipe_phv_out_data_101; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_102 = ipsa_io_pipe_phv_out_data_102; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_103 = ipsa_io_pipe_phv_out_data_103; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_104 = ipsa_io_pipe_phv_out_data_104; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_105 = ipsa_io_pipe_phv_out_data_105; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_106 = ipsa_io_pipe_phv_out_data_106; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_107 = ipsa_io_pipe_phv_out_data_107; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_108 = ipsa_io_pipe_phv_out_data_108; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_109 = ipsa_io_pipe_phv_out_data_109; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_110 = ipsa_io_pipe_phv_out_data_110; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_111 = ipsa_io_pipe_phv_out_data_111; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_112 = ipsa_io_pipe_phv_out_data_112; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_113 = ipsa_io_pipe_phv_out_data_113; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_114 = ipsa_io_pipe_phv_out_data_114; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_115 = ipsa_io_pipe_phv_out_data_115; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_116 = ipsa_io_pipe_phv_out_data_116; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_117 = ipsa_io_pipe_phv_out_data_117; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_118 = ipsa_io_pipe_phv_out_data_118; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_119 = ipsa_io_pipe_phv_out_data_119; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_120 = ipsa_io_pipe_phv_out_data_120; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_121 = ipsa_io_pipe_phv_out_data_121; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_122 = ipsa_io_pipe_phv_out_data_122; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_123 = ipsa_io_pipe_phv_out_data_123; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_124 = ipsa_io_pipe_phv_out_data_124; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_125 = ipsa_io_pipe_phv_out_data_125; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_126 = ipsa_io_pipe_phv_out_data_126; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_127 = ipsa_io_pipe_phv_out_data_127; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_128 = ipsa_io_pipe_phv_out_data_128; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_129 = ipsa_io_pipe_phv_out_data_129; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_130 = ipsa_io_pipe_phv_out_data_130; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_131 = ipsa_io_pipe_phv_out_data_131; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_132 = ipsa_io_pipe_phv_out_data_132; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_133 = ipsa_io_pipe_phv_out_data_133; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_134 = ipsa_io_pipe_phv_out_data_134; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_135 = ipsa_io_pipe_phv_out_data_135; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_136 = ipsa_io_pipe_phv_out_data_136; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_137 = ipsa_io_pipe_phv_out_data_137; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_138 = ipsa_io_pipe_phv_out_data_138; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_139 = ipsa_io_pipe_phv_out_data_139; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_140 = ipsa_io_pipe_phv_out_data_140; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_141 = ipsa_io_pipe_phv_out_data_141; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_142 = ipsa_io_pipe_phv_out_data_142; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_143 = ipsa_io_pipe_phv_out_data_143; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_144 = ipsa_io_pipe_phv_out_data_144; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_145 = ipsa_io_pipe_phv_out_data_145; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_146 = ipsa_io_pipe_phv_out_data_146; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_147 = ipsa_io_pipe_phv_out_data_147; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_148 = ipsa_io_pipe_phv_out_data_148; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_149 = ipsa_io_pipe_phv_out_data_149; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_150 = ipsa_io_pipe_phv_out_data_150; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_151 = ipsa_io_pipe_phv_out_data_151; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_152 = ipsa_io_pipe_phv_out_data_152; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_153 = ipsa_io_pipe_phv_out_data_153; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_154 = ipsa_io_pipe_phv_out_data_154; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_155 = ipsa_io_pipe_phv_out_data_155; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_156 = ipsa_io_pipe_phv_out_data_156; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_157 = ipsa_io_pipe_phv_out_data_157; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_158 = ipsa_io_pipe_phv_out_data_158; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_159 = ipsa_io_pipe_phv_out_data_159; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_160 = ipsa_io_pipe_phv_out_data_160; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_161 = ipsa_io_pipe_phv_out_data_161; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_162 = ipsa_io_pipe_phv_out_data_162; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_163 = ipsa_io_pipe_phv_out_data_163; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_164 = ipsa_io_pipe_phv_out_data_164; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_165 = ipsa_io_pipe_phv_out_data_165; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_166 = ipsa_io_pipe_phv_out_data_166; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_167 = ipsa_io_pipe_phv_out_data_167; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_168 = ipsa_io_pipe_phv_out_data_168; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_169 = ipsa_io_pipe_phv_out_data_169; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_170 = ipsa_io_pipe_phv_out_data_170; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_171 = ipsa_io_pipe_phv_out_data_171; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_172 = ipsa_io_pipe_phv_out_data_172; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_173 = ipsa_io_pipe_phv_out_data_173; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_174 = ipsa_io_pipe_phv_out_data_174; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_175 = ipsa_io_pipe_phv_out_data_175; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_176 = ipsa_io_pipe_phv_out_data_176; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_177 = ipsa_io_pipe_phv_out_data_177; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_178 = ipsa_io_pipe_phv_out_data_178; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_179 = ipsa_io_pipe_phv_out_data_179; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_180 = ipsa_io_pipe_phv_out_data_180; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_181 = ipsa_io_pipe_phv_out_data_181; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_182 = ipsa_io_pipe_phv_out_data_182; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_183 = ipsa_io_pipe_phv_out_data_183; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_184 = ipsa_io_pipe_phv_out_data_184; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_185 = ipsa_io_pipe_phv_out_data_185; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_186 = ipsa_io_pipe_phv_out_data_186; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_187 = ipsa_io_pipe_phv_out_data_187; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_188 = ipsa_io_pipe_phv_out_data_188; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_189 = ipsa_io_pipe_phv_out_data_189; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_190 = ipsa_io_pipe_phv_out_data_190; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_191 = ipsa_io_pipe_phv_out_data_191; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_192 = ipsa_io_pipe_phv_out_data_192; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_193 = ipsa_io_pipe_phv_out_data_193; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_194 = ipsa_io_pipe_phv_out_data_194; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_195 = ipsa_io_pipe_phv_out_data_195; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_196 = ipsa_io_pipe_phv_out_data_196; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_197 = ipsa_io_pipe_phv_out_data_197; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_198 = ipsa_io_pipe_phv_out_data_198; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_199 = ipsa_io_pipe_phv_out_data_199; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_200 = ipsa_io_pipe_phv_out_data_200; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_201 = ipsa_io_pipe_phv_out_data_201; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_202 = ipsa_io_pipe_phv_out_data_202; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_203 = ipsa_io_pipe_phv_out_data_203; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_204 = ipsa_io_pipe_phv_out_data_204; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_205 = ipsa_io_pipe_phv_out_data_205; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_206 = ipsa_io_pipe_phv_out_data_206; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_207 = ipsa_io_pipe_phv_out_data_207; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_208 = ipsa_io_pipe_phv_out_data_208; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_209 = ipsa_io_pipe_phv_out_data_209; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_210 = ipsa_io_pipe_phv_out_data_210; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_211 = ipsa_io_pipe_phv_out_data_211; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_212 = ipsa_io_pipe_phv_out_data_212; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_213 = ipsa_io_pipe_phv_out_data_213; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_214 = ipsa_io_pipe_phv_out_data_214; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_215 = ipsa_io_pipe_phv_out_data_215; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_216 = ipsa_io_pipe_phv_out_data_216; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_217 = ipsa_io_pipe_phv_out_data_217; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_218 = ipsa_io_pipe_phv_out_data_218; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_219 = ipsa_io_pipe_phv_out_data_219; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_220 = ipsa_io_pipe_phv_out_data_220; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_221 = ipsa_io_pipe_phv_out_data_221; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_222 = ipsa_io_pipe_phv_out_data_222; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_223 = ipsa_io_pipe_phv_out_data_223; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_224 = ipsa_io_pipe_phv_out_data_224; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_225 = ipsa_io_pipe_phv_out_data_225; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_226 = ipsa_io_pipe_phv_out_data_226; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_227 = ipsa_io_pipe_phv_out_data_227; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_228 = ipsa_io_pipe_phv_out_data_228; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_229 = ipsa_io_pipe_phv_out_data_229; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_230 = ipsa_io_pipe_phv_out_data_230; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_231 = ipsa_io_pipe_phv_out_data_231; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_232 = ipsa_io_pipe_phv_out_data_232; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_233 = ipsa_io_pipe_phv_out_data_233; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_234 = ipsa_io_pipe_phv_out_data_234; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_235 = ipsa_io_pipe_phv_out_data_235; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_236 = ipsa_io_pipe_phv_out_data_236; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_237 = ipsa_io_pipe_phv_out_data_237; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_238 = ipsa_io_pipe_phv_out_data_238; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_239 = ipsa_io_pipe_phv_out_data_239; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_240 = ipsa_io_pipe_phv_out_data_240; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_241 = ipsa_io_pipe_phv_out_data_241; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_242 = ipsa_io_pipe_phv_out_data_242; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_243 = ipsa_io_pipe_phv_out_data_243; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_244 = ipsa_io_pipe_phv_out_data_244; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_245 = ipsa_io_pipe_phv_out_data_245; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_246 = ipsa_io_pipe_phv_out_data_246; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_247 = ipsa_io_pipe_phv_out_data_247; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_248 = ipsa_io_pipe_phv_out_data_248; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_249 = ipsa_io_pipe_phv_out_data_249; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_250 = ipsa_io_pipe_phv_out_data_250; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_251 = ipsa_io_pipe_phv_out_data_251; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_252 = ipsa_io_pipe_phv_out_data_252; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_253 = ipsa_io_pipe_phv_out_data_253; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_254 = ipsa_io_pipe_phv_out_data_254; // @[ipsa_pcie.scala 25:26]
  assign outp_io_phv_in_data_255 = ipsa_io_pipe_phv_out_data_255; // @[ipsa_pcie.scala 25:26]
  assign outp_io_pcie_o_cs = pcie_io_pcie_o_cs; // @[ipsa_pcie.scala 26:26]
  assign outp_io_pcie_o_r_en = pcie_io_pcie_o_r_en; // @[ipsa_pcie.scala 26:26]
  assign outp_io_pcie_o_r_addr = pcie_io_pcie_o_r_addr; // @[ipsa_pcie.scala 26:26]
  assign inp_clock = clock;
  assign inp_reset = reset;
endmodule
