module MatchGetKeyRaw(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [7:0]  io_key_config_0_key_length,
  input  [7:0]  io_key_config_1_key_length,
  input  [7:0]  io_key_offset_in,
  output [1:0]  io_bias_out,
  output [7:0]  io_match_key_bytes_0,
  output [7:0]  io_match_key_bytes_1,
  output [7:0]  io_match_key_bytes_2,
  output [7:0]  io_match_key_bytes_3,
  output [7:0]  io_match_key_bytes_4,
  output [7:0]  io_match_key_bytes_5,
  output [7:0]  io_match_key_bytes_6,
  output [7:0]  io_match_key_bytes_7,
  output [7:0]  io_match_key_bytes_8,
  output [7:0]  io_match_key_bytes_9,
  output [7:0]  io_match_key_bytes_10,
  output [7:0]  io_match_key_bytes_11,
  output [7:0]  io_match_key_bytes_12,
  output [7:0]  io_match_key_bytes_13,
  output [7:0]  io_match_key_bytes_14,
  output [7:0]  io_match_key_bytes_15,
  output [7:0]  io_match_key_bytes_16,
  output [7:0]  io_match_key_bytes_17,
  output [7:0]  io_match_key_bytes_18,
  output [7:0]  io_match_key_bytes_19,
  output [7:0]  io_match_key_bytes_20,
  output [7:0]  io_match_key_bytes_21,
  output [7:0]  io_match_key_bytes_22,
  output [7:0]  io_match_key_bytes_23
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 67:26]
  reg [7:0] phv_data_1; // @[matcher.scala 67:26]
  reg [7:0] phv_data_2; // @[matcher.scala 67:26]
  reg [7:0] phv_data_3; // @[matcher.scala 67:26]
  reg [7:0] phv_data_4; // @[matcher.scala 67:26]
  reg [7:0] phv_data_5; // @[matcher.scala 67:26]
  reg [7:0] phv_data_6; // @[matcher.scala 67:26]
  reg [7:0] phv_data_7; // @[matcher.scala 67:26]
  reg [7:0] phv_data_8; // @[matcher.scala 67:26]
  reg [7:0] phv_data_9; // @[matcher.scala 67:26]
  reg [7:0] phv_data_10; // @[matcher.scala 67:26]
  reg [7:0] phv_data_11; // @[matcher.scala 67:26]
  reg [7:0] phv_data_12; // @[matcher.scala 67:26]
  reg [7:0] phv_data_13; // @[matcher.scala 67:26]
  reg [7:0] phv_data_14; // @[matcher.scala 67:26]
  reg [7:0] phv_data_15; // @[matcher.scala 67:26]
  reg [7:0] phv_data_16; // @[matcher.scala 67:26]
  reg [7:0] phv_data_17; // @[matcher.scala 67:26]
  reg [7:0] phv_data_18; // @[matcher.scala 67:26]
  reg [7:0] phv_data_19; // @[matcher.scala 67:26]
  reg [7:0] phv_data_20; // @[matcher.scala 67:26]
  reg [7:0] phv_data_21; // @[matcher.scala 67:26]
  reg [7:0] phv_data_22; // @[matcher.scala 67:26]
  reg [7:0] phv_data_23; // @[matcher.scala 67:26]
  reg [7:0] phv_data_24; // @[matcher.scala 67:26]
  reg [7:0] phv_data_25; // @[matcher.scala 67:26]
  reg [7:0] phv_data_26; // @[matcher.scala 67:26]
  reg [7:0] phv_data_27; // @[matcher.scala 67:26]
  reg [7:0] phv_data_28; // @[matcher.scala 67:26]
  reg [7:0] phv_data_29; // @[matcher.scala 67:26]
  reg [7:0] phv_data_30; // @[matcher.scala 67:26]
  reg [7:0] phv_data_31; // @[matcher.scala 67:26]
  reg [7:0] phv_data_32; // @[matcher.scala 67:26]
  reg [7:0] phv_data_33; // @[matcher.scala 67:26]
  reg [7:0] phv_data_34; // @[matcher.scala 67:26]
  reg [7:0] phv_data_35; // @[matcher.scala 67:26]
  reg [7:0] phv_data_36; // @[matcher.scala 67:26]
  reg [7:0] phv_data_37; // @[matcher.scala 67:26]
  reg [7:0] phv_data_38; // @[matcher.scala 67:26]
  reg [7:0] phv_data_39; // @[matcher.scala 67:26]
  reg [7:0] phv_data_40; // @[matcher.scala 67:26]
  reg [7:0] phv_data_41; // @[matcher.scala 67:26]
  reg [7:0] phv_data_42; // @[matcher.scala 67:26]
  reg [7:0] phv_data_43; // @[matcher.scala 67:26]
  reg [7:0] phv_data_44; // @[matcher.scala 67:26]
  reg [7:0] phv_data_45; // @[matcher.scala 67:26]
  reg [7:0] phv_data_46; // @[matcher.scala 67:26]
  reg [7:0] phv_data_47; // @[matcher.scala 67:26]
  reg [7:0] phv_data_48; // @[matcher.scala 67:26]
  reg [7:0] phv_data_49; // @[matcher.scala 67:26]
  reg [7:0] phv_data_50; // @[matcher.scala 67:26]
  reg [7:0] phv_data_51; // @[matcher.scala 67:26]
  reg [7:0] phv_data_52; // @[matcher.scala 67:26]
  reg [7:0] phv_data_53; // @[matcher.scala 67:26]
  reg [7:0] phv_data_54; // @[matcher.scala 67:26]
  reg [7:0] phv_data_55; // @[matcher.scala 67:26]
  reg [7:0] phv_data_56; // @[matcher.scala 67:26]
  reg [7:0] phv_data_57; // @[matcher.scala 67:26]
  reg [7:0] phv_data_58; // @[matcher.scala 67:26]
  reg [7:0] phv_data_59; // @[matcher.scala 67:26]
  reg [7:0] phv_data_60; // @[matcher.scala 67:26]
  reg [7:0] phv_data_61; // @[matcher.scala 67:26]
  reg [7:0] phv_data_62; // @[matcher.scala 67:26]
  reg [7:0] phv_data_63; // @[matcher.scala 67:26]
  reg [7:0] phv_data_64; // @[matcher.scala 67:26]
  reg [7:0] phv_data_65; // @[matcher.scala 67:26]
  reg [7:0] phv_data_66; // @[matcher.scala 67:26]
  reg [7:0] phv_data_67; // @[matcher.scala 67:26]
  reg [7:0] phv_data_68; // @[matcher.scala 67:26]
  reg [7:0] phv_data_69; // @[matcher.scala 67:26]
  reg [7:0] phv_data_70; // @[matcher.scala 67:26]
  reg [7:0] phv_data_71; // @[matcher.scala 67:26]
  reg [7:0] phv_data_72; // @[matcher.scala 67:26]
  reg [7:0] phv_data_73; // @[matcher.scala 67:26]
  reg [7:0] phv_data_74; // @[matcher.scala 67:26]
  reg [7:0] phv_data_75; // @[matcher.scala 67:26]
  reg [7:0] phv_data_76; // @[matcher.scala 67:26]
  reg [7:0] phv_data_77; // @[matcher.scala 67:26]
  reg [7:0] phv_data_78; // @[matcher.scala 67:26]
  reg [7:0] phv_data_79; // @[matcher.scala 67:26]
  reg [7:0] phv_data_80; // @[matcher.scala 67:26]
  reg [7:0] phv_data_81; // @[matcher.scala 67:26]
  reg [7:0] phv_data_82; // @[matcher.scala 67:26]
  reg [7:0] phv_data_83; // @[matcher.scala 67:26]
  reg [7:0] phv_data_84; // @[matcher.scala 67:26]
  reg [7:0] phv_data_85; // @[matcher.scala 67:26]
  reg [7:0] phv_data_86; // @[matcher.scala 67:26]
  reg [7:0] phv_data_87; // @[matcher.scala 67:26]
  reg [7:0] phv_data_88; // @[matcher.scala 67:26]
  reg [7:0] phv_data_89; // @[matcher.scala 67:26]
  reg [7:0] phv_data_90; // @[matcher.scala 67:26]
  reg [7:0] phv_data_91; // @[matcher.scala 67:26]
  reg [7:0] phv_data_92; // @[matcher.scala 67:26]
  reg [7:0] phv_data_93; // @[matcher.scala 67:26]
  reg [7:0] phv_data_94; // @[matcher.scala 67:26]
  reg [7:0] phv_data_95; // @[matcher.scala 67:26]
  reg [7:0] phv_data_96; // @[matcher.scala 67:26]
  reg [7:0] phv_data_97; // @[matcher.scala 67:26]
  reg [7:0] phv_data_98; // @[matcher.scala 67:26]
  reg [7:0] phv_data_99; // @[matcher.scala 67:26]
  reg [7:0] phv_data_100; // @[matcher.scala 67:26]
  reg [7:0] phv_data_101; // @[matcher.scala 67:26]
  reg [7:0] phv_data_102; // @[matcher.scala 67:26]
  reg [7:0] phv_data_103; // @[matcher.scala 67:26]
  reg [7:0] phv_data_104; // @[matcher.scala 67:26]
  reg [7:0] phv_data_105; // @[matcher.scala 67:26]
  reg [7:0] phv_data_106; // @[matcher.scala 67:26]
  reg [7:0] phv_data_107; // @[matcher.scala 67:26]
  reg [7:0] phv_data_108; // @[matcher.scala 67:26]
  reg [7:0] phv_data_109; // @[matcher.scala 67:26]
  reg [7:0] phv_data_110; // @[matcher.scala 67:26]
  reg [7:0] phv_data_111; // @[matcher.scala 67:26]
  reg [7:0] phv_data_112; // @[matcher.scala 67:26]
  reg [7:0] phv_data_113; // @[matcher.scala 67:26]
  reg [7:0] phv_data_114; // @[matcher.scala 67:26]
  reg [7:0] phv_data_115; // @[matcher.scala 67:26]
  reg [7:0] phv_data_116; // @[matcher.scala 67:26]
  reg [7:0] phv_data_117; // @[matcher.scala 67:26]
  reg [7:0] phv_data_118; // @[matcher.scala 67:26]
  reg [7:0] phv_data_119; // @[matcher.scala 67:26]
  reg [7:0] phv_data_120; // @[matcher.scala 67:26]
  reg [7:0] phv_data_121; // @[matcher.scala 67:26]
  reg [7:0] phv_data_122; // @[matcher.scala 67:26]
  reg [7:0] phv_data_123; // @[matcher.scala 67:26]
  reg [7:0] phv_data_124; // @[matcher.scala 67:26]
  reg [7:0] phv_data_125; // @[matcher.scala 67:26]
  reg [7:0] phv_data_126; // @[matcher.scala 67:26]
  reg [7:0] phv_data_127; // @[matcher.scala 67:26]
  reg [7:0] phv_data_128; // @[matcher.scala 67:26]
  reg [7:0] phv_data_129; // @[matcher.scala 67:26]
  reg [7:0] phv_data_130; // @[matcher.scala 67:26]
  reg [7:0] phv_data_131; // @[matcher.scala 67:26]
  reg [7:0] phv_data_132; // @[matcher.scala 67:26]
  reg [7:0] phv_data_133; // @[matcher.scala 67:26]
  reg [7:0] phv_data_134; // @[matcher.scala 67:26]
  reg [7:0] phv_data_135; // @[matcher.scala 67:26]
  reg [7:0] phv_data_136; // @[matcher.scala 67:26]
  reg [7:0] phv_data_137; // @[matcher.scala 67:26]
  reg [7:0] phv_data_138; // @[matcher.scala 67:26]
  reg [7:0] phv_data_139; // @[matcher.scala 67:26]
  reg [7:0] phv_data_140; // @[matcher.scala 67:26]
  reg [7:0] phv_data_141; // @[matcher.scala 67:26]
  reg [7:0] phv_data_142; // @[matcher.scala 67:26]
  reg [7:0] phv_data_143; // @[matcher.scala 67:26]
  reg [7:0] phv_data_144; // @[matcher.scala 67:26]
  reg [7:0] phv_data_145; // @[matcher.scala 67:26]
  reg [7:0] phv_data_146; // @[matcher.scala 67:26]
  reg [7:0] phv_data_147; // @[matcher.scala 67:26]
  reg [7:0] phv_data_148; // @[matcher.scala 67:26]
  reg [7:0] phv_data_149; // @[matcher.scala 67:26]
  reg [7:0] phv_data_150; // @[matcher.scala 67:26]
  reg [7:0] phv_data_151; // @[matcher.scala 67:26]
  reg [7:0] phv_data_152; // @[matcher.scala 67:26]
  reg [7:0] phv_data_153; // @[matcher.scala 67:26]
  reg [7:0] phv_data_154; // @[matcher.scala 67:26]
  reg [7:0] phv_data_155; // @[matcher.scala 67:26]
  reg [7:0] phv_data_156; // @[matcher.scala 67:26]
  reg [7:0] phv_data_157; // @[matcher.scala 67:26]
  reg [7:0] phv_data_158; // @[matcher.scala 67:26]
  reg [7:0] phv_data_159; // @[matcher.scala 67:26]
  reg [7:0] phv_data_160; // @[matcher.scala 67:26]
  reg [7:0] phv_data_161; // @[matcher.scala 67:26]
  reg [7:0] phv_data_162; // @[matcher.scala 67:26]
  reg [7:0] phv_data_163; // @[matcher.scala 67:26]
  reg [7:0] phv_data_164; // @[matcher.scala 67:26]
  reg [7:0] phv_data_165; // @[matcher.scala 67:26]
  reg [7:0] phv_data_166; // @[matcher.scala 67:26]
  reg [7:0] phv_data_167; // @[matcher.scala 67:26]
  reg [7:0] phv_data_168; // @[matcher.scala 67:26]
  reg [7:0] phv_data_169; // @[matcher.scala 67:26]
  reg [7:0] phv_data_170; // @[matcher.scala 67:26]
  reg [7:0] phv_data_171; // @[matcher.scala 67:26]
  reg [7:0] phv_data_172; // @[matcher.scala 67:26]
  reg [7:0] phv_data_173; // @[matcher.scala 67:26]
  reg [7:0] phv_data_174; // @[matcher.scala 67:26]
  reg [7:0] phv_data_175; // @[matcher.scala 67:26]
  reg [7:0] phv_data_176; // @[matcher.scala 67:26]
  reg [7:0] phv_data_177; // @[matcher.scala 67:26]
  reg [7:0] phv_data_178; // @[matcher.scala 67:26]
  reg [7:0] phv_data_179; // @[matcher.scala 67:26]
  reg [7:0] phv_data_180; // @[matcher.scala 67:26]
  reg [7:0] phv_data_181; // @[matcher.scala 67:26]
  reg [7:0] phv_data_182; // @[matcher.scala 67:26]
  reg [7:0] phv_data_183; // @[matcher.scala 67:26]
  reg [7:0] phv_data_184; // @[matcher.scala 67:26]
  reg [7:0] phv_data_185; // @[matcher.scala 67:26]
  reg [7:0] phv_data_186; // @[matcher.scala 67:26]
  reg [7:0] phv_data_187; // @[matcher.scala 67:26]
  reg [7:0] phv_data_188; // @[matcher.scala 67:26]
  reg [7:0] phv_data_189; // @[matcher.scala 67:26]
  reg [7:0] phv_data_190; // @[matcher.scala 67:26]
  reg [7:0] phv_data_191; // @[matcher.scala 67:26]
  reg [7:0] phv_data_192; // @[matcher.scala 67:26]
  reg [7:0] phv_data_193; // @[matcher.scala 67:26]
  reg [7:0] phv_data_194; // @[matcher.scala 67:26]
  reg [7:0] phv_data_195; // @[matcher.scala 67:26]
  reg [7:0] phv_data_196; // @[matcher.scala 67:26]
  reg [7:0] phv_data_197; // @[matcher.scala 67:26]
  reg [7:0] phv_data_198; // @[matcher.scala 67:26]
  reg [7:0] phv_data_199; // @[matcher.scala 67:26]
  reg [7:0] phv_data_200; // @[matcher.scala 67:26]
  reg [7:0] phv_data_201; // @[matcher.scala 67:26]
  reg [7:0] phv_data_202; // @[matcher.scala 67:26]
  reg [7:0] phv_data_203; // @[matcher.scala 67:26]
  reg [7:0] phv_data_204; // @[matcher.scala 67:26]
  reg [7:0] phv_data_205; // @[matcher.scala 67:26]
  reg [7:0] phv_data_206; // @[matcher.scala 67:26]
  reg [7:0] phv_data_207; // @[matcher.scala 67:26]
  reg [7:0] phv_data_208; // @[matcher.scala 67:26]
  reg [7:0] phv_data_209; // @[matcher.scala 67:26]
  reg [7:0] phv_data_210; // @[matcher.scala 67:26]
  reg [7:0] phv_data_211; // @[matcher.scala 67:26]
  reg [7:0] phv_data_212; // @[matcher.scala 67:26]
  reg [7:0] phv_data_213; // @[matcher.scala 67:26]
  reg [7:0] phv_data_214; // @[matcher.scala 67:26]
  reg [7:0] phv_data_215; // @[matcher.scala 67:26]
  reg [7:0] phv_data_216; // @[matcher.scala 67:26]
  reg [7:0] phv_data_217; // @[matcher.scala 67:26]
  reg [7:0] phv_data_218; // @[matcher.scala 67:26]
  reg [7:0] phv_data_219; // @[matcher.scala 67:26]
  reg [7:0] phv_data_220; // @[matcher.scala 67:26]
  reg [7:0] phv_data_221; // @[matcher.scala 67:26]
  reg [7:0] phv_data_222; // @[matcher.scala 67:26]
  reg [7:0] phv_data_223; // @[matcher.scala 67:26]
  reg [7:0] phv_data_224; // @[matcher.scala 67:26]
  reg [7:0] phv_data_225; // @[matcher.scala 67:26]
  reg [7:0] phv_data_226; // @[matcher.scala 67:26]
  reg [7:0] phv_data_227; // @[matcher.scala 67:26]
  reg [7:0] phv_data_228; // @[matcher.scala 67:26]
  reg [7:0] phv_data_229; // @[matcher.scala 67:26]
  reg [7:0] phv_data_230; // @[matcher.scala 67:26]
  reg [7:0] phv_data_231; // @[matcher.scala 67:26]
  reg [7:0] phv_data_232; // @[matcher.scala 67:26]
  reg [7:0] phv_data_233; // @[matcher.scala 67:26]
  reg [7:0] phv_data_234; // @[matcher.scala 67:26]
  reg [7:0] phv_data_235; // @[matcher.scala 67:26]
  reg [7:0] phv_data_236; // @[matcher.scala 67:26]
  reg [7:0] phv_data_237; // @[matcher.scala 67:26]
  reg [7:0] phv_data_238; // @[matcher.scala 67:26]
  reg [7:0] phv_data_239; // @[matcher.scala 67:26]
  reg [7:0] phv_data_240; // @[matcher.scala 67:26]
  reg [7:0] phv_data_241; // @[matcher.scala 67:26]
  reg [7:0] phv_data_242; // @[matcher.scala 67:26]
  reg [7:0] phv_data_243; // @[matcher.scala 67:26]
  reg [7:0] phv_data_244; // @[matcher.scala 67:26]
  reg [7:0] phv_data_245; // @[matcher.scala 67:26]
  reg [7:0] phv_data_246; // @[matcher.scala 67:26]
  reg [7:0] phv_data_247; // @[matcher.scala 67:26]
  reg [7:0] phv_data_248; // @[matcher.scala 67:26]
  reg [7:0] phv_data_249; // @[matcher.scala 67:26]
  reg [7:0] phv_data_250; // @[matcher.scala 67:26]
  reg [7:0] phv_data_251; // @[matcher.scala 67:26]
  reg [7:0] phv_data_252; // @[matcher.scala 67:26]
  reg [7:0] phv_data_253; // @[matcher.scala 67:26]
  reg [7:0] phv_data_254; // @[matcher.scala 67:26]
  reg [7:0] phv_data_255; // @[matcher.scala 67:26]
  reg [15:0] phv_header_0; // @[matcher.scala 67:26]
  reg [15:0] phv_header_1; // @[matcher.scala 67:26]
  reg [15:0] phv_header_2; // @[matcher.scala 67:26]
  reg [15:0] phv_header_3; // @[matcher.scala 67:26]
  reg [15:0] phv_header_4; // @[matcher.scala 67:26]
  reg [15:0] phv_header_5; // @[matcher.scala 67:26]
  reg [15:0] phv_header_6; // @[matcher.scala 67:26]
  reg [15:0] phv_header_7; // @[matcher.scala 67:26]
  reg [15:0] phv_header_8; // @[matcher.scala 67:26]
  reg [15:0] phv_header_9; // @[matcher.scala 67:26]
  reg [15:0] phv_header_10; // @[matcher.scala 67:26]
  reg [15:0] phv_header_11; // @[matcher.scala 67:26]
  reg [15:0] phv_header_12; // @[matcher.scala 67:26]
  reg [15:0] phv_header_13; // @[matcher.scala 67:26]
  reg [15:0] phv_header_14; // @[matcher.scala 67:26]
  reg [15:0] phv_header_15; // @[matcher.scala 67:26]
  reg  phv_next_config_id; // @[matcher.scala 67:26]
  reg  phv_is_valid_processor; // @[matcher.scala 67:26]
  reg [7:0] key_offset; // @[matcher.scala 71:33]
  wire [5:0] read_key_offset_hi = key_offset[7:2]; // @[matcher.scala 73:49]
  wire [7:0] read_key_offset = {read_key_offset_hi,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 84:85 matcher.scala 84:85]
  wire [7:0] end_offset = _GEN_6 + key_offset; // @[matcher.scala 84:85]
  wire [8:0] _local_offset_T = {{1'd0}, read_key_offset}; // @[matcher.scala 87:77]
  wire [7:0] local_offset = _local_offset_T[7:0]; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_0_hi = local_offset[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_0_T = {match_key_qbytes_0_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_0_T_1 = {match_key_qbytes_0_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_0_T_2 = {match_key_qbytes_0_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_9 = 8'h1 == _match_key_qbytes_0_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10 = 8'h2 == _match_key_qbytes_0_T_2 ? phv_data_2 : _GEN_9; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11 = 8'h3 == _match_key_qbytes_0_T_2 ? phv_data_3 : _GEN_10; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12 = 8'h4 == _match_key_qbytes_0_T_2 ? phv_data_4 : _GEN_11; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_13 = 8'h5 == _match_key_qbytes_0_T_2 ? phv_data_5 : _GEN_12; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_14 = 8'h6 == _match_key_qbytes_0_T_2 ? phv_data_6 : _GEN_13; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_15 = 8'h7 == _match_key_qbytes_0_T_2 ? phv_data_7 : _GEN_14; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_16 = 8'h8 == _match_key_qbytes_0_T_2 ? phv_data_8 : _GEN_15; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_17 = 8'h9 == _match_key_qbytes_0_T_2 ? phv_data_9 : _GEN_16; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_18 = 8'ha == _match_key_qbytes_0_T_2 ? phv_data_10 : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_19 = 8'hb == _match_key_qbytes_0_T_2 ? phv_data_11 : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_20 = 8'hc == _match_key_qbytes_0_T_2 ? phv_data_12 : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_21 = 8'hd == _match_key_qbytes_0_T_2 ? phv_data_13 : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_22 = 8'he == _match_key_qbytes_0_T_2 ? phv_data_14 : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_23 = 8'hf == _match_key_qbytes_0_T_2 ? phv_data_15 : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_24 = 8'h10 == _match_key_qbytes_0_T_2 ? phv_data_16 : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_25 = 8'h11 == _match_key_qbytes_0_T_2 ? phv_data_17 : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_26 = 8'h12 == _match_key_qbytes_0_T_2 ? phv_data_18 : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_27 = 8'h13 == _match_key_qbytes_0_T_2 ? phv_data_19 : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_28 = 8'h14 == _match_key_qbytes_0_T_2 ? phv_data_20 : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_29 = 8'h15 == _match_key_qbytes_0_T_2 ? phv_data_21 : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_30 = 8'h16 == _match_key_qbytes_0_T_2 ? phv_data_22 : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_31 = 8'h17 == _match_key_qbytes_0_T_2 ? phv_data_23 : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_32 = 8'h18 == _match_key_qbytes_0_T_2 ? phv_data_24 : _GEN_31; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_33 = 8'h19 == _match_key_qbytes_0_T_2 ? phv_data_25 : _GEN_32; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_34 = 8'h1a == _match_key_qbytes_0_T_2 ? phv_data_26 : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_35 = 8'h1b == _match_key_qbytes_0_T_2 ? phv_data_27 : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_36 = 8'h1c == _match_key_qbytes_0_T_2 ? phv_data_28 : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_37 = 8'h1d == _match_key_qbytes_0_T_2 ? phv_data_29 : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_38 = 8'h1e == _match_key_qbytes_0_T_2 ? phv_data_30 : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_39 = 8'h1f == _match_key_qbytes_0_T_2 ? phv_data_31 : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_40 = 8'h20 == _match_key_qbytes_0_T_2 ? phv_data_32 : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_41 = 8'h21 == _match_key_qbytes_0_T_2 ? phv_data_33 : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_42 = 8'h22 == _match_key_qbytes_0_T_2 ? phv_data_34 : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_43 = 8'h23 == _match_key_qbytes_0_T_2 ? phv_data_35 : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_44 = 8'h24 == _match_key_qbytes_0_T_2 ? phv_data_36 : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_45 = 8'h25 == _match_key_qbytes_0_T_2 ? phv_data_37 : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_46 = 8'h26 == _match_key_qbytes_0_T_2 ? phv_data_38 : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_47 = 8'h27 == _match_key_qbytes_0_T_2 ? phv_data_39 : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_48 = 8'h28 == _match_key_qbytes_0_T_2 ? phv_data_40 : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_49 = 8'h29 == _match_key_qbytes_0_T_2 ? phv_data_41 : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_50 = 8'h2a == _match_key_qbytes_0_T_2 ? phv_data_42 : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 8'h2b == _match_key_qbytes_0_T_2 ? phv_data_43 : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 8'h2c == _match_key_qbytes_0_T_2 ? phv_data_44 : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 8'h2d == _match_key_qbytes_0_T_2 ? phv_data_45 : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 8'h2e == _match_key_qbytes_0_T_2 ? phv_data_46 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 8'h2f == _match_key_qbytes_0_T_2 ? phv_data_47 : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 8'h30 == _match_key_qbytes_0_T_2 ? phv_data_48 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 8'h31 == _match_key_qbytes_0_T_2 ? phv_data_49 : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 8'h32 == _match_key_qbytes_0_T_2 ? phv_data_50 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 8'h33 == _match_key_qbytes_0_T_2 ? phv_data_51 : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 8'h34 == _match_key_qbytes_0_T_2 ? phv_data_52 : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 8'h35 == _match_key_qbytes_0_T_2 ? phv_data_53 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 8'h36 == _match_key_qbytes_0_T_2 ? phv_data_54 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 8'h37 == _match_key_qbytes_0_T_2 ? phv_data_55 : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_64 = 8'h38 == _match_key_qbytes_0_T_2 ? phv_data_56 : _GEN_63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_65 = 8'h39 == _match_key_qbytes_0_T_2 ? phv_data_57 : _GEN_64; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_66 = 8'h3a == _match_key_qbytes_0_T_2 ? phv_data_58 : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_67 = 8'h3b == _match_key_qbytes_0_T_2 ? phv_data_59 : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_68 = 8'h3c == _match_key_qbytes_0_T_2 ? phv_data_60 : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_69 = 8'h3d == _match_key_qbytes_0_T_2 ? phv_data_61 : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_70 = 8'h3e == _match_key_qbytes_0_T_2 ? phv_data_62 : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_71 = 8'h3f == _match_key_qbytes_0_T_2 ? phv_data_63 : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_72 = 8'h40 == _match_key_qbytes_0_T_2 ? phv_data_64 : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_73 = 8'h41 == _match_key_qbytes_0_T_2 ? phv_data_65 : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_74 = 8'h42 == _match_key_qbytes_0_T_2 ? phv_data_66 : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_75 = 8'h43 == _match_key_qbytes_0_T_2 ? phv_data_67 : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_76 = 8'h44 == _match_key_qbytes_0_T_2 ? phv_data_68 : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_77 = 8'h45 == _match_key_qbytes_0_T_2 ? phv_data_69 : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_78 = 8'h46 == _match_key_qbytes_0_T_2 ? phv_data_70 : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_79 = 8'h47 == _match_key_qbytes_0_T_2 ? phv_data_71 : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_80 = 8'h48 == _match_key_qbytes_0_T_2 ? phv_data_72 : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_81 = 8'h49 == _match_key_qbytes_0_T_2 ? phv_data_73 : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_82 = 8'h4a == _match_key_qbytes_0_T_2 ? phv_data_74 : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_83 = 8'h4b == _match_key_qbytes_0_T_2 ? phv_data_75 : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_84 = 8'h4c == _match_key_qbytes_0_T_2 ? phv_data_76 : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_85 = 8'h4d == _match_key_qbytes_0_T_2 ? phv_data_77 : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_86 = 8'h4e == _match_key_qbytes_0_T_2 ? phv_data_78 : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_87 = 8'h4f == _match_key_qbytes_0_T_2 ? phv_data_79 : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_88 = 8'h50 == _match_key_qbytes_0_T_2 ? phv_data_80 : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_89 = 8'h51 == _match_key_qbytes_0_T_2 ? phv_data_81 : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_90 = 8'h52 == _match_key_qbytes_0_T_2 ? phv_data_82 : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_91 = 8'h53 == _match_key_qbytes_0_T_2 ? phv_data_83 : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_92 = 8'h54 == _match_key_qbytes_0_T_2 ? phv_data_84 : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_93 = 8'h55 == _match_key_qbytes_0_T_2 ? phv_data_85 : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_94 = 8'h56 == _match_key_qbytes_0_T_2 ? phv_data_86 : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_95 = 8'h57 == _match_key_qbytes_0_T_2 ? phv_data_87 : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_96 = 8'h58 == _match_key_qbytes_0_T_2 ? phv_data_88 : _GEN_95; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_97 = 8'h59 == _match_key_qbytes_0_T_2 ? phv_data_89 : _GEN_96; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_98 = 8'h5a == _match_key_qbytes_0_T_2 ? phv_data_90 : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_99 = 8'h5b == _match_key_qbytes_0_T_2 ? phv_data_91 : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_100 = 8'h5c == _match_key_qbytes_0_T_2 ? phv_data_92 : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_101 = 8'h5d == _match_key_qbytes_0_T_2 ? phv_data_93 : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_102 = 8'h5e == _match_key_qbytes_0_T_2 ? phv_data_94 : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_103 = 8'h5f == _match_key_qbytes_0_T_2 ? phv_data_95 : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_104 = 8'h60 == _match_key_qbytes_0_T_2 ? phv_data_96 : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_105 = 8'h61 == _match_key_qbytes_0_T_2 ? phv_data_97 : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_106 = 8'h62 == _match_key_qbytes_0_T_2 ? phv_data_98 : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_107 = 8'h63 == _match_key_qbytes_0_T_2 ? phv_data_99 : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_108 = 8'h64 == _match_key_qbytes_0_T_2 ? phv_data_100 : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_109 = 8'h65 == _match_key_qbytes_0_T_2 ? phv_data_101 : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_110 = 8'h66 == _match_key_qbytes_0_T_2 ? phv_data_102 : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_111 = 8'h67 == _match_key_qbytes_0_T_2 ? phv_data_103 : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_112 = 8'h68 == _match_key_qbytes_0_T_2 ? phv_data_104 : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_113 = 8'h69 == _match_key_qbytes_0_T_2 ? phv_data_105 : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_114 = 8'h6a == _match_key_qbytes_0_T_2 ? phv_data_106 : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_115 = 8'h6b == _match_key_qbytes_0_T_2 ? phv_data_107 : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_116 = 8'h6c == _match_key_qbytes_0_T_2 ? phv_data_108 : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_117 = 8'h6d == _match_key_qbytes_0_T_2 ? phv_data_109 : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_118 = 8'h6e == _match_key_qbytes_0_T_2 ? phv_data_110 : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_119 = 8'h6f == _match_key_qbytes_0_T_2 ? phv_data_111 : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_120 = 8'h70 == _match_key_qbytes_0_T_2 ? phv_data_112 : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_121 = 8'h71 == _match_key_qbytes_0_T_2 ? phv_data_113 : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_122 = 8'h72 == _match_key_qbytes_0_T_2 ? phv_data_114 : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_123 = 8'h73 == _match_key_qbytes_0_T_2 ? phv_data_115 : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_124 = 8'h74 == _match_key_qbytes_0_T_2 ? phv_data_116 : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_125 = 8'h75 == _match_key_qbytes_0_T_2 ? phv_data_117 : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_126 = 8'h76 == _match_key_qbytes_0_T_2 ? phv_data_118 : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_127 = 8'h77 == _match_key_qbytes_0_T_2 ? phv_data_119 : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_128 = 8'h78 == _match_key_qbytes_0_T_2 ? phv_data_120 : _GEN_127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_129 = 8'h79 == _match_key_qbytes_0_T_2 ? phv_data_121 : _GEN_128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_130 = 8'h7a == _match_key_qbytes_0_T_2 ? phv_data_122 : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_131 = 8'h7b == _match_key_qbytes_0_T_2 ? phv_data_123 : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_132 = 8'h7c == _match_key_qbytes_0_T_2 ? phv_data_124 : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_133 = 8'h7d == _match_key_qbytes_0_T_2 ? phv_data_125 : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_134 = 8'h7e == _match_key_qbytes_0_T_2 ? phv_data_126 : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_135 = 8'h7f == _match_key_qbytes_0_T_2 ? phv_data_127 : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_136 = 8'h80 == _match_key_qbytes_0_T_2 ? phv_data_128 : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_137 = 8'h81 == _match_key_qbytes_0_T_2 ? phv_data_129 : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_138 = 8'h82 == _match_key_qbytes_0_T_2 ? phv_data_130 : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_139 = 8'h83 == _match_key_qbytes_0_T_2 ? phv_data_131 : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_140 = 8'h84 == _match_key_qbytes_0_T_2 ? phv_data_132 : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_141 = 8'h85 == _match_key_qbytes_0_T_2 ? phv_data_133 : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_142 = 8'h86 == _match_key_qbytes_0_T_2 ? phv_data_134 : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_143 = 8'h87 == _match_key_qbytes_0_T_2 ? phv_data_135 : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_144 = 8'h88 == _match_key_qbytes_0_T_2 ? phv_data_136 : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_145 = 8'h89 == _match_key_qbytes_0_T_2 ? phv_data_137 : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_146 = 8'h8a == _match_key_qbytes_0_T_2 ? phv_data_138 : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_147 = 8'h8b == _match_key_qbytes_0_T_2 ? phv_data_139 : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_148 = 8'h8c == _match_key_qbytes_0_T_2 ? phv_data_140 : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_149 = 8'h8d == _match_key_qbytes_0_T_2 ? phv_data_141 : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_150 = 8'h8e == _match_key_qbytes_0_T_2 ? phv_data_142 : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_151 = 8'h8f == _match_key_qbytes_0_T_2 ? phv_data_143 : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_152 = 8'h90 == _match_key_qbytes_0_T_2 ? phv_data_144 : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_153 = 8'h91 == _match_key_qbytes_0_T_2 ? phv_data_145 : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_154 = 8'h92 == _match_key_qbytes_0_T_2 ? phv_data_146 : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_155 = 8'h93 == _match_key_qbytes_0_T_2 ? phv_data_147 : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_156 = 8'h94 == _match_key_qbytes_0_T_2 ? phv_data_148 : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_157 = 8'h95 == _match_key_qbytes_0_T_2 ? phv_data_149 : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_158 = 8'h96 == _match_key_qbytes_0_T_2 ? phv_data_150 : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_159 = 8'h97 == _match_key_qbytes_0_T_2 ? phv_data_151 : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_160 = 8'h98 == _match_key_qbytes_0_T_2 ? phv_data_152 : _GEN_159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_161 = 8'h99 == _match_key_qbytes_0_T_2 ? phv_data_153 : _GEN_160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_162 = 8'h9a == _match_key_qbytes_0_T_2 ? phv_data_154 : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_163 = 8'h9b == _match_key_qbytes_0_T_2 ? phv_data_155 : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_164 = 8'h9c == _match_key_qbytes_0_T_2 ? phv_data_156 : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_165 = 8'h9d == _match_key_qbytes_0_T_2 ? phv_data_157 : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_166 = 8'h9e == _match_key_qbytes_0_T_2 ? phv_data_158 : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_167 = 8'h9f == _match_key_qbytes_0_T_2 ? phv_data_159 : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_168 = 8'ha0 == _match_key_qbytes_0_T_2 ? phv_data_160 : _GEN_167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_169 = 8'ha1 == _match_key_qbytes_0_T_2 ? phv_data_161 : _GEN_168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_170 = 8'ha2 == _match_key_qbytes_0_T_2 ? phv_data_162 : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_171 = 8'ha3 == _match_key_qbytes_0_T_2 ? phv_data_163 : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_172 = 8'ha4 == _match_key_qbytes_0_T_2 ? phv_data_164 : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_173 = 8'ha5 == _match_key_qbytes_0_T_2 ? phv_data_165 : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_174 = 8'ha6 == _match_key_qbytes_0_T_2 ? phv_data_166 : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_175 = 8'ha7 == _match_key_qbytes_0_T_2 ? phv_data_167 : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_176 = 8'ha8 == _match_key_qbytes_0_T_2 ? phv_data_168 : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_177 = 8'ha9 == _match_key_qbytes_0_T_2 ? phv_data_169 : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_178 = 8'haa == _match_key_qbytes_0_T_2 ? phv_data_170 : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_179 = 8'hab == _match_key_qbytes_0_T_2 ? phv_data_171 : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_180 = 8'hac == _match_key_qbytes_0_T_2 ? phv_data_172 : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_181 = 8'had == _match_key_qbytes_0_T_2 ? phv_data_173 : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_182 = 8'hae == _match_key_qbytes_0_T_2 ? phv_data_174 : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_183 = 8'haf == _match_key_qbytes_0_T_2 ? phv_data_175 : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_184 = 8'hb0 == _match_key_qbytes_0_T_2 ? phv_data_176 : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_185 = 8'hb1 == _match_key_qbytes_0_T_2 ? phv_data_177 : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_186 = 8'hb2 == _match_key_qbytes_0_T_2 ? phv_data_178 : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_187 = 8'hb3 == _match_key_qbytes_0_T_2 ? phv_data_179 : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_188 = 8'hb4 == _match_key_qbytes_0_T_2 ? phv_data_180 : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_189 = 8'hb5 == _match_key_qbytes_0_T_2 ? phv_data_181 : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_190 = 8'hb6 == _match_key_qbytes_0_T_2 ? phv_data_182 : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_191 = 8'hb7 == _match_key_qbytes_0_T_2 ? phv_data_183 : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_192 = 8'hb8 == _match_key_qbytes_0_T_2 ? phv_data_184 : _GEN_191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_193 = 8'hb9 == _match_key_qbytes_0_T_2 ? phv_data_185 : _GEN_192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_194 = 8'hba == _match_key_qbytes_0_T_2 ? phv_data_186 : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_195 = 8'hbb == _match_key_qbytes_0_T_2 ? phv_data_187 : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_196 = 8'hbc == _match_key_qbytes_0_T_2 ? phv_data_188 : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_197 = 8'hbd == _match_key_qbytes_0_T_2 ? phv_data_189 : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_198 = 8'hbe == _match_key_qbytes_0_T_2 ? phv_data_190 : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_199 = 8'hbf == _match_key_qbytes_0_T_2 ? phv_data_191 : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_200 = 8'hc0 == _match_key_qbytes_0_T_2 ? phv_data_192 : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_201 = 8'hc1 == _match_key_qbytes_0_T_2 ? phv_data_193 : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_202 = 8'hc2 == _match_key_qbytes_0_T_2 ? phv_data_194 : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_203 = 8'hc3 == _match_key_qbytes_0_T_2 ? phv_data_195 : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_204 = 8'hc4 == _match_key_qbytes_0_T_2 ? phv_data_196 : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_205 = 8'hc5 == _match_key_qbytes_0_T_2 ? phv_data_197 : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_206 = 8'hc6 == _match_key_qbytes_0_T_2 ? phv_data_198 : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_207 = 8'hc7 == _match_key_qbytes_0_T_2 ? phv_data_199 : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_208 = 8'hc8 == _match_key_qbytes_0_T_2 ? phv_data_200 : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_209 = 8'hc9 == _match_key_qbytes_0_T_2 ? phv_data_201 : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_210 = 8'hca == _match_key_qbytes_0_T_2 ? phv_data_202 : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_211 = 8'hcb == _match_key_qbytes_0_T_2 ? phv_data_203 : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_212 = 8'hcc == _match_key_qbytes_0_T_2 ? phv_data_204 : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_213 = 8'hcd == _match_key_qbytes_0_T_2 ? phv_data_205 : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_214 = 8'hce == _match_key_qbytes_0_T_2 ? phv_data_206 : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_215 = 8'hcf == _match_key_qbytes_0_T_2 ? phv_data_207 : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_216 = 8'hd0 == _match_key_qbytes_0_T_2 ? phv_data_208 : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_217 = 8'hd1 == _match_key_qbytes_0_T_2 ? phv_data_209 : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_218 = 8'hd2 == _match_key_qbytes_0_T_2 ? phv_data_210 : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_219 = 8'hd3 == _match_key_qbytes_0_T_2 ? phv_data_211 : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_220 = 8'hd4 == _match_key_qbytes_0_T_2 ? phv_data_212 : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_221 = 8'hd5 == _match_key_qbytes_0_T_2 ? phv_data_213 : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_222 = 8'hd6 == _match_key_qbytes_0_T_2 ? phv_data_214 : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_223 = 8'hd7 == _match_key_qbytes_0_T_2 ? phv_data_215 : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_224 = 8'hd8 == _match_key_qbytes_0_T_2 ? phv_data_216 : _GEN_223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_225 = 8'hd9 == _match_key_qbytes_0_T_2 ? phv_data_217 : _GEN_224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_226 = 8'hda == _match_key_qbytes_0_T_2 ? phv_data_218 : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_227 = 8'hdb == _match_key_qbytes_0_T_2 ? phv_data_219 : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_228 = 8'hdc == _match_key_qbytes_0_T_2 ? phv_data_220 : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_229 = 8'hdd == _match_key_qbytes_0_T_2 ? phv_data_221 : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_230 = 8'hde == _match_key_qbytes_0_T_2 ? phv_data_222 : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_231 = 8'hdf == _match_key_qbytes_0_T_2 ? phv_data_223 : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_232 = 8'he0 == _match_key_qbytes_0_T_2 ? phv_data_224 : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_233 = 8'he1 == _match_key_qbytes_0_T_2 ? phv_data_225 : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_234 = 8'he2 == _match_key_qbytes_0_T_2 ? phv_data_226 : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_235 = 8'he3 == _match_key_qbytes_0_T_2 ? phv_data_227 : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_236 = 8'he4 == _match_key_qbytes_0_T_2 ? phv_data_228 : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_237 = 8'he5 == _match_key_qbytes_0_T_2 ? phv_data_229 : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_238 = 8'he6 == _match_key_qbytes_0_T_2 ? phv_data_230 : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_239 = 8'he7 == _match_key_qbytes_0_T_2 ? phv_data_231 : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_240 = 8'he8 == _match_key_qbytes_0_T_2 ? phv_data_232 : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_241 = 8'he9 == _match_key_qbytes_0_T_2 ? phv_data_233 : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_242 = 8'hea == _match_key_qbytes_0_T_2 ? phv_data_234 : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_243 = 8'heb == _match_key_qbytes_0_T_2 ? phv_data_235 : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_244 = 8'hec == _match_key_qbytes_0_T_2 ? phv_data_236 : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_245 = 8'hed == _match_key_qbytes_0_T_2 ? phv_data_237 : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_246 = 8'hee == _match_key_qbytes_0_T_2 ? phv_data_238 : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_247 = 8'hef == _match_key_qbytes_0_T_2 ? phv_data_239 : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_248 = 8'hf0 == _match_key_qbytes_0_T_2 ? phv_data_240 : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_249 = 8'hf1 == _match_key_qbytes_0_T_2 ? phv_data_241 : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_250 = 8'hf2 == _match_key_qbytes_0_T_2 ? phv_data_242 : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_251 = 8'hf3 == _match_key_qbytes_0_T_2 ? phv_data_243 : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_252 = 8'hf4 == _match_key_qbytes_0_T_2 ? phv_data_244 : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_253 = 8'hf5 == _match_key_qbytes_0_T_2 ? phv_data_245 : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_254 = 8'hf6 == _match_key_qbytes_0_T_2 ? phv_data_246 : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_255 = 8'hf7 == _match_key_qbytes_0_T_2 ? phv_data_247 : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_256 = 8'hf8 == _match_key_qbytes_0_T_2 ? phv_data_248 : _GEN_255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_257 = 8'hf9 == _match_key_qbytes_0_T_2 ? phv_data_249 : _GEN_256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_258 = 8'hfa == _match_key_qbytes_0_T_2 ? phv_data_250 : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_259 = 8'hfb == _match_key_qbytes_0_T_2 ? phv_data_251 : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_260 = 8'hfc == _match_key_qbytes_0_T_2 ? phv_data_252 : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_261 = 8'hfd == _match_key_qbytes_0_T_2 ? phv_data_253 : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_262 = 8'hfe == _match_key_qbytes_0_T_2 ? phv_data_254 : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_263 = 8'hff == _match_key_qbytes_0_T_2 ? phv_data_255 : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_265 = 8'h1 == local_offset ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_266 = 8'h2 == local_offset ? phv_data_2 : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_267 = 8'h3 == local_offset ? phv_data_3 : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_268 = 8'h4 == local_offset ? phv_data_4 : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_269 = 8'h5 == local_offset ? phv_data_5 : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_270 = 8'h6 == local_offset ? phv_data_6 : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_271 = 8'h7 == local_offset ? phv_data_7 : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_272 = 8'h8 == local_offset ? phv_data_8 : _GEN_271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_273 = 8'h9 == local_offset ? phv_data_9 : _GEN_272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_274 = 8'ha == local_offset ? phv_data_10 : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_275 = 8'hb == local_offset ? phv_data_11 : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_276 = 8'hc == local_offset ? phv_data_12 : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_277 = 8'hd == local_offset ? phv_data_13 : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_278 = 8'he == local_offset ? phv_data_14 : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_279 = 8'hf == local_offset ? phv_data_15 : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_280 = 8'h10 == local_offset ? phv_data_16 : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_281 = 8'h11 == local_offset ? phv_data_17 : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_282 = 8'h12 == local_offset ? phv_data_18 : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_283 = 8'h13 == local_offset ? phv_data_19 : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_284 = 8'h14 == local_offset ? phv_data_20 : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_285 = 8'h15 == local_offset ? phv_data_21 : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_286 = 8'h16 == local_offset ? phv_data_22 : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_287 = 8'h17 == local_offset ? phv_data_23 : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_288 = 8'h18 == local_offset ? phv_data_24 : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_289 = 8'h19 == local_offset ? phv_data_25 : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_290 = 8'h1a == local_offset ? phv_data_26 : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_291 = 8'h1b == local_offset ? phv_data_27 : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_292 = 8'h1c == local_offset ? phv_data_28 : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_293 = 8'h1d == local_offset ? phv_data_29 : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_294 = 8'h1e == local_offset ? phv_data_30 : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_295 = 8'h1f == local_offset ? phv_data_31 : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_296 = 8'h20 == local_offset ? phv_data_32 : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_297 = 8'h21 == local_offset ? phv_data_33 : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_298 = 8'h22 == local_offset ? phv_data_34 : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_299 = 8'h23 == local_offset ? phv_data_35 : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_300 = 8'h24 == local_offset ? phv_data_36 : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_301 = 8'h25 == local_offset ? phv_data_37 : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_302 = 8'h26 == local_offset ? phv_data_38 : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_303 = 8'h27 == local_offset ? phv_data_39 : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_304 = 8'h28 == local_offset ? phv_data_40 : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_305 = 8'h29 == local_offset ? phv_data_41 : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_306 = 8'h2a == local_offset ? phv_data_42 : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_307 = 8'h2b == local_offset ? phv_data_43 : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_308 = 8'h2c == local_offset ? phv_data_44 : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_309 = 8'h2d == local_offset ? phv_data_45 : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_310 = 8'h2e == local_offset ? phv_data_46 : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_311 = 8'h2f == local_offset ? phv_data_47 : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_312 = 8'h30 == local_offset ? phv_data_48 : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_313 = 8'h31 == local_offset ? phv_data_49 : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_314 = 8'h32 == local_offset ? phv_data_50 : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_315 = 8'h33 == local_offset ? phv_data_51 : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_316 = 8'h34 == local_offset ? phv_data_52 : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_317 = 8'h35 == local_offset ? phv_data_53 : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_318 = 8'h36 == local_offset ? phv_data_54 : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_319 = 8'h37 == local_offset ? phv_data_55 : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_320 = 8'h38 == local_offset ? phv_data_56 : _GEN_319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_321 = 8'h39 == local_offset ? phv_data_57 : _GEN_320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_322 = 8'h3a == local_offset ? phv_data_58 : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_323 = 8'h3b == local_offset ? phv_data_59 : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_324 = 8'h3c == local_offset ? phv_data_60 : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_325 = 8'h3d == local_offset ? phv_data_61 : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_326 = 8'h3e == local_offset ? phv_data_62 : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_327 = 8'h3f == local_offset ? phv_data_63 : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_328 = 8'h40 == local_offset ? phv_data_64 : _GEN_327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_329 = 8'h41 == local_offset ? phv_data_65 : _GEN_328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_330 = 8'h42 == local_offset ? phv_data_66 : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_331 = 8'h43 == local_offset ? phv_data_67 : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_332 = 8'h44 == local_offset ? phv_data_68 : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_333 = 8'h45 == local_offset ? phv_data_69 : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_334 = 8'h46 == local_offset ? phv_data_70 : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_335 = 8'h47 == local_offset ? phv_data_71 : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_336 = 8'h48 == local_offset ? phv_data_72 : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_337 = 8'h49 == local_offset ? phv_data_73 : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_338 = 8'h4a == local_offset ? phv_data_74 : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_339 = 8'h4b == local_offset ? phv_data_75 : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_340 = 8'h4c == local_offset ? phv_data_76 : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_341 = 8'h4d == local_offset ? phv_data_77 : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_342 = 8'h4e == local_offset ? phv_data_78 : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_343 = 8'h4f == local_offset ? phv_data_79 : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_344 = 8'h50 == local_offset ? phv_data_80 : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_345 = 8'h51 == local_offset ? phv_data_81 : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_346 = 8'h52 == local_offset ? phv_data_82 : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_347 = 8'h53 == local_offset ? phv_data_83 : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_348 = 8'h54 == local_offset ? phv_data_84 : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_349 = 8'h55 == local_offset ? phv_data_85 : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_350 = 8'h56 == local_offset ? phv_data_86 : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_351 = 8'h57 == local_offset ? phv_data_87 : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_352 = 8'h58 == local_offset ? phv_data_88 : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_353 = 8'h59 == local_offset ? phv_data_89 : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_354 = 8'h5a == local_offset ? phv_data_90 : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_355 = 8'h5b == local_offset ? phv_data_91 : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_356 = 8'h5c == local_offset ? phv_data_92 : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_357 = 8'h5d == local_offset ? phv_data_93 : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_358 = 8'h5e == local_offset ? phv_data_94 : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_359 = 8'h5f == local_offset ? phv_data_95 : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_360 = 8'h60 == local_offset ? phv_data_96 : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_361 = 8'h61 == local_offset ? phv_data_97 : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_362 = 8'h62 == local_offset ? phv_data_98 : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_363 = 8'h63 == local_offset ? phv_data_99 : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_364 = 8'h64 == local_offset ? phv_data_100 : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_365 = 8'h65 == local_offset ? phv_data_101 : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_366 = 8'h66 == local_offset ? phv_data_102 : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_367 = 8'h67 == local_offset ? phv_data_103 : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_368 = 8'h68 == local_offset ? phv_data_104 : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_369 = 8'h69 == local_offset ? phv_data_105 : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_370 = 8'h6a == local_offset ? phv_data_106 : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_371 = 8'h6b == local_offset ? phv_data_107 : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_372 = 8'h6c == local_offset ? phv_data_108 : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_373 = 8'h6d == local_offset ? phv_data_109 : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_374 = 8'h6e == local_offset ? phv_data_110 : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_375 = 8'h6f == local_offset ? phv_data_111 : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_376 = 8'h70 == local_offset ? phv_data_112 : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_377 = 8'h71 == local_offset ? phv_data_113 : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_378 = 8'h72 == local_offset ? phv_data_114 : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_379 = 8'h73 == local_offset ? phv_data_115 : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_380 = 8'h74 == local_offset ? phv_data_116 : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_381 = 8'h75 == local_offset ? phv_data_117 : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_382 = 8'h76 == local_offset ? phv_data_118 : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_383 = 8'h77 == local_offset ? phv_data_119 : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_384 = 8'h78 == local_offset ? phv_data_120 : _GEN_383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_385 = 8'h79 == local_offset ? phv_data_121 : _GEN_384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_386 = 8'h7a == local_offset ? phv_data_122 : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_387 = 8'h7b == local_offset ? phv_data_123 : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_388 = 8'h7c == local_offset ? phv_data_124 : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_389 = 8'h7d == local_offset ? phv_data_125 : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_390 = 8'h7e == local_offset ? phv_data_126 : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_391 = 8'h7f == local_offset ? phv_data_127 : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_392 = 8'h80 == local_offset ? phv_data_128 : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_393 = 8'h81 == local_offset ? phv_data_129 : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_394 = 8'h82 == local_offset ? phv_data_130 : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_395 = 8'h83 == local_offset ? phv_data_131 : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_396 = 8'h84 == local_offset ? phv_data_132 : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_397 = 8'h85 == local_offset ? phv_data_133 : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_398 = 8'h86 == local_offset ? phv_data_134 : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_399 = 8'h87 == local_offset ? phv_data_135 : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_400 = 8'h88 == local_offset ? phv_data_136 : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_401 = 8'h89 == local_offset ? phv_data_137 : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_402 = 8'h8a == local_offset ? phv_data_138 : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_403 = 8'h8b == local_offset ? phv_data_139 : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_404 = 8'h8c == local_offset ? phv_data_140 : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_405 = 8'h8d == local_offset ? phv_data_141 : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_406 = 8'h8e == local_offset ? phv_data_142 : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_407 = 8'h8f == local_offset ? phv_data_143 : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_408 = 8'h90 == local_offset ? phv_data_144 : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_409 = 8'h91 == local_offset ? phv_data_145 : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_410 = 8'h92 == local_offset ? phv_data_146 : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_411 = 8'h93 == local_offset ? phv_data_147 : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_412 = 8'h94 == local_offset ? phv_data_148 : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_413 = 8'h95 == local_offset ? phv_data_149 : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_414 = 8'h96 == local_offset ? phv_data_150 : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_415 = 8'h97 == local_offset ? phv_data_151 : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_416 = 8'h98 == local_offset ? phv_data_152 : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_417 = 8'h99 == local_offset ? phv_data_153 : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_418 = 8'h9a == local_offset ? phv_data_154 : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_419 = 8'h9b == local_offset ? phv_data_155 : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_420 = 8'h9c == local_offset ? phv_data_156 : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_421 = 8'h9d == local_offset ? phv_data_157 : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_422 = 8'h9e == local_offset ? phv_data_158 : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_423 = 8'h9f == local_offset ? phv_data_159 : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_424 = 8'ha0 == local_offset ? phv_data_160 : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_425 = 8'ha1 == local_offset ? phv_data_161 : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_426 = 8'ha2 == local_offset ? phv_data_162 : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_427 = 8'ha3 == local_offset ? phv_data_163 : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_428 = 8'ha4 == local_offset ? phv_data_164 : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_429 = 8'ha5 == local_offset ? phv_data_165 : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_430 = 8'ha6 == local_offset ? phv_data_166 : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_431 = 8'ha7 == local_offset ? phv_data_167 : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_432 = 8'ha8 == local_offset ? phv_data_168 : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_433 = 8'ha9 == local_offset ? phv_data_169 : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_434 = 8'haa == local_offset ? phv_data_170 : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_435 = 8'hab == local_offset ? phv_data_171 : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_436 = 8'hac == local_offset ? phv_data_172 : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_437 = 8'had == local_offset ? phv_data_173 : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_438 = 8'hae == local_offset ? phv_data_174 : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_439 = 8'haf == local_offset ? phv_data_175 : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_440 = 8'hb0 == local_offset ? phv_data_176 : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_441 = 8'hb1 == local_offset ? phv_data_177 : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_442 = 8'hb2 == local_offset ? phv_data_178 : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_443 = 8'hb3 == local_offset ? phv_data_179 : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_444 = 8'hb4 == local_offset ? phv_data_180 : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_445 = 8'hb5 == local_offset ? phv_data_181 : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_446 = 8'hb6 == local_offset ? phv_data_182 : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_447 = 8'hb7 == local_offset ? phv_data_183 : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_448 = 8'hb8 == local_offset ? phv_data_184 : _GEN_447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_449 = 8'hb9 == local_offset ? phv_data_185 : _GEN_448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_450 = 8'hba == local_offset ? phv_data_186 : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_451 = 8'hbb == local_offset ? phv_data_187 : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_452 = 8'hbc == local_offset ? phv_data_188 : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_453 = 8'hbd == local_offset ? phv_data_189 : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_454 = 8'hbe == local_offset ? phv_data_190 : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_455 = 8'hbf == local_offset ? phv_data_191 : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_456 = 8'hc0 == local_offset ? phv_data_192 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_457 = 8'hc1 == local_offset ? phv_data_193 : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_458 = 8'hc2 == local_offset ? phv_data_194 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_459 = 8'hc3 == local_offset ? phv_data_195 : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_460 = 8'hc4 == local_offset ? phv_data_196 : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_461 = 8'hc5 == local_offset ? phv_data_197 : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_462 = 8'hc6 == local_offset ? phv_data_198 : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_463 = 8'hc7 == local_offset ? phv_data_199 : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_464 = 8'hc8 == local_offset ? phv_data_200 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_465 = 8'hc9 == local_offset ? phv_data_201 : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_466 = 8'hca == local_offset ? phv_data_202 : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_467 = 8'hcb == local_offset ? phv_data_203 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_468 = 8'hcc == local_offset ? phv_data_204 : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_469 = 8'hcd == local_offset ? phv_data_205 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_470 = 8'hce == local_offset ? phv_data_206 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_471 = 8'hcf == local_offset ? phv_data_207 : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_472 = 8'hd0 == local_offset ? phv_data_208 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_473 = 8'hd1 == local_offset ? phv_data_209 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_474 = 8'hd2 == local_offset ? phv_data_210 : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_475 = 8'hd3 == local_offset ? phv_data_211 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_476 = 8'hd4 == local_offset ? phv_data_212 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_477 = 8'hd5 == local_offset ? phv_data_213 : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_478 = 8'hd6 == local_offset ? phv_data_214 : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_479 = 8'hd7 == local_offset ? phv_data_215 : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_480 = 8'hd8 == local_offset ? phv_data_216 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_481 = 8'hd9 == local_offset ? phv_data_217 : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_482 = 8'hda == local_offset ? phv_data_218 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_483 = 8'hdb == local_offset ? phv_data_219 : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_484 = 8'hdc == local_offset ? phv_data_220 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_485 = 8'hdd == local_offset ? phv_data_221 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_486 = 8'hde == local_offset ? phv_data_222 : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_487 = 8'hdf == local_offset ? phv_data_223 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_488 = 8'he0 == local_offset ? phv_data_224 : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_489 = 8'he1 == local_offset ? phv_data_225 : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_490 = 8'he2 == local_offset ? phv_data_226 : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_491 = 8'he3 == local_offset ? phv_data_227 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_492 = 8'he4 == local_offset ? phv_data_228 : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_493 = 8'he5 == local_offset ? phv_data_229 : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_494 = 8'he6 == local_offset ? phv_data_230 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_495 = 8'he7 == local_offset ? phv_data_231 : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_496 = 8'he8 == local_offset ? phv_data_232 : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_497 = 8'he9 == local_offset ? phv_data_233 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_498 = 8'hea == local_offset ? phv_data_234 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_499 = 8'heb == local_offset ? phv_data_235 : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_500 = 8'hec == local_offset ? phv_data_236 : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_501 = 8'hed == local_offset ? phv_data_237 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_502 = 8'hee == local_offset ? phv_data_238 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_503 = 8'hef == local_offset ? phv_data_239 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_504 = 8'hf0 == local_offset ? phv_data_240 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_505 = 8'hf1 == local_offset ? phv_data_241 : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_506 = 8'hf2 == local_offset ? phv_data_242 : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_507 = 8'hf3 == local_offset ? phv_data_243 : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_508 = 8'hf4 == local_offset ? phv_data_244 : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_509 = 8'hf5 == local_offset ? phv_data_245 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_510 = 8'hf6 == local_offset ? phv_data_246 : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_511 = 8'hf7 == local_offset ? phv_data_247 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_512 = 8'hf8 == local_offset ? phv_data_248 : _GEN_511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_513 = 8'hf9 == local_offset ? phv_data_249 : _GEN_512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_514 = 8'hfa == local_offset ? phv_data_250 : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_515 = 8'hfb == local_offset ? phv_data_251 : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_516 = 8'hfc == local_offset ? phv_data_252 : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_517 = 8'hfd == local_offset ? phv_data_253 : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_518 = 8'hfe == local_offset ? phv_data_254 : _GEN_517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_519 = 8'hff == local_offset ? phv_data_255 : _GEN_518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_521 = 8'h1 == _match_key_qbytes_0_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_522 = 8'h2 == _match_key_qbytes_0_T ? phv_data_2 : _GEN_521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_523 = 8'h3 == _match_key_qbytes_0_T ? phv_data_3 : _GEN_522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_524 = 8'h4 == _match_key_qbytes_0_T ? phv_data_4 : _GEN_523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_525 = 8'h5 == _match_key_qbytes_0_T ? phv_data_5 : _GEN_524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_526 = 8'h6 == _match_key_qbytes_0_T ? phv_data_6 : _GEN_525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_527 = 8'h7 == _match_key_qbytes_0_T ? phv_data_7 : _GEN_526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_528 = 8'h8 == _match_key_qbytes_0_T ? phv_data_8 : _GEN_527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_529 = 8'h9 == _match_key_qbytes_0_T ? phv_data_9 : _GEN_528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_530 = 8'ha == _match_key_qbytes_0_T ? phv_data_10 : _GEN_529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_531 = 8'hb == _match_key_qbytes_0_T ? phv_data_11 : _GEN_530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_532 = 8'hc == _match_key_qbytes_0_T ? phv_data_12 : _GEN_531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_533 = 8'hd == _match_key_qbytes_0_T ? phv_data_13 : _GEN_532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_534 = 8'he == _match_key_qbytes_0_T ? phv_data_14 : _GEN_533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_535 = 8'hf == _match_key_qbytes_0_T ? phv_data_15 : _GEN_534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_536 = 8'h10 == _match_key_qbytes_0_T ? phv_data_16 : _GEN_535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_537 = 8'h11 == _match_key_qbytes_0_T ? phv_data_17 : _GEN_536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_538 = 8'h12 == _match_key_qbytes_0_T ? phv_data_18 : _GEN_537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_539 = 8'h13 == _match_key_qbytes_0_T ? phv_data_19 : _GEN_538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_540 = 8'h14 == _match_key_qbytes_0_T ? phv_data_20 : _GEN_539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_541 = 8'h15 == _match_key_qbytes_0_T ? phv_data_21 : _GEN_540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_542 = 8'h16 == _match_key_qbytes_0_T ? phv_data_22 : _GEN_541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_543 = 8'h17 == _match_key_qbytes_0_T ? phv_data_23 : _GEN_542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_544 = 8'h18 == _match_key_qbytes_0_T ? phv_data_24 : _GEN_543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_545 = 8'h19 == _match_key_qbytes_0_T ? phv_data_25 : _GEN_544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_546 = 8'h1a == _match_key_qbytes_0_T ? phv_data_26 : _GEN_545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_547 = 8'h1b == _match_key_qbytes_0_T ? phv_data_27 : _GEN_546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_548 = 8'h1c == _match_key_qbytes_0_T ? phv_data_28 : _GEN_547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_549 = 8'h1d == _match_key_qbytes_0_T ? phv_data_29 : _GEN_548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_550 = 8'h1e == _match_key_qbytes_0_T ? phv_data_30 : _GEN_549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_551 = 8'h1f == _match_key_qbytes_0_T ? phv_data_31 : _GEN_550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_552 = 8'h20 == _match_key_qbytes_0_T ? phv_data_32 : _GEN_551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_553 = 8'h21 == _match_key_qbytes_0_T ? phv_data_33 : _GEN_552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_554 = 8'h22 == _match_key_qbytes_0_T ? phv_data_34 : _GEN_553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_555 = 8'h23 == _match_key_qbytes_0_T ? phv_data_35 : _GEN_554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_556 = 8'h24 == _match_key_qbytes_0_T ? phv_data_36 : _GEN_555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_557 = 8'h25 == _match_key_qbytes_0_T ? phv_data_37 : _GEN_556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_558 = 8'h26 == _match_key_qbytes_0_T ? phv_data_38 : _GEN_557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_559 = 8'h27 == _match_key_qbytes_0_T ? phv_data_39 : _GEN_558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_560 = 8'h28 == _match_key_qbytes_0_T ? phv_data_40 : _GEN_559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_561 = 8'h29 == _match_key_qbytes_0_T ? phv_data_41 : _GEN_560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_562 = 8'h2a == _match_key_qbytes_0_T ? phv_data_42 : _GEN_561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_563 = 8'h2b == _match_key_qbytes_0_T ? phv_data_43 : _GEN_562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_564 = 8'h2c == _match_key_qbytes_0_T ? phv_data_44 : _GEN_563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_565 = 8'h2d == _match_key_qbytes_0_T ? phv_data_45 : _GEN_564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_566 = 8'h2e == _match_key_qbytes_0_T ? phv_data_46 : _GEN_565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_567 = 8'h2f == _match_key_qbytes_0_T ? phv_data_47 : _GEN_566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_568 = 8'h30 == _match_key_qbytes_0_T ? phv_data_48 : _GEN_567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_569 = 8'h31 == _match_key_qbytes_0_T ? phv_data_49 : _GEN_568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_570 = 8'h32 == _match_key_qbytes_0_T ? phv_data_50 : _GEN_569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_571 = 8'h33 == _match_key_qbytes_0_T ? phv_data_51 : _GEN_570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_572 = 8'h34 == _match_key_qbytes_0_T ? phv_data_52 : _GEN_571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_573 = 8'h35 == _match_key_qbytes_0_T ? phv_data_53 : _GEN_572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_574 = 8'h36 == _match_key_qbytes_0_T ? phv_data_54 : _GEN_573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_575 = 8'h37 == _match_key_qbytes_0_T ? phv_data_55 : _GEN_574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_576 = 8'h38 == _match_key_qbytes_0_T ? phv_data_56 : _GEN_575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_577 = 8'h39 == _match_key_qbytes_0_T ? phv_data_57 : _GEN_576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_578 = 8'h3a == _match_key_qbytes_0_T ? phv_data_58 : _GEN_577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_579 = 8'h3b == _match_key_qbytes_0_T ? phv_data_59 : _GEN_578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_580 = 8'h3c == _match_key_qbytes_0_T ? phv_data_60 : _GEN_579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_581 = 8'h3d == _match_key_qbytes_0_T ? phv_data_61 : _GEN_580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_582 = 8'h3e == _match_key_qbytes_0_T ? phv_data_62 : _GEN_581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_583 = 8'h3f == _match_key_qbytes_0_T ? phv_data_63 : _GEN_582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_584 = 8'h40 == _match_key_qbytes_0_T ? phv_data_64 : _GEN_583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_585 = 8'h41 == _match_key_qbytes_0_T ? phv_data_65 : _GEN_584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_586 = 8'h42 == _match_key_qbytes_0_T ? phv_data_66 : _GEN_585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_587 = 8'h43 == _match_key_qbytes_0_T ? phv_data_67 : _GEN_586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_588 = 8'h44 == _match_key_qbytes_0_T ? phv_data_68 : _GEN_587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_589 = 8'h45 == _match_key_qbytes_0_T ? phv_data_69 : _GEN_588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_590 = 8'h46 == _match_key_qbytes_0_T ? phv_data_70 : _GEN_589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_591 = 8'h47 == _match_key_qbytes_0_T ? phv_data_71 : _GEN_590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_592 = 8'h48 == _match_key_qbytes_0_T ? phv_data_72 : _GEN_591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_593 = 8'h49 == _match_key_qbytes_0_T ? phv_data_73 : _GEN_592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_594 = 8'h4a == _match_key_qbytes_0_T ? phv_data_74 : _GEN_593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_595 = 8'h4b == _match_key_qbytes_0_T ? phv_data_75 : _GEN_594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_596 = 8'h4c == _match_key_qbytes_0_T ? phv_data_76 : _GEN_595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_597 = 8'h4d == _match_key_qbytes_0_T ? phv_data_77 : _GEN_596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_598 = 8'h4e == _match_key_qbytes_0_T ? phv_data_78 : _GEN_597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_599 = 8'h4f == _match_key_qbytes_0_T ? phv_data_79 : _GEN_598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_600 = 8'h50 == _match_key_qbytes_0_T ? phv_data_80 : _GEN_599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_601 = 8'h51 == _match_key_qbytes_0_T ? phv_data_81 : _GEN_600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_602 = 8'h52 == _match_key_qbytes_0_T ? phv_data_82 : _GEN_601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_603 = 8'h53 == _match_key_qbytes_0_T ? phv_data_83 : _GEN_602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_604 = 8'h54 == _match_key_qbytes_0_T ? phv_data_84 : _GEN_603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_605 = 8'h55 == _match_key_qbytes_0_T ? phv_data_85 : _GEN_604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_606 = 8'h56 == _match_key_qbytes_0_T ? phv_data_86 : _GEN_605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_607 = 8'h57 == _match_key_qbytes_0_T ? phv_data_87 : _GEN_606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_608 = 8'h58 == _match_key_qbytes_0_T ? phv_data_88 : _GEN_607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_609 = 8'h59 == _match_key_qbytes_0_T ? phv_data_89 : _GEN_608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_610 = 8'h5a == _match_key_qbytes_0_T ? phv_data_90 : _GEN_609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_611 = 8'h5b == _match_key_qbytes_0_T ? phv_data_91 : _GEN_610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_612 = 8'h5c == _match_key_qbytes_0_T ? phv_data_92 : _GEN_611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_613 = 8'h5d == _match_key_qbytes_0_T ? phv_data_93 : _GEN_612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_614 = 8'h5e == _match_key_qbytes_0_T ? phv_data_94 : _GEN_613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_615 = 8'h5f == _match_key_qbytes_0_T ? phv_data_95 : _GEN_614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_616 = 8'h60 == _match_key_qbytes_0_T ? phv_data_96 : _GEN_615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_617 = 8'h61 == _match_key_qbytes_0_T ? phv_data_97 : _GEN_616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_618 = 8'h62 == _match_key_qbytes_0_T ? phv_data_98 : _GEN_617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_619 = 8'h63 == _match_key_qbytes_0_T ? phv_data_99 : _GEN_618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_620 = 8'h64 == _match_key_qbytes_0_T ? phv_data_100 : _GEN_619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_621 = 8'h65 == _match_key_qbytes_0_T ? phv_data_101 : _GEN_620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_622 = 8'h66 == _match_key_qbytes_0_T ? phv_data_102 : _GEN_621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_623 = 8'h67 == _match_key_qbytes_0_T ? phv_data_103 : _GEN_622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_624 = 8'h68 == _match_key_qbytes_0_T ? phv_data_104 : _GEN_623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_625 = 8'h69 == _match_key_qbytes_0_T ? phv_data_105 : _GEN_624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_626 = 8'h6a == _match_key_qbytes_0_T ? phv_data_106 : _GEN_625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_627 = 8'h6b == _match_key_qbytes_0_T ? phv_data_107 : _GEN_626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_628 = 8'h6c == _match_key_qbytes_0_T ? phv_data_108 : _GEN_627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_629 = 8'h6d == _match_key_qbytes_0_T ? phv_data_109 : _GEN_628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_630 = 8'h6e == _match_key_qbytes_0_T ? phv_data_110 : _GEN_629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_631 = 8'h6f == _match_key_qbytes_0_T ? phv_data_111 : _GEN_630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_632 = 8'h70 == _match_key_qbytes_0_T ? phv_data_112 : _GEN_631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_633 = 8'h71 == _match_key_qbytes_0_T ? phv_data_113 : _GEN_632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_634 = 8'h72 == _match_key_qbytes_0_T ? phv_data_114 : _GEN_633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_635 = 8'h73 == _match_key_qbytes_0_T ? phv_data_115 : _GEN_634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_636 = 8'h74 == _match_key_qbytes_0_T ? phv_data_116 : _GEN_635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_637 = 8'h75 == _match_key_qbytes_0_T ? phv_data_117 : _GEN_636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_638 = 8'h76 == _match_key_qbytes_0_T ? phv_data_118 : _GEN_637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_639 = 8'h77 == _match_key_qbytes_0_T ? phv_data_119 : _GEN_638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_640 = 8'h78 == _match_key_qbytes_0_T ? phv_data_120 : _GEN_639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_641 = 8'h79 == _match_key_qbytes_0_T ? phv_data_121 : _GEN_640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_642 = 8'h7a == _match_key_qbytes_0_T ? phv_data_122 : _GEN_641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_643 = 8'h7b == _match_key_qbytes_0_T ? phv_data_123 : _GEN_642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_644 = 8'h7c == _match_key_qbytes_0_T ? phv_data_124 : _GEN_643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_645 = 8'h7d == _match_key_qbytes_0_T ? phv_data_125 : _GEN_644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_646 = 8'h7e == _match_key_qbytes_0_T ? phv_data_126 : _GEN_645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_647 = 8'h7f == _match_key_qbytes_0_T ? phv_data_127 : _GEN_646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_648 = 8'h80 == _match_key_qbytes_0_T ? phv_data_128 : _GEN_647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_649 = 8'h81 == _match_key_qbytes_0_T ? phv_data_129 : _GEN_648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_650 = 8'h82 == _match_key_qbytes_0_T ? phv_data_130 : _GEN_649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_651 = 8'h83 == _match_key_qbytes_0_T ? phv_data_131 : _GEN_650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_652 = 8'h84 == _match_key_qbytes_0_T ? phv_data_132 : _GEN_651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_653 = 8'h85 == _match_key_qbytes_0_T ? phv_data_133 : _GEN_652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_654 = 8'h86 == _match_key_qbytes_0_T ? phv_data_134 : _GEN_653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_655 = 8'h87 == _match_key_qbytes_0_T ? phv_data_135 : _GEN_654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_656 = 8'h88 == _match_key_qbytes_0_T ? phv_data_136 : _GEN_655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_657 = 8'h89 == _match_key_qbytes_0_T ? phv_data_137 : _GEN_656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_658 = 8'h8a == _match_key_qbytes_0_T ? phv_data_138 : _GEN_657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_659 = 8'h8b == _match_key_qbytes_0_T ? phv_data_139 : _GEN_658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_660 = 8'h8c == _match_key_qbytes_0_T ? phv_data_140 : _GEN_659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_661 = 8'h8d == _match_key_qbytes_0_T ? phv_data_141 : _GEN_660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_662 = 8'h8e == _match_key_qbytes_0_T ? phv_data_142 : _GEN_661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_663 = 8'h8f == _match_key_qbytes_0_T ? phv_data_143 : _GEN_662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_664 = 8'h90 == _match_key_qbytes_0_T ? phv_data_144 : _GEN_663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_665 = 8'h91 == _match_key_qbytes_0_T ? phv_data_145 : _GEN_664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_666 = 8'h92 == _match_key_qbytes_0_T ? phv_data_146 : _GEN_665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_667 = 8'h93 == _match_key_qbytes_0_T ? phv_data_147 : _GEN_666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_668 = 8'h94 == _match_key_qbytes_0_T ? phv_data_148 : _GEN_667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_669 = 8'h95 == _match_key_qbytes_0_T ? phv_data_149 : _GEN_668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_670 = 8'h96 == _match_key_qbytes_0_T ? phv_data_150 : _GEN_669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_671 = 8'h97 == _match_key_qbytes_0_T ? phv_data_151 : _GEN_670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_672 = 8'h98 == _match_key_qbytes_0_T ? phv_data_152 : _GEN_671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_673 = 8'h99 == _match_key_qbytes_0_T ? phv_data_153 : _GEN_672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_674 = 8'h9a == _match_key_qbytes_0_T ? phv_data_154 : _GEN_673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_675 = 8'h9b == _match_key_qbytes_0_T ? phv_data_155 : _GEN_674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_676 = 8'h9c == _match_key_qbytes_0_T ? phv_data_156 : _GEN_675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_677 = 8'h9d == _match_key_qbytes_0_T ? phv_data_157 : _GEN_676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_678 = 8'h9e == _match_key_qbytes_0_T ? phv_data_158 : _GEN_677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_679 = 8'h9f == _match_key_qbytes_0_T ? phv_data_159 : _GEN_678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_680 = 8'ha0 == _match_key_qbytes_0_T ? phv_data_160 : _GEN_679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_681 = 8'ha1 == _match_key_qbytes_0_T ? phv_data_161 : _GEN_680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_682 = 8'ha2 == _match_key_qbytes_0_T ? phv_data_162 : _GEN_681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_683 = 8'ha3 == _match_key_qbytes_0_T ? phv_data_163 : _GEN_682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_684 = 8'ha4 == _match_key_qbytes_0_T ? phv_data_164 : _GEN_683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_685 = 8'ha5 == _match_key_qbytes_0_T ? phv_data_165 : _GEN_684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_686 = 8'ha6 == _match_key_qbytes_0_T ? phv_data_166 : _GEN_685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_687 = 8'ha7 == _match_key_qbytes_0_T ? phv_data_167 : _GEN_686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_688 = 8'ha8 == _match_key_qbytes_0_T ? phv_data_168 : _GEN_687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_689 = 8'ha9 == _match_key_qbytes_0_T ? phv_data_169 : _GEN_688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_690 = 8'haa == _match_key_qbytes_0_T ? phv_data_170 : _GEN_689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_691 = 8'hab == _match_key_qbytes_0_T ? phv_data_171 : _GEN_690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_692 = 8'hac == _match_key_qbytes_0_T ? phv_data_172 : _GEN_691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_693 = 8'had == _match_key_qbytes_0_T ? phv_data_173 : _GEN_692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_694 = 8'hae == _match_key_qbytes_0_T ? phv_data_174 : _GEN_693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_695 = 8'haf == _match_key_qbytes_0_T ? phv_data_175 : _GEN_694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_696 = 8'hb0 == _match_key_qbytes_0_T ? phv_data_176 : _GEN_695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_697 = 8'hb1 == _match_key_qbytes_0_T ? phv_data_177 : _GEN_696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_698 = 8'hb2 == _match_key_qbytes_0_T ? phv_data_178 : _GEN_697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_699 = 8'hb3 == _match_key_qbytes_0_T ? phv_data_179 : _GEN_698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_700 = 8'hb4 == _match_key_qbytes_0_T ? phv_data_180 : _GEN_699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_701 = 8'hb5 == _match_key_qbytes_0_T ? phv_data_181 : _GEN_700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_702 = 8'hb6 == _match_key_qbytes_0_T ? phv_data_182 : _GEN_701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_703 = 8'hb7 == _match_key_qbytes_0_T ? phv_data_183 : _GEN_702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_704 = 8'hb8 == _match_key_qbytes_0_T ? phv_data_184 : _GEN_703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_705 = 8'hb9 == _match_key_qbytes_0_T ? phv_data_185 : _GEN_704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_706 = 8'hba == _match_key_qbytes_0_T ? phv_data_186 : _GEN_705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_707 = 8'hbb == _match_key_qbytes_0_T ? phv_data_187 : _GEN_706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_708 = 8'hbc == _match_key_qbytes_0_T ? phv_data_188 : _GEN_707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_709 = 8'hbd == _match_key_qbytes_0_T ? phv_data_189 : _GEN_708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_710 = 8'hbe == _match_key_qbytes_0_T ? phv_data_190 : _GEN_709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_711 = 8'hbf == _match_key_qbytes_0_T ? phv_data_191 : _GEN_710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_712 = 8'hc0 == _match_key_qbytes_0_T ? phv_data_192 : _GEN_711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_713 = 8'hc1 == _match_key_qbytes_0_T ? phv_data_193 : _GEN_712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_714 = 8'hc2 == _match_key_qbytes_0_T ? phv_data_194 : _GEN_713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_715 = 8'hc3 == _match_key_qbytes_0_T ? phv_data_195 : _GEN_714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_716 = 8'hc4 == _match_key_qbytes_0_T ? phv_data_196 : _GEN_715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_717 = 8'hc5 == _match_key_qbytes_0_T ? phv_data_197 : _GEN_716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_718 = 8'hc6 == _match_key_qbytes_0_T ? phv_data_198 : _GEN_717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_719 = 8'hc7 == _match_key_qbytes_0_T ? phv_data_199 : _GEN_718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_720 = 8'hc8 == _match_key_qbytes_0_T ? phv_data_200 : _GEN_719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_721 = 8'hc9 == _match_key_qbytes_0_T ? phv_data_201 : _GEN_720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_722 = 8'hca == _match_key_qbytes_0_T ? phv_data_202 : _GEN_721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_723 = 8'hcb == _match_key_qbytes_0_T ? phv_data_203 : _GEN_722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_724 = 8'hcc == _match_key_qbytes_0_T ? phv_data_204 : _GEN_723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_725 = 8'hcd == _match_key_qbytes_0_T ? phv_data_205 : _GEN_724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_726 = 8'hce == _match_key_qbytes_0_T ? phv_data_206 : _GEN_725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_727 = 8'hcf == _match_key_qbytes_0_T ? phv_data_207 : _GEN_726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_728 = 8'hd0 == _match_key_qbytes_0_T ? phv_data_208 : _GEN_727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_729 = 8'hd1 == _match_key_qbytes_0_T ? phv_data_209 : _GEN_728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_730 = 8'hd2 == _match_key_qbytes_0_T ? phv_data_210 : _GEN_729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_731 = 8'hd3 == _match_key_qbytes_0_T ? phv_data_211 : _GEN_730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_732 = 8'hd4 == _match_key_qbytes_0_T ? phv_data_212 : _GEN_731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_733 = 8'hd5 == _match_key_qbytes_0_T ? phv_data_213 : _GEN_732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_734 = 8'hd6 == _match_key_qbytes_0_T ? phv_data_214 : _GEN_733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_735 = 8'hd7 == _match_key_qbytes_0_T ? phv_data_215 : _GEN_734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_736 = 8'hd8 == _match_key_qbytes_0_T ? phv_data_216 : _GEN_735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_737 = 8'hd9 == _match_key_qbytes_0_T ? phv_data_217 : _GEN_736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_738 = 8'hda == _match_key_qbytes_0_T ? phv_data_218 : _GEN_737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_739 = 8'hdb == _match_key_qbytes_0_T ? phv_data_219 : _GEN_738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_740 = 8'hdc == _match_key_qbytes_0_T ? phv_data_220 : _GEN_739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_741 = 8'hdd == _match_key_qbytes_0_T ? phv_data_221 : _GEN_740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_742 = 8'hde == _match_key_qbytes_0_T ? phv_data_222 : _GEN_741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_743 = 8'hdf == _match_key_qbytes_0_T ? phv_data_223 : _GEN_742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_744 = 8'he0 == _match_key_qbytes_0_T ? phv_data_224 : _GEN_743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_745 = 8'he1 == _match_key_qbytes_0_T ? phv_data_225 : _GEN_744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_746 = 8'he2 == _match_key_qbytes_0_T ? phv_data_226 : _GEN_745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_747 = 8'he3 == _match_key_qbytes_0_T ? phv_data_227 : _GEN_746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_748 = 8'he4 == _match_key_qbytes_0_T ? phv_data_228 : _GEN_747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_749 = 8'he5 == _match_key_qbytes_0_T ? phv_data_229 : _GEN_748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_750 = 8'he6 == _match_key_qbytes_0_T ? phv_data_230 : _GEN_749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_751 = 8'he7 == _match_key_qbytes_0_T ? phv_data_231 : _GEN_750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_752 = 8'he8 == _match_key_qbytes_0_T ? phv_data_232 : _GEN_751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_753 = 8'he9 == _match_key_qbytes_0_T ? phv_data_233 : _GEN_752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_754 = 8'hea == _match_key_qbytes_0_T ? phv_data_234 : _GEN_753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_755 = 8'heb == _match_key_qbytes_0_T ? phv_data_235 : _GEN_754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_756 = 8'hec == _match_key_qbytes_0_T ? phv_data_236 : _GEN_755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_757 = 8'hed == _match_key_qbytes_0_T ? phv_data_237 : _GEN_756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_758 = 8'hee == _match_key_qbytes_0_T ? phv_data_238 : _GEN_757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_759 = 8'hef == _match_key_qbytes_0_T ? phv_data_239 : _GEN_758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_760 = 8'hf0 == _match_key_qbytes_0_T ? phv_data_240 : _GEN_759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_761 = 8'hf1 == _match_key_qbytes_0_T ? phv_data_241 : _GEN_760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_762 = 8'hf2 == _match_key_qbytes_0_T ? phv_data_242 : _GEN_761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_763 = 8'hf3 == _match_key_qbytes_0_T ? phv_data_243 : _GEN_762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_764 = 8'hf4 == _match_key_qbytes_0_T ? phv_data_244 : _GEN_763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_765 = 8'hf5 == _match_key_qbytes_0_T ? phv_data_245 : _GEN_764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_766 = 8'hf6 == _match_key_qbytes_0_T ? phv_data_246 : _GEN_765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_767 = 8'hf7 == _match_key_qbytes_0_T ? phv_data_247 : _GEN_766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_768 = 8'hf8 == _match_key_qbytes_0_T ? phv_data_248 : _GEN_767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_769 = 8'hf9 == _match_key_qbytes_0_T ? phv_data_249 : _GEN_768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_770 = 8'hfa == _match_key_qbytes_0_T ? phv_data_250 : _GEN_769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_771 = 8'hfb == _match_key_qbytes_0_T ? phv_data_251 : _GEN_770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_772 = 8'hfc == _match_key_qbytes_0_T ? phv_data_252 : _GEN_771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_773 = 8'hfd == _match_key_qbytes_0_T ? phv_data_253 : _GEN_772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_774 = 8'hfe == _match_key_qbytes_0_T ? phv_data_254 : _GEN_773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_775 = 8'hff == _match_key_qbytes_0_T ? phv_data_255 : _GEN_774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_777 = 8'h1 == _match_key_qbytes_0_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_778 = 8'h2 == _match_key_qbytes_0_T_1 ? phv_data_2 : _GEN_777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_779 = 8'h3 == _match_key_qbytes_0_T_1 ? phv_data_3 : _GEN_778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_780 = 8'h4 == _match_key_qbytes_0_T_1 ? phv_data_4 : _GEN_779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_781 = 8'h5 == _match_key_qbytes_0_T_1 ? phv_data_5 : _GEN_780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_782 = 8'h6 == _match_key_qbytes_0_T_1 ? phv_data_6 : _GEN_781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_783 = 8'h7 == _match_key_qbytes_0_T_1 ? phv_data_7 : _GEN_782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_784 = 8'h8 == _match_key_qbytes_0_T_1 ? phv_data_8 : _GEN_783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_785 = 8'h9 == _match_key_qbytes_0_T_1 ? phv_data_9 : _GEN_784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_786 = 8'ha == _match_key_qbytes_0_T_1 ? phv_data_10 : _GEN_785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_787 = 8'hb == _match_key_qbytes_0_T_1 ? phv_data_11 : _GEN_786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_788 = 8'hc == _match_key_qbytes_0_T_1 ? phv_data_12 : _GEN_787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_789 = 8'hd == _match_key_qbytes_0_T_1 ? phv_data_13 : _GEN_788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_790 = 8'he == _match_key_qbytes_0_T_1 ? phv_data_14 : _GEN_789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_791 = 8'hf == _match_key_qbytes_0_T_1 ? phv_data_15 : _GEN_790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_792 = 8'h10 == _match_key_qbytes_0_T_1 ? phv_data_16 : _GEN_791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_793 = 8'h11 == _match_key_qbytes_0_T_1 ? phv_data_17 : _GEN_792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_794 = 8'h12 == _match_key_qbytes_0_T_1 ? phv_data_18 : _GEN_793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_795 = 8'h13 == _match_key_qbytes_0_T_1 ? phv_data_19 : _GEN_794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_796 = 8'h14 == _match_key_qbytes_0_T_1 ? phv_data_20 : _GEN_795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_797 = 8'h15 == _match_key_qbytes_0_T_1 ? phv_data_21 : _GEN_796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_798 = 8'h16 == _match_key_qbytes_0_T_1 ? phv_data_22 : _GEN_797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_799 = 8'h17 == _match_key_qbytes_0_T_1 ? phv_data_23 : _GEN_798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_800 = 8'h18 == _match_key_qbytes_0_T_1 ? phv_data_24 : _GEN_799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_801 = 8'h19 == _match_key_qbytes_0_T_1 ? phv_data_25 : _GEN_800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_802 = 8'h1a == _match_key_qbytes_0_T_1 ? phv_data_26 : _GEN_801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_803 = 8'h1b == _match_key_qbytes_0_T_1 ? phv_data_27 : _GEN_802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_804 = 8'h1c == _match_key_qbytes_0_T_1 ? phv_data_28 : _GEN_803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_805 = 8'h1d == _match_key_qbytes_0_T_1 ? phv_data_29 : _GEN_804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_806 = 8'h1e == _match_key_qbytes_0_T_1 ? phv_data_30 : _GEN_805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_807 = 8'h1f == _match_key_qbytes_0_T_1 ? phv_data_31 : _GEN_806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_808 = 8'h20 == _match_key_qbytes_0_T_1 ? phv_data_32 : _GEN_807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_809 = 8'h21 == _match_key_qbytes_0_T_1 ? phv_data_33 : _GEN_808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_810 = 8'h22 == _match_key_qbytes_0_T_1 ? phv_data_34 : _GEN_809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_811 = 8'h23 == _match_key_qbytes_0_T_1 ? phv_data_35 : _GEN_810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_812 = 8'h24 == _match_key_qbytes_0_T_1 ? phv_data_36 : _GEN_811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_813 = 8'h25 == _match_key_qbytes_0_T_1 ? phv_data_37 : _GEN_812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_814 = 8'h26 == _match_key_qbytes_0_T_1 ? phv_data_38 : _GEN_813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_815 = 8'h27 == _match_key_qbytes_0_T_1 ? phv_data_39 : _GEN_814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_816 = 8'h28 == _match_key_qbytes_0_T_1 ? phv_data_40 : _GEN_815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_817 = 8'h29 == _match_key_qbytes_0_T_1 ? phv_data_41 : _GEN_816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_818 = 8'h2a == _match_key_qbytes_0_T_1 ? phv_data_42 : _GEN_817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_819 = 8'h2b == _match_key_qbytes_0_T_1 ? phv_data_43 : _GEN_818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_820 = 8'h2c == _match_key_qbytes_0_T_1 ? phv_data_44 : _GEN_819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_821 = 8'h2d == _match_key_qbytes_0_T_1 ? phv_data_45 : _GEN_820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_822 = 8'h2e == _match_key_qbytes_0_T_1 ? phv_data_46 : _GEN_821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_823 = 8'h2f == _match_key_qbytes_0_T_1 ? phv_data_47 : _GEN_822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_824 = 8'h30 == _match_key_qbytes_0_T_1 ? phv_data_48 : _GEN_823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_825 = 8'h31 == _match_key_qbytes_0_T_1 ? phv_data_49 : _GEN_824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_826 = 8'h32 == _match_key_qbytes_0_T_1 ? phv_data_50 : _GEN_825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_827 = 8'h33 == _match_key_qbytes_0_T_1 ? phv_data_51 : _GEN_826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_828 = 8'h34 == _match_key_qbytes_0_T_1 ? phv_data_52 : _GEN_827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_829 = 8'h35 == _match_key_qbytes_0_T_1 ? phv_data_53 : _GEN_828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_830 = 8'h36 == _match_key_qbytes_0_T_1 ? phv_data_54 : _GEN_829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_831 = 8'h37 == _match_key_qbytes_0_T_1 ? phv_data_55 : _GEN_830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_832 = 8'h38 == _match_key_qbytes_0_T_1 ? phv_data_56 : _GEN_831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_833 = 8'h39 == _match_key_qbytes_0_T_1 ? phv_data_57 : _GEN_832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_834 = 8'h3a == _match_key_qbytes_0_T_1 ? phv_data_58 : _GEN_833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_835 = 8'h3b == _match_key_qbytes_0_T_1 ? phv_data_59 : _GEN_834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_836 = 8'h3c == _match_key_qbytes_0_T_1 ? phv_data_60 : _GEN_835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_837 = 8'h3d == _match_key_qbytes_0_T_1 ? phv_data_61 : _GEN_836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_838 = 8'h3e == _match_key_qbytes_0_T_1 ? phv_data_62 : _GEN_837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_839 = 8'h3f == _match_key_qbytes_0_T_1 ? phv_data_63 : _GEN_838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_840 = 8'h40 == _match_key_qbytes_0_T_1 ? phv_data_64 : _GEN_839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_841 = 8'h41 == _match_key_qbytes_0_T_1 ? phv_data_65 : _GEN_840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_842 = 8'h42 == _match_key_qbytes_0_T_1 ? phv_data_66 : _GEN_841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_843 = 8'h43 == _match_key_qbytes_0_T_1 ? phv_data_67 : _GEN_842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_844 = 8'h44 == _match_key_qbytes_0_T_1 ? phv_data_68 : _GEN_843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_845 = 8'h45 == _match_key_qbytes_0_T_1 ? phv_data_69 : _GEN_844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_846 = 8'h46 == _match_key_qbytes_0_T_1 ? phv_data_70 : _GEN_845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_847 = 8'h47 == _match_key_qbytes_0_T_1 ? phv_data_71 : _GEN_846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_848 = 8'h48 == _match_key_qbytes_0_T_1 ? phv_data_72 : _GEN_847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_849 = 8'h49 == _match_key_qbytes_0_T_1 ? phv_data_73 : _GEN_848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_850 = 8'h4a == _match_key_qbytes_0_T_1 ? phv_data_74 : _GEN_849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_851 = 8'h4b == _match_key_qbytes_0_T_1 ? phv_data_75 : _GEN_850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_852 = 8'h4c == _match_key_qbytes_0_T_1 ? phv_data_76 : _GEN_851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_853 = 8'h4d == _match_key_qbytes_0_T_1 ? phv_data_77 : _GEN_852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_854 = 8'h4e == _match_key_qbytes_0_T_1 ? phv_data_78 : _GEN_853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_855 = 8'h4f == _match_key_qbytes_0_T_1 ? phv_data_79 : _GEN_854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_856 = 8'h50 == _match_key_qbytes_0_T_1 ? phv_data_80 : _GEN_855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_857 = 8'h51 == _match_key_qbytes_0_T_1 ? phv_data_81 : _GEN_856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_858 = 8'h52 == _match_key_qbytes_0_T_1 ? phv_data_82 : _GEN_857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_859 = 8'h53 == _match_key_qbytes_0_T_1 ? phv_data_83 : _GEN_858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_860 = 8'h54 == _match_key_qbytes_0_T_1 ? phv_data_84 : _GEN_859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_861 = 8'h55 == _match_key_qbytes_0_T_1 ? phv_data_85 : _GEN_860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_862 = 8'h56 == _match_key_qbytes_0_T_1 ? phv_data_86 : _GEN_861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_863 = 8'h57 == _match_key_qbytes_0_T_1 ? phv_data_87 : _GEN_862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_864 = 8'h58 == _match_key_qbytes_0_T_1 ? phv_data_88 : _GEN_863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_865 = 8'h59 == _match_key_qbytes_0_T_1 ? phv_data_89 : _GEN_864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_866 = 8'h5a == _match_key_qbytes_0_T_1 ? phv_data_90 : _GEN_865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_867 = 8'h5b == _match_key_qbytes_0_T_1 ? phv_data_91 : _GEN_866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_868 = 8'h5c == _match_key_qbytes_0_T_1 ? phv_data_92 : _GEN_867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_869 = 8'h5d == _match_key_qbytes_0_T_1 ? phv_data_93 : _GEN_868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_870 = 8'h5e == _match_key_qbytes_0_T_1 ? phv_data_94 : _GEN_869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_871 = 8'h5f == _match_key_qbytes_0_T_1 ? phv_data_95 : _GEN_870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_872 = 8'h60 == _match_key_qbytes_0_T_1 ? phv_data_96 : _GEN_871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_873 = 8'h61 == _match_key_qbytes_0_T_1 ? phv_data_97 : _GEN_872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_874 = 8'h62 == _match_key_qbytes_0_T_1 ? phv_data_98 : _GEN_873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_875 = 8'h63 == _match_key_qbytes_0_T_1 ? phv_data_99 : _GEN_874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_876 = 8'h64 == _match_key_qbytes_0_T_1 ? phv_data_100 : _GEN_875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_877 = 8'h65 == _match_key_qbytes_0_T_1 ? phv_data_101 : _GEN_876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_878 = 8'h66 == _match_key_qbytes_0_T_1 ? phv_data_102 : _GEN_877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_879 = 8'h67 == _match_key_qbytes_0_T_1 ? phv_data_103 : _GEN_878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_880 = 8'h68 == _match_key_qbytes_0_T_1 ? phv_data_104 : _GEN_879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_881 = 8'h69 == _match_key_qbytes_0_T_1 ? phv_data_105 : _GEN_880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_882 = 8'h6a == _match_key_qbytes_0_T_1 ? phv_data_106 : _GEN_881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_883 = 8'h6b == _match_key_qbytes_0_T_1 ? phv_data_107 : _GEN_882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_884 = 8'h6c == _match_key_qbytes_0_T_1 ? phv_data_108 : _GEN_883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_885 = 8'h6d == _match_key_qbytes_0_T_1 ? phv_data_109 : _GEN_884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_886 = 8'h6e == _match_key_qbytes_0_T_1 ? phv_data_110 : _GEN_885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_887 = 8'h6f == _match_key_qbytes_0_T_1 ? phv_data_111 : _GEN_886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_888 = 8'h70 == _match_key_qbytes_0_T_1 ? phv_data_112 : _GEN_887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_889 = 8'h71 == _match_key_qbytes_0_T_1 ? phv_data_113 : _GEN_888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_890 = 8'h72 == _match_key_qbytes_0_T_1 ? phv_data_114 : _GEN_889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_891 = 8'h73 == _match_key_qbytes_0_T_1 ? phv_data_115 : _GEN_890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_892 = 8'h74 == _match_key_qbytes_0_T_1 ? phv_data_116 : _GEN_891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_893 = 8'h75 == _match_key_qbytes_0_T_1 ? phv_data_117 : _GEN_892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_894 = 8'h76 == _match_key_qbytes_0_T_1 ? phv_data_118 : _GEN_893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_895 = 8'h77 == _match_key_qbytes_0_T_1 ? phv_data_119 : _GEN_894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_896 = 8'h78 == _match_key_qbytes_0_T_1 ? phv_data_120 : _GEN_895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_897 = 8'h79 == _match_key_qbytes_0_T_1 ? phv_data_121 : _GEN_896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_898 = 8'h7a == _match_key_qbytes_0_T_1 ? phv_data_122 : _GEN_897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_899 = 8'h7b == _match_key_qbytes_0_T_1 ? phv_data_123 : _GEN_898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_900 = 8'h7c == _match_key_qbytes_0_T_1 ? phv_data_124 : _GEN_899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_901 = 8'h7d == _match_key_qbytes_0_T_1 ? phv_data_125 : _GEN_900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_902 = 8'h7e == _match_key_qbytes_0_T_1 ? phv_data_126 : _GEN_901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_903 = 8'h7f == _match_key_qbytes_0_T_1 ? phv_data_127 : _GEN_902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_904 = 8'h80 == _match_key_qbytes_0_T_1 ? phv_data_128 : _GEN_903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_905 = 8'h81 == _match_key_qbytes_0_T_1 ? phv_data_129 : _GEN_904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_906 = 8'h82 == _match_key_qbytes_0_T_1 ? phv_data_130 : _GEN_905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_907 = 8'h83 == _match_key_qbytes_0_T_1 ? phv_data_131 : _GEN_906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_908 = 8'h84 == _match_key_qbytes_0_T_1 ? phv_data_132 : _GEN_907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_909 = 8'h85 == _match_key_qbytes_0_T_1 ? phv_data_133 : _GEN_908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_910 = 8'h86 == _match_key_qbytes_0_T_1 ? phv_data_134 : _GEN_909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_911 = 8'h87 == _match_key_qbytes_0_T_1 ? phv_data_135 : _GEN_910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_912 = 8'h88 == _match_key_qbytes_0_T_1 ? phv_data_136 : _GEN_911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_913 = 8'h89 == _match_key_qbytes_0_T_1 ? phv_data_137 : _GEN_912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_914 = 8'h8a == _match_key_qbytes_0_T_1 ? phv_data_138 : _GEN_913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_915 = 8'h8b == _match_key_qbytes_0_T_1 ? phv_data_139 : _GEN_914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_916 = 8'h8c == _match_key_qbytes_0_T_1 ? phv_data_140 : _GEN_915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_917 = 8'h8d == _match_key_qbytes_0_T_1 ? phv_data_141 : _GEN_916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_918 = 8'h8e == _match_key_qbytes_0_T_1 ? phv_data_142 : _GEN_917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_919 = 8'h8f == _match_key_qbytes_0_T_1 ? phv_data_143 : _GEN_918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_920 = 8'h90 == _match_key_qbytes_0_T_1 ? phv_data_144 : _GEN_919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_921 = 8'h91 == _match_key_qbytes_0_T_1 ? phv_data_145 : _GEN_920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_922 = 8'h92 == _match_key_qbytes_0_T_1 ? phv_data_146 : _GEN_921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_923 = 8'h93 == _match_key_qbytes_0_T_1 ? phv_data_147 : _GEN_922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_924 = 8'h94 == _match_key_qbytes_0_T_1 ? phv_data_148 : _GEN_923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_925 = 8'h95 == _match_key_qbytes_0_T_1 ? phv_data_149 : _GEN_924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_926 = 8'h96 == _match_key_qbytes_0_T_1 ? phv_data_150 : _GEN_925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_927 = 8'h97 == _match_key_qbytes_0_T_1 ? phv_data_151 : _GEN_926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_928 = 8'h98 == _match_key_qbytes_0_T_1 ? phv_data_152 : _GEN_927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_929 = 8'h99 == _match_key_qbytes_0_T_1 ? phv_data_153 : _GEN_928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_930 = 8'h9a == _match_key_qbytes_0_T_1 ? phv_data_154 : _GEN_929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_931 = 8'h9b == _match_key_qbytes_0_T_1 ? phv_data_155 : _GEN_930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_932 = 8'h9c == _match_key_qbytes_0_T_1 ? phv_data_156 : _GEN_931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_933 = 8'h9d == _match_key_qbytes_0_T_1 ? phv_data_157 : _GEN_932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_934 = 8'h9e == _match_key_qbytes_0_T_1 ? phv_data_158 : _GEN_933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_935 = 8'h9f == _match_key_qbytes_0_T_1 ? phv_data_159 : _GEN_934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_936 = 8'ha0 == _match_key_qbytes_0_T_1 ? phv_data_160 : _GEN_935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_937 = 8'ha1 == _match_key_qbytes_0_T_1 ? phv_data_161 : _GEN_936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_938 = 8'ha2 == _match_key_qbytes_0_T_1 ? phv_data_162 : _GEN_937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_939 = 8'ha3 == _match_key_qbytes_0_T_1 ? phv_data_163 : _GEN_938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_940 = 8'ha4 == _match_key_qbytes_0_T_1 ? phv_data_164 : _GEN_939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_941 = 8'ha5 == _match_key_qbytes_0_T_1 ? phv_data_165 : _GEN_940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_942 = 8'ha6 == _match_key_qbytes_0_T_1 ? phv_data_166 : _GEN_941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_943 = 8'ha7 == _match_key_qbytes_0_T_1 ? phv_data_167 : _GEN_942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_944 = 8'ha8 == _match_key_qbytes_0_T_1 ? phv_data_168 : _GEN_943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_945 = 8'ha9 == _match_key_qbytes_0_T_1 ? phv_data_169 : _GEN_944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_946 = 8'haa == _match_key_qbytes_0_T_1 ? phv_data_170 : _GEN_945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_947 = 8'hab == _match_key_qbytes_0_T_1 ? phv_data_171 : _GEN_946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_948 = 8'hac == _match_key_qbytes_0_T_1 ? phv_data_172 : _GEN_947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_949 = 8'had == _match_key_qbytes_0_T_1 ? phv_data_173 : _GEN_948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_950 = 8'hae == _match_key_qbytes_0_T_1 ? phv_data_174 : _GEN_949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_951 = 8'haf == _match_key_qbytes_0_T_1 ? phv_data_175 : _GEN_950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_952 = 8'hb0 == _match_key_qbytes_0_T_1 ? phv_data_176 : _GEN_951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_953 = 8'hb1 == _match_key_qbytes_0_T_1 ? phv_data_177 : _GEN_952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_954 = 8'hb2 == _match_key_qbytes_0_T_1 ? phv_data_178 : _GEN_953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_955 = 8'hb3 == _match_key_qbytes_0_T_1 ? phv_data_179 : _GEN_954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_956 = 8'hb4 == _match_key_qbytes_0_T_1 ? phv_data_180 : _GEN_955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_957 = 8'hb5 == _match_key_qbytes_0_T_1 ? phv_data_181 : _GEN_956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_958 = 8'hb6 == _match_key_qbytes_0_T_1 ? phv_data_182 : _GEN_957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_959 = 8'hb7 == _match_key_qbytes_0_T_1 ? phv_data_183 : _GEN_958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_960 = 8'hb8 == _match_key_qbytes_0_T_1 ? phv_data_184 : _GEN_959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_961 = 8'hb9 == _match_key_qbytes_0_T_1 ? phv_data_185 : _GEN_960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_962 = 8'hba == _match_key_qbytes_0_T_1 ? phv_data_186 : _GEN_961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_963 = 8'hbb == _match_key_qbytes_0_T_1 ? phv_data_187 : _GEN_962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_964 = 8'hbc == _match_key_qbytes_0_T_1 ? phv_data_188 : _GEN_963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_965 = 8'hbd == _match_key_qbytes_0_T_1 ? phv_data_189 : _GEN_964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_966 = 8'hbe == _match_key_qbytes_0_T_1 ? phv_data_190 : _GEN_965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_967 = 8'hbf == _match_key_qbytes_0_T_1 ? phv_data_191 : _GEN_966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_968 = 8'hc0 == _match_key_qbytes_0_T_1 ? phv_data_192 : _GEN_967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_969 = 8'hc1 == _match_key_qbytes_0_T_1 ? phv_data_193 : _GEN_968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_970 = 8'hc2 == _match_key_qbytes_0_T_1 ? phv_data_194 : _GEN_969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_971 = 8'hc3 == _match_key_qbytes_0_T_1 ? phv_data_195 : _GEN_970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_972 = 8'hc4 == _match_key_qbytes_0_T_1 ? phv_data_196 : _GEN_971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_973 = 8'hc5 == _match_key_qbytes_0_T_1 ? phv_data_197 : _GEN_972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_974 = 8'hc6 == _match_key_qbytes_0_T_1 ? phv_data_198 : _GEN_973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_975 = 8'hc7 == _match_key_qbytes_0_T_1 ? phv_data_199 : _GEN_974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_976 = 8'hc8 == _match_key_qbytes_0_T_1 ? phv_data_200 : _GEN_975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_977 = 8'hc9 == _match_key_qbytes_0_T_1 ? phv_data_201 : _GEN_976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_978 = 8'hca == _match_key_qbytes_0_T_1 ? phv_data_202 : _GEN_977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_979 = 8'hcb == _match_key_qbytes_0_T_1 ? phv_data_203 : _GEN_978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_980 = 8'hcc == _match_key_qbytes_0_T_1 ? phv_data_204 : _GEN_979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_981 = 8'hcd == _match_key_qbytes_0_T_1 ? phv_data_205 : _GEN_980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_982 = 8'hce == _match_key_qbytes_0_T_1 ? phv_data_206 : _GEN_981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_983 = 8'hcf == _match_key_qbytes_0_T_1 ? phv_data_207 : _GEN_982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_984 = 8'hd0 == _match_key_qbytes_0_T_1 ? phv_data_208 : _GEN_983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_985 = 8'hd1 == _match_key_qbytes_0_T_1 ? phv_data_209 : _GEN_984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_986 = 8'hd2 == _match_key_qbytes_0_T_1 ? phv_data_210 : _GEN_985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_987 = 8'hd3 == _match_key_qbytes_0_T_1 ? phv_data_211 : _GEN_986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_988 = 8'hd4 == _match_key_qbytes_0_T_1 ? phv_data_212 : _GEN_987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_989 = 8'hd5 == _match_key_qbytes_0_T_1 ? phv_data_213 : _GEN_988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_990 = 8'hd6 == _match_key_qbytes_0_T_1 ? phv_data_214 : _GEN_989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_991 = 8'hd7 == _match_key_qbytes_0_T_1 ? phv_data_215 : _GEN_990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_992 = 8'hd8 == _match_key_qbytes_0_T_1 ? phv_data_216 : _GEN_991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_993 = 8'hd9 == _match_key_qbytes_0_T_1 ? phv_data_217 : _GEN_992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_994 = 8'hda == _match_key_qbytes_0_T_1 ? phv_data_218 : _GEN_993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_995 = 8'hdb == _match_key_qbytes_0_T_1 ? phv_data_219 : _GEN_994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_996 = 8'hdc == _match_key_qbytes_0_T_1 ? phv_data_220 : _GEN_995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_997 = 8'hdd == _match_key_qbytes_0_T_1 ? phv_data_221 : _GEN_996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_998 = 8'hde == _match_key_qbytes_0_T_1 ? phv_data_222 : _GEN_997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_999 = 8'hdf == _match_key_qbytes_0_T_1 ? phv_data_223 : _GEN_998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1000 = 8'he0 == _match_key_qbytes_0_T_1 ? phv_data_224 : _GEN_999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1001 = 8'he1 == _match_key_qbytes_0_T_1 ? phv_data_225 : _GEN_1000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1002 = 8'he2 == _match_key_qbytes_0_T_1 ? phv_data_226 : _GEN_1001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1003 = 8'he3 == _match_key_qbytes_0_T_1 ? phv_data_227 : _GEN_1002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1004 = 8'he4 == _match_key_qbytes_0_T_1 ? phv_data_228 : _GEN_1003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1005 = 8'he5 == _match_key_qbytes_0_T_1 ? phv_data_229 : _GEN_1004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1006 = 8'he6 == _match_key_qbytes_0_T_1 ? phv_data_230 : _GEN_1005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1007 = 8'he7 == _match_key_qbytes_0_T_1 ? phv_data_231 : _GEN_1006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1008 = 8'he8 == _match_key_qbytes_0_T_1 ? phv_data_232 : _GEN_1007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1009 = 8'he9 == _match_key_qbytes_0_T_1 ? phv_data_233 : _GEN_1008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1010 = 8'hea == _match_key_qbytes_0_T_1 ? phv_data_234 : _GEN_1009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1011 = 8'heb == _match_key_qbytes_0_T_1 ? phv_data_235 : _GEN_1010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1012 = 8'hec == _match_key_qbytes_0_T_1 ? phv_data_236 : _GEN_1011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1013 = 8'hed == _match_key_qbytes_0_T_1 ? phv_data_237 : _GEN_1012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1014 = 8'hee == _match_key_qbytes_0_T_1 ? phv_data_238 : _GEN_1013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1015 = 8'hef == _match_key_qbytes_0_T_1 ? phv_data_239 : _GEN_1014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1016 = 8'hf0 == _match_key_qbytes_0_T_1 ? phv_data_240 : _GEN_1015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1017 = 8'hf1 == _match_key_qbytes_0_T_1 ? phv_data_241 : _GEN_1016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1018 = 8'hf2 == _match_key_qbytes_0_T_1 ? phv_data_242 : _GEN_1017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1019 = 8'hf3 == _match_key_qbytes_0_T_1 ? phv_data_243 : _GEN_1018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1020 = 8'hf4 == _match_key_qbytes_0_T_1 ? phv_data_244 : _GEN_1019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1021 = 8'hf5 == _match_key_qbytes_0_T_1 ? phv_data_245 : _GEN_1020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1022 = 8'hf6 == _match_key_qbytes_0_T_1 ? phv_data_246 : _GEN_1021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1023 = 8'hf7 == _match_key_qbytes_0_T_1 ? phv_data_247 : _GEN_1022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1024 = 8'hf8 == _match_key_qbytes_0_T_1 ? phv_data_248 : _GEN_1023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1025 = 8'hf9 == _match_key_qbytes_0_T_1 ? phv_data_249 : _GEN_1024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1026 = 8'hfa == _match_key_qbytes_0_T_1 ? phv_data_250 : _GEN_1025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1027 = 8'hfb == _match_key_qbytes_0_T_1 ? phv_data_251 : _GEN_1026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1028 = 8'hfc == _match_key_qbytes_0_T_1 ? phv_data_252 : _GEN_1027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1029 = 8'hfd == _match_key_qbytes_0_T_1 ? phv_data_253 : _GEN_1028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1030 = 8'hfe == _match_key_qbytes_0_T_1 ? phv_data_254 : _GEN_1029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1031 = 8'hff == _match_key_qbytes_0_T_1 ? phv_data_255 : _GEN_1030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_0_T_3 = {_GEN_775,_GEN_1031,_GEN_263,_GEN_519}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_0 = local_offset < end_offset ? _match_key_qbytes_0_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_1 = 8'h4 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_1_hi = local_offset_1[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_1_T = {match_key_qbytes_1_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_1_T_1 = {match_key_qbytes_1_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_1_T_2 = {match_key_qbytes_1_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1034 = 8'h1 == _match_key_qbytes_1_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1035 = 8'h2 == _match_key_qbytes_1_T_2 ? phv_data_2 : _GEN_1034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1036 = 8'h3 == _match_key_qbytes_1_T_2 ? phv_data_3 : _GEN_1035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1037 = 8'h4 == _match_key_qbytes_1_T_2 ? phv_data_4 : _GEN_1036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1038 = 8'h5 == _match_key_qbytes_1_T_2 ? phv_data_5 : _GEN_1037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1039 = 8'h6 == _match_key_qbytes_1_T_2 ? phv_data_6 : _GEN_1038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1040 = 8'h7 == _match_key_qbytes_1_T_2 ? phv_data_7 : _GEN_1039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1041 = 8'h8 == _match_key_qbytes_1_T_2 ? phv_data_8 : _GEN_1040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1042 = 8'h9 == _match_key_qbytes_1_T_2 ? phv_data_9 : _GEN_1041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1043 = 8'ha == _match_key_qbytes_1_T_2 ? phv_data_10 : _GEN_1042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1044 = 8'hb == _match_key_qbytes_1_T_2 ? phv_data_11 : _GEN_1043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1045 = 8'hc == _match_key_qbytes_1_T_2 ? phv_data_12 : _GEN_1044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1046 = 8'hd == _match_key_qbytes_1_T_2 ? phv_data_13 : _GEN_1045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1047 = 8'he == _match_key_qbytes_1_T_2 ? phv_data_14 : _GEN_1046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1048 = 8'hf == _match_key_qbytes_1_T_2 ? phv_data_15 : _GEN_1047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1049 = 8'h10 == _match_key_qbytes_1_T_2 ? phv_data_16 : _GEN_1048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1050 = 8'h11 == _match_key_qbytes_1_T_2 ? phv_data_17 : _GEN_1049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1051 = 8'h12 == _match_key_qbytes_1_T_2 ? phv_data_18 : _GEN_1050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1052 = 8'h13 == _match_key_qbytes_1_T_2 ? phv_data_19 : _GEN_1051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1053 = 8'h14 == _match_key_qbytes_1_T_2 ? phv_data_20 : _GEN_1052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1054 = 8'h15 == _match_key_qbytes_1_T_2 ? phv_data_21 : _GEN_1053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1055 = 8'h16 == _match_key_qbytes_1_T_2 ? phv_data_22 : _GEN_1054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1056 = 8'h17 == _match_key_qbytes_1_T_2 ? phv_data_23 : _GEN_1055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1057 = 8'h18 == _match_key_qbytes_1_T_2 ? phv_data_24 : _GEN_1056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1058 = 8'h19 == _match_key_qbytes_1_T_2 ? phv_data_25 : _GEN_1057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1059 = 8'h1a == _match_key_qbytes_1_T_2 ? phv_data_26 : _GEN_1058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1060 = 8'h1b == _match_key_qbytes_1_T_2 ? phv_data_27 : _GEN_1059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1061 = 8'h1c == _match_key_qbytes_1_T_2 ? phv_data_28 : _GEN_1060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1062 = 8'h1d == _match_key_qbytes_1_T_2 ? phv_data_29 : _GEN_1061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1063 = 8'h1e == _match_key_qbytes_1_T_2 ? phv_data_30 : _GEN_1062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1064 = 8'h1f == _match_key_qbytes_1_T_2 ? phv_data_31 : _GEN_1063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1065 = 8'h20 == _match_key_qbytes_1_T_2 ? phv_data_32 : _GEN_1064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1066 = 8'h21 == _match_key_qbytes_1_T_2 ? phv_data_33 : _GEN_1065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1067 = 8'h22 == _match_key_qbytes_1_T_2 ? phv_data_34 : _GEN_1066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1068 = 8'h23 == _match_key_qbytes_1_T_2 ? phv_data_35 : _GEN_1067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1069 = 8'h24 == _match_key_qbytes_1_T_2 ? phv_data_36 : _GEN_1068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1070 = 8'h25 == _match_key_qbytes_1_T_2 ? phv_data_37 : _GEN_1069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1071 = 8'h26 == _match_key_qbytes_1_T_2 ? phv_data_38 : _GEN_1070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1072 = 8'h27 == _match_key_qbytes_1_T_2 ? phv_data_39 : _GEN_1071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1073 = 8'h28 == _match_key_qbytes_1_T_2 ? phv_data_40 : _GEN_1072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1074 = 8'h29 == _match_key_qbytes_1_T_2 ? phv_data_41 : _GEN_1073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1075 = 8'h2a == _match_key_qbytes_1_T_2 ? phv_data_42 : _GEN_1074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1076 = 8'h2b == _match_key_qbytes_1_T_2 ? phv_data_43 : _GEN_1075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1077 = 8'h2c == _match_key_qbytes_1_T_2 ? phv_data_44 : _GEN_1076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1078 = 8'h2d == _match_key_qbytes_1_T_2 ? phv_data_45 : _GEN_1077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1079 = 8'h2e == _match_key_qbytes_1_T_2 ? phv_data_46 : _GEN_1078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1080 = 8'h2f == _match_key_qbytes_1_T_2 ? phv_data_47 : _GEN_1079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1081 = 8'h30 == _match_key_qbytes_1_T_2 ? phv_data_48 : _GEN_1080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1082 = 8'h31 == _match_key_qbytes_1_T_2 ? phv_data_49 : _GEN_1081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1083 = 8'h32 == _match_key_qbytes_1_T_2 ? phv_data_50 : _GEN_1082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1084 = 8'h33 == _match_key_qbytes_1_T_2 ? phv_data_51 : _GEN_1083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1085 = 8'h34 == _match_key_qbytes_1_T_2 ? phv_data_52 : _GEN_1084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1086 = 8'h35 == _match_key_qbytes_1_T_2 ? phv_data_53 : _GEN_1085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1087 = 8'h36 == _match_key_qbytes_1_T_2 ? phv_data_54 : _GEN_1086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1088 = 8'h37 == _match_key_qbytes_1_T_2 ? phv_data_55 : _GEN_1087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1089 = 8'h38 == _match_key_qbytes_1_T_2 ? phv_data_56 : _GEN_1088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1090 = 8'h39 == _match_key_qbytes_1_T_2 ? phv_data_57 : _GEN_1089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1091 = 8'h3a == _match_key_qbytes_1_T_2 ? phv_data_58 : _GEN_1090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1092 = 8'h3b == _match_key_qbytes_1_T_2 ? phv_data_59 : _GEN_1091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1093 = 8'h3c == _match_key_qbytes_1_T_2 ? phv_data_60 : _GEN_1092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1094 = 8'h3d == _match_key_qbytes_1_T_2 ? phv_data_61 : _GEN_1093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1095 = 8'h3e == _match_key_qbytes_1_T_2 ? phv_data_62 : _GEN_1094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1096 = 8'h3f == _match_key_qbytes_1_T_2 ? phv_data_63 : _GEN_1095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1097 = 8'h40 == _match_key_qbytes_1_T_2 ? phv_data_64 : _GEN_1096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1098 = 8'h41 == _match_key_qbytes_1_T_2 ? phv_data_65 : _GEN_1097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1099 = 8'h42 == _match_key_qbytes_1_T_2 ? phv_data_66 : _GEN_1098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1100 = 8'h43 == _match_key_qbytes_1_T_2 ? phv_data_67 : _GEN_1099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1101 = 8'h44 == _match_key_qbytes_1_T_2 ? phv_data_68 : _GEN_1100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1102 = 8'h45 == _match_key_qbytes_1_T_2 ? phv_data_69 : _GEN_1101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1103 = 8'h46 == _match_key_qbytes_1_T_2 ? phv_data_70 : _GEN_1102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1104 = 8'h47 == _match_key_qbytes_1_T_2 ? phv_data_71 : _GEN_1103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1105 = 8'h48 == _match_key_qbytes_1_T_2 ? phv_data_72 : _GEN_1104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1106 = 8'h49 == _match_key_qbytes_1_T_2 ? phv_data_73 : _GEN_1105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1107 = 8'h4a == _match_key_qbytes_1_T_2 ? phv_data_74 : _GEN_1106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1108 = 8'h4b == _match_key_qbytes_1_T_2 ? phv_data_75 : _GEN_1107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1109 = 8'h4c == _match_key_qbytes_1_T_2 ? phv_data_76 : _GEN_1108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1110 = 8'h4d == _match_key_qbytes_1_T_2 ? phv_data_77 : _GEN_1109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1111 = 8'h4e == _match_key_qbytes_1_T_2 ? phv_data_78 : _GEN_1110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1112 = 8'h4f == _match_key_qbytes_1_T_2 ? phv_data_79 : _GEN_1111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1113 = 8'h50 == _match_key_qbytes_1_T_2 ? phv_data_80 : _GEN_1112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1114 = 8'h51 == _match_key_qbytes_1_T_2 ? phv_data_81 : _GEN_1113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1115 = 8'h52 == _match_key_qbytes_1_T_2 ? phv_data_82 : _GEN_1114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1116 = 8'h53 == _match_key_qbytes_1_T_2 ? phv_data_83 : _GEN_1115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1117 = 8'h54 == _match_key_qbytes_1_T_2 ? phv_data_84 : _GEN_1116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1118 = 8'h55 == _match_key_qbytes_1_T_2 ? phv_data_85 : _GEN_1117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1119 = 8'h56 == _match_key_qbytes_1_T_2 ? phv_data_86 : _GEN_1118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1120 = 8'h57 == _match_key_qbytes_1_T_2 ? phv_data_87 : _GEN_1119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1121 = 8'h58 == _match_key_qbytes_1_T_2 ? phv_data_88 : _GEN_1120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1122 = 8'h59 == _match_key_qbytes_1_T_2 ? phv_data_89 : _GEN_1121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1123 = 8'h5a == _match_key_qbytes_1_T_2 ? phv_data_90 : _GEN_1122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1124 = 8'h5b == _match_key_qbytes_1_T_2 ? phv_data_91 : _GEN_1123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1125 = 8'h5c == _match_key_qbytes_1_T_2 ? phv_data_92 : _GEN_1124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1126 = 8'h5d == _match_key_qbytes_1_T_2 ? phv_data_93 : _GEN_1125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1127 = 8'h5e == _match_key_qbytes_1_T_2 ? phv_data_94 : _GEN_1126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1128 = 8'h5f == _match_key_qbytes_1_T_2 ? phv_data_95 : _GEN_1127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1129 = 8'h60 == _match_key_qbytes_1_T_2 ? phv_data_96 : _GEN_1128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1130 = 8'h61 == _match_key_qbytes_1_T_2 ? phv_data_97 : _GEN_1129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1131 = 8'h62 == _match_key_qbytes_1_T_2 ? phv_data_98 : _GEN_1130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1132 = 8'h63 == _match_key_qbytes_1_T_2 ? phv_data_99 : _GEN_1131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1133 = 8'h64 == _match_key_qbytes_1_T_2 ? phv_data_100 : _GEN_1132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1134 = 8'h65 == _match_key_qbytes_1_T_2 ? phv_data_101 : _GEN_1133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1135 = 8'h66 == _match_key_qbytes_1_T_2 ? phv_data_102 : _GEN_1134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1136 = 8'h67 == _match_key_qbytes_1_T_2 ? phv_data_103 : _GEN_1135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1137 = 8'h68 == _match_key_qbytes_1_T_2 ? phv_data_104 : _GEN_1136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1138 = 8'h69 == _match_key_qbytes_1_T_2 ? phv_data_105 : _GEN_1137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1139 = 8'h6a == _match_key_qbytes_1_T_2 ? phv_data_106 : _GEN_1138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1140 = 8'h6b == _match_key_qbytes_1_T_2 ? phv_data_107 : _GEN_1139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1141 = 8'h6c == _match_key_qbytes_1_T_2 ? phv_data_108 : _GEN_1140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1142 = 8'h6d == _match_key_qbytes_1_T_2 ? phv_data_109 : _GEN_1141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1143 = 8'h6e == _match_key_qbytes_1_T_2 ? phv_data_110 : _GEN_1142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1144 = 8'h6f == _match_key_qbytes_1_T_2 ? phv_data_111 : _GEN_1143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1145 = 8'h70 == _match_key_qbytes_1_T_2 ? phv_data_112 : _GEN_1144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1146 = 8'h71 == _match_key_qbytes_1_T_2 ? phv_data_113 : _GEN_1145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1147 = 8'h72 == _match_key_qbytes_1_T_2 ? phv_data_114 : _GEN_1146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1148 = 8'h73 == _match_key_qbytes_1_T_2 ? phv_data_115 : _GEN_1147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1149 = 8'h74 == _match_key_qbytes_1_T_2 ? phv_data_116 : _GEN_1148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1150 = 8'h75 == _match_key_qbytes_1_T_2 ? phv_data_117 : _GEN_1149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1151 = 8'h76 == _match_key_qbytes_1_T_2 ? phv_data_118 : _GEN_1150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1152 = 8'h77 == _match_key_qbytes_1_T_2 ? phv_data_119 : _GEN_1151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1153 = 8'h78 == _match_key_qbytes_1_T_2 ? phv_data_120 : _GEN_1152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1154 = 8'h79 == _match_key_qbytes_1_T_2 ? phv_data_121 : _GEN_1153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1155 = 8'h7a == _match_key_qbytes_1_T_2 ? phv_data_122 : _GEN_1154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1156 = 8'h7b == _match_key_qbytes_1_T_2 ? phv_data_123 : _GEN_1155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1157 = 8'h7c == _match_key_qbytes_1_T_2 ? phv_data_124 : _GEN_1156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1158 = 8'h7d == _match_key_qbytes_1_T_2 ? phv_data_125 : _GEN_1157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1159 = 8'h7e == _match_key_qbytes_1_T_2 ? phv_data_126 : _GEN_1158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1160 = 8'h7f == _match_key_qbytes_1_T_2 ? phv_data_127 : _GEN_1159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1161 = 8'h80 == _match_key_qbytes_1_T_2 ? phv_data_128 : _GEN_1160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1162 = 8'h81 == _match_key_qbytes_1_T_2 ? phv_data_129 : _GEN_1161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1163 = 8'h82 == _match_key_qbytes_1_T_2 ? phv_data_130 : _GEN_1162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1164 = 8'h83 == _match_key_qbytes_1_T_2 ? phv_data_131 : _GEN_1163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1165 = 8'h84 == _match_key_qbytes_1_T_2 ? phv_data_132 : _GEN_1164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1166 = 8'h85 == _match_key_qbytes_1_T_2 ? phv_data_133 : _GEN_1165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1167 = 8'h86 == _match_key_qbytes_1_T_2 ? phv_data_134 : _GEN_1166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1168 = 8'h87 == _match_key_qbytes_1_T_2 ? phv_data_135 : _GEN_1167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1169 = 8'h88 == _match_key_qbytes_1_T_2 ? phv_data_136 : _GEN_1168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1170 = 8'h89 == _match_key_qbytes_1_T_2 ? phv_data_137 : _GEN_1169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1171 = 8'h8a == _match_key_qbytes_1_T_2 ? phv_data_138 : _GEN_1170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1172 = 8'h8b == _match_key_qbytes_1_T_2 ? phv_data_139 : _GEN_1171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1173 = 8'h8c == _match_key_qbytes_1_T_2 ? phv_data_140 : _GEN_1172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1174 = 8'h8d == _match_key_qbytes_1_T_2 ? phv_data_141 : _GEN_1173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1175 = 8'h8e == _match_key_qbytes_1_T_2 ? phv_data_142 : _GEN_1174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1176 = 8'h8f == _match_key_qbytes_1_T_2 ? phv_data_143 : _GEN_1175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1177 = 8'h90 == _match_key_qbytes_1_T_2 ? phv_data_144 : _GEN_1176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1178 = 8'h91 == _match_key_qbytes_1_T_2 ? phv_data_145 : _GEN_1177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1179 = 8'h92 == _match_key_qbytes_1_T_2 ? phv_data_146 : _GEN_1178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1180 = 8'h93 == _match_key_qbytes_1_T_2 ? phv_data_147 : _GEN_1179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1181 = 8'h94 == _match_key_qbytes_1_T_2 ? phv_data_148 : _GEN_1180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1182 = 8'h95 == _match_key_qbytes_1_T_2 ? phv_data_149 : _GEN_1181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1183 = 8'h96 == _match_key_qbytes_1_T_2 ? phv_data_150 : _GEN_1182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1184 = 8'h97 == _match_key_qbytes_1_T_2 ? phv_data_151 : _GEN_1183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1185 = 8'h98 == _match_key_qbytes_1_T_2 ? phv_data_152 : _GEN_1184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1186 = 8'h99 == _match_key_qbytes_1_T_2 ? phv_data_153 : _GEN_1185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1187 = 8'h9a == _match_key_qbytes_1_T_2 ? phv_data_154 : _GEN_1186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1188 = 8'h9b == _match_key_qbytes_1_T_2 ? phv_data_155 : _GEN_1187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1189 = 8'h9c == _match_key_qbytes_1_T_2 ? phv_data_156 : _GEN_1188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1190 = 8'h9d == _match_key_qbytes_1_T_2 ? phv_data_157 : _GEN_1189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1191 = 8'h9e == _match_key_qbytes_1_T_2 ? phv_data_158 : _GEN_1190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1192 = 8'h9f == _match_key_qbytes_1_T_2 ? phv_data_159 : _GEN_1191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1193 = 8'ha0 == _match_key_qbytes_1_T_2 ? phv_data_160 : _GEN_1192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1194 = 8'ha1 == _match_key_qbytes_1_T_2 ? phv_data_161 : _GEN_1193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1195 = 8'ha2 == _match_key_qbytes_1_T_2 ? phv_data_162 : _GEN_1194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1196 = 8'ha3 == _match_key_qbytes_1_T_2 ? phv_data_163 : _GEN_1195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1197 = 8'ha4 == _match_key_qbytes_1_T_2 ? phv_data_164 : _GEN_1196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1198 = 8'ha5 == _match_key_qbytes_1_T_2 ? phv_data_165 : _GEN_1197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1199 = 8'ha6 == _match_key_qbytes_1_T_2 ? phv_data_166 : _GEN_1198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1200 = 8'ha7 == _match_key_qbytes_1_T_2 ? phv_data_167 : _GEN_1199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1201 = 8'ha8 == _match_key_qbytes_1_T_2 ? phv_data_168 : _GEN_1200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1202 = 8'ha9 == _match_key_qbytes_1_T_2 ? phv_data_169 : _GEN_1201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1203 = 8'haa == _match_key_qbytes_1_T_2 ? phv_data_170 : _GEN_1202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1204 = 8'hab == _match_key_qbytes_1_T_2 ? phv_data_171 : _GEN_1203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1205 = 8'hac == _match_key_qbytes_1_T_2 ? phv_data_172 : _GEN_1204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1206 = 8'had == _match_key_qbytes_1_T_2 ? phv_data_173 : _GEN_1205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1207 = 8'hae == _match_key_qbytes_1_T_2 ? phv_data_174 : _GEN_1206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1208 = 8'haf == _match_key_qbytes_1_T_2 ? phv_data_175 : _GEN_1207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1209 = 8'hb0 == _match_key_qbytes_1_T_2 ? phv_data_176 : _GEN_1208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1210 = 8'hb1 == _match_key_qbytes_1_T_2 ? phv_data_177 : _GEN_1209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1211 = 8'hb2 == _match_key_qbytes_1_T_2 ? phv_data_178 : _GEN_1210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1212 = 8'hb3 == _match_key_qbytes_1_T_2 ? phv_data_179 : _GEN_1211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1213 = 8'hb4 == _match_key_qbytes_1_T_2 ? phv_data_180 : _GEN_1212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1214 = 8'hb5 == _match_key_qbytes_1_T_2 ? phv_data_181 : _GEN_1213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1215 = 8'hb6 == _match_key_qbytes_1_T_2 ? phv_data_182 : _GEN_1214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1216 = 8'hb7 == _match_key_qbytes_1_T_2 ? phv_data_183 : _GEN_1215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1217 = 8'hb8 == _match_key_qbytes_1_T_2 ? phv_data_184 : _GEN_1216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1218 = 8'hb9 == _match_key_qbytes_1_T_2 ? phv_data_185 : _GEN_1217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1219 = 8'hba == _match_key_qbytes_1_T_2 ? phv_data_186 : _GEN_1218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1220 = 8'hbb == _match_key_qbytes_1_T_2 ? phv_data_187 : _GEN_1219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1221 = 8'hbc == _match_key_qbytes_1_T_2 ? phv_data_188 : _GEN_1220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1222 = 8'hbd == _match_key_qbytes_1_T_2 ? phv_data_189 : _GEN_1221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1223 = 8'hbe == _match_key_qbytes_1_T_2 ? phv_data_190 : _GEN_1222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1224 = 8'hbf == _match_key_qbytes_1_T_2 ? phv_data_191 : _GEN_1223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1225 = 8'hc0 == _match_key_qbytes_1_T_2 ? phv_data_192 : _GEN_1224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1226 = 8'hc1 == _match_key_qbytes_1_T_2 ? phv_data_193 : _GEN_1225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1227 = 8'hc2 == _match_key_qbytes_1_T_2 ? phv_data_194 : _GEN_1226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1228 = 8'hc3 == _match_key_qbytes_1_T_2 ? phv_data_195 : _GEN_1227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1229 = 8'hc4 == _match_key_qbytes_1_T_2 ? phv_data_196 : _GEN_1228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1230 = 8'hc5 == _match_key_qbytes_1_T_2 ? phv_data_197 : _GEN_1229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1231 = 8'hc6 == _match_key_qbytes_1_T_2 ? phv_data_198 : _GEN_1230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1232 = 8'hc7 == _match_key_qbytes_1_T_2 ? phv_data_199 : _GEN_1231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1233 = 8'hc8 == _match_key_qbytes_1_T_2 ? phv_data_200 : _GEN_1232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1234 = 8'hc9 == _match_key_qbytes_1_T_2 ? phv_data_201 : _GEN_1233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1235 = 8'hca == _match_key_qbytes_1_T_2 ? phv_data_202 : _GEN_1234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1236 = 8'hcb == _match_key_qbytes_1_T_2 ? phv_data_203 : _GEN_1235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1237 = 8'hcc == _match_key_qbytes_1_T_2 ? phv_data_204 : _GEN_1236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1238 = 8'hcd == _match_key_qbytes_1_T_2 ? phv_data_205 : _GEN_1237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1239 = 8'hce == _match_key_qbytes_1_T_2 ? phv_data_206 : _GEN_1238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1240 = 8'hcf == _match_key_qbytes_1_T_2 ? phv_data_207 : _GEN_1239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1241 = 8'hd0 == _match_key_qbytes_1_T_2 ? phv_data_208 : _GEN_1240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1242 = 8'hd1 == _match_key_qbytes_1_T_2 ? phv_data_209 : _GEN_1241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1243 = 8'hd2 == _match_key_qbytes_1_T_2 ? phv_data_210 : _GEN_1242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1244 = 8'hd3 == _match_key_qbytes_1_T_2 ? phv_data_211 : _GEN_1243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1245 = 8'hd4 == _match_key_qbytes_1_T_2 ? phv_data_212 : _GEN_1244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1246 = 8'hd5 == _match_key_qbytes_1_T_2 ? phv_data_213 : _GEN_1245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1247 = 8'hd6 == _match_key_qbytes_1_T_2 ? phv_data_214 : _GEN_1246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1248 = 8'hd7 == _match_key_qbytes_1_T_2 ? phv_data_215 : _GEN_1247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1249 = 8'hd8 == _match_key_qbytes_1_T_2 ? phv_data_216 : _GEN_1248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1250 = 8'hd9 == _match_key_qbytes_1_T_2 ? phv_data_217 : _GEN_1249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1251 = 8'hda == _match_key_qbytes_1_T_2 ? phv_data_218 : _GEN_1250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1252 = 8'hdb == _match_key_qbytes_1_T_2 ? phv_data_219 : _GEN_1251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1253 = 8'hdc == _match_key_qbytes_1_T_2 ? phv_data_220 : _GEN_1252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1254 = 8'hdd == _match_key_qbytes_1_T_2 ? phv_data_221 : _GEN_1253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1255 = 8'hde == _match_key_qbytes_1_T_2 ? phv_data_222 : _GEN_1254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1256 = 8'hdf == _match_key_qbytes_1_T_2 ? phv_data_223 : _GEN_1255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1257 = 8'he0 == _match_key_qbytes_1_T_2 ? phv_data_224 : _GEN_1256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1258 = 8'he1 == _match_key_qbytes_1_T_2 ? phv_data_225 : _GEN_1257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1259 = 8'he2 == _match_key_qbytes_1_T_2 ? phv_data_226 : _GEN_1258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1260 = 8'he3 == _match_key_qbytes_1_T_2 ? phv_data_227 : _GEN_1259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1261 = 8'he4 == _match_key_qbytes_1_T_2 ? phv_data_228 : _GEN_1260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1262 = 8'he5 == _match_key_qbytes_1_T_2 ? phv_data_229 : _GEN_1261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1263 = 8'he6 == _match_key_qbytes_1_T_2 ? phv_data_230 : _GEN_1262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1264 = 8'he7 == _match_key_qbytes_1_T_2 ? phv_data_231 : _GEN_1263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1265 = 8'he8 == _match_key_qbytes_1_T_2 ? phv_data_232 : _GEN_1264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1266 = 8'he9 == _match_key_qbytes_1_T_2 ? phv_data_233 : _GEN_1265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1267 = 8'hea == _match_key_qbytes_1_T_2 ? phv_data_234 : _GEN_1266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1268 = 8'heb == _match_key_qbytes_1_T_2 ? phv_data_235 : _GEN_1267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1269 = 8'hec == _match_key_qbytes_1_T_2 ? phv_data_236 : _GEN_1268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1270 = 8'hed == _match_key_qbytes_1_T_2 ? phv_data_237 : _GEN_1269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1271 = 8'hee == _match_key_qbytes_1_T_2 ? phv_data_238 : _GEN_1270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1272 = 8'hef == _match_key_qbytes_1_T_2 ? phv_data_239 : _GEN_1271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1273 = 8'hf0 == _match_key_qbytes_1_T_2 ? phv_data_240 : _GEN_1272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1274 = 8'hf1 == _match_key_qbytes_1_T_2 ? phv_data_241 : _GEN_1273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1275 = 8'hf2 == _match_key_qbytes_1_T_2 ? phv_data_242 : _GEN_1274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1276 = 8'hf3 == _match_key_qbytes_1_T_2 ? phv_data_243 : _GEN_1275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1277 = 8'hf4 == _match_key_qbytes_1_T_2 ? phv_data_244 : _GEN_1276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1278 = 8'hf5 == _match_key_qbytes_1_T_2 ? phv_data_245 : _GEN_1277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1279 = 8'hf6 == _match_key_qbytes_1_T_2 ? phv_data_246 : _GEN_1278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1280 = 8'hf7 == _match_key_qbytes_1_T_2 ? phv_data_247 : _GEN_1279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1281 = 8'hf8 == _match_key_qbytes_1_T_2 ? phv_data_248 : _GEN_1280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1282 = 8'hf9 == _match_key_qbytes_1_T_2 ? phv_data_249 : _GEN_1281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1283 = 8'hfa == _match_key_qbytes_1_T_2 ? phv_data_250 : _GEN_1282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1284 = 8'hfb == _match_key_qbytes_1_T_2 ? phv_data_251 : _GEN_1283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1285 = 8'hfc == _match_key_qbytes_1_T_2 ? phv_data_252 : _GEN_1284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1286 = 8'hfd == _match_key_qbytes_1_T_2 ? phv_data_253 : _GEN_1285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1287 = 8'hfe == _match_key_qbytes_1_T_2 ? phv_data_254 : _GEN_1286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1288 = 8'hff == _match_key_qbytes_1_T_2 ? phv_data_255 : _GEN_1287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1290 = 8'h1 == local_offset_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1291 = 8'h2 == local_offset_1 ? phv_data_2 : _GEN_1290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1292 = 8'h3 == local_offset_1 ? phv_data_3 : _GEN_1291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1293 = 8'h4 == local_offset_1 ? phv_data_4 : _GEN_1292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1294 = 8'h5 == local_offset_1 ? phv_data_5 : _GEN_1293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1295 = 8'h6 == local_offset_1 ? phv_data_6 : _GEN_1294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1296 = 8'h7 == local_offset_1 ? phv_data_7 : _GEN_1295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1297 = 8'h8 == local_offset_1 ? phv_data_8 : _GEN_1296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1298 = 8'h9 == local_offset_1 ? phv_data_9 : _GEN_1297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1299 = 8'ha == local_offset_1 ? phv_data_10 : _GEN_1298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1300 = 8'hb == local_offset_1 ? phv_data_11 : _GEN_1299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1301 = 8'hc == local_offset_1 ? phv_data_12 : _GEN_1300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1302 = 8'hd == local_offset_1 ? phv_data_13 : _GEN_1301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1303 = 8'he == local_offset_1 ? phv_data_14 : _GEN_1302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1304 = 8'hf == local_offset_1 ? phv_data_15 : _GEN_1303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1305 = 8'h10 == local_offset_1 ? phv_data_16 : _GEN_1304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1306 = 8'h11 == local_offset_1 ? phv_data_17 : _GEN_1305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1307 = 8'h12 == local_offset_1 ? phv_data_18 : _GEN_1306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1308 = 8'h13 == local_offset_1 ? phv_data_19 : _GEN_1307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1309 = 8'h14 == local_offset_1 ? phv_data_20 : _GEN_1308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1310 = 8'h15 == local_offset_1 ? phv_data_21 : _GEN_1309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1311 = 8'h16 == local_offset_1 ? phv_data_22 : _GEN_1310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1312 = 8'h17 == local_offset_1 ? phv_data_23 : _GEN_1311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1313 = 8'h18 == local_offset_1 ? phv_data_24 : _GEN_1312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1314 = 8'h19 == local_offset_1 ? phv_data_25 : _GEN_1313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1315 = 8'h1a == local_offset_1 ? phv_data_26 : _GEN_1314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1316 = 8'h1b == local_offset_1 ? phv_data_27 : _GEN_1315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1317 = 8'h1c == local_offset_1 ? phv_data_28 : _GEN_1316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1318 = 8'h1d == local_offset_1 ? phv_data_29 : _GEN_1317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1319 = 8'h1e == local_offset_1 ? phv_data_30 : _GEN_1318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1320 = 8'h1f == local_offset_1 ? phv_data_31 : _GEN_1319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1321 = 8'h20 == local_offset_1 ? phv_data_32 : _GEN_1320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1322 = 8'h21 == local_offset_1 ? phv_data_33 : _GEN_1321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1323 = 8'h22 == local_offset_1 ? phv_data_34 : _GEN_1322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1324 = 8'h23 == local_offset_1 ? phv_data_35 : _GEN_1323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1325 = 8'h24 == local_offset_1 ? phv_data_36 : _GEN_1324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1326 = 8'h25 == local_offset_1 ? phv_data_37 : _GEN_1325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1327 = 8'h26 == local_offset_1 ? phv_data_38 : _GEN_1326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1328 = 8'h27 == local_offset_1 ? phv_data_39 : _GEN_1327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1329 = 8'h28 == local_offset_1 ? phv_data_40 : _GEN_1328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1330 = 8'h29 == local_offset_1 ? phv_data_41 : _GEN_1329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1331 = 8'h2a == local_offset_1 ? phv_data_42 : _GEN_1330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1332 = 8'h2b == local_offset_1 ? phv_data_43 : _GEN_1331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1333 = 8'h2c == local_offset_1 ? phv_data_44 : _GEN_1332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1334 = 8'h2d == local_offset_1 ? phv_data_45 : _GEN_1333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1335 = 8'h2e == local_offset_1 ? phv_data_46 : _GEN_1334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1336 = 8'h2f == local_offset_1 ? phv_data_47 : _GEN_1335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1337 = 8'h30 == local_offset_1 ? phv_data_48 : _GEN_1336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1338 = 8'h31 == local_offset_1 ? phv_data_49 : _GEN_1337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1339 = 8'h32 == local_offset_1 ? phv_data_50 : _GEN_1338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1340 = 8'h33 == local_offset_1 ? phv_data_51 : _GEN_1339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1341 = 8'h34 == local_offset_1 ? phv_data_52 : _GEN_1340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1342 = 8'h35 == local_offset_1 ? phv_data_53 : _GEN_1341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1343 = 8'h36 == local_offset_1 ? phv_data_54 : _GEN_1342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1344 = 8'h37 == local_offset_1 ? phv_data_55 : _GEN_1343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1345 = 8'h38 == local_offset_1 ? phv_data_56 : _GEN_1344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1346 = 8'h39 == local_offset_1 ? phv_data_57 : _GEN_1345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1347 = 8'h3a == local_offset_1 ? phv_data_58 : _GEN_1346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1348 = 8'h3b == local_offset_1 ? phv_data_59 : _GEN_1347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1349 = 8'h3c == local_offset_1 ? phv_data_60 : _GEN_1348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1350 = 8'h3d == local_offset_1 ? phv_data_61 : _GEN_1349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1351 = 8'h3e == local_offset_1 ? phv_data_62 : _GEN_1350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1352 = 8'h3f == local_offset_1 ? phv_data_63 : _GEN_1351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1353 = 8'h40 == local_offset_1 ? phv_data_64 : _GEN_1352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1354 = 8'h41 == local_offset_1 ? phv_data_65 : _GEN_1353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1355 = 8'h42 == local_offset_1 ? phv_data_66 : _GEN_1354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1356 = 8'h43 == local_offset_1 ? phv_data_67 : _GEN_1355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1357 = 8'h44 == local_offset_1 ? phv_data_68 : _GEN_1356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1358 = 8'h45 == local_offset_1 ? phv_data_69 : _GEN_1357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1359 = 8'h46 == local_offset_1 ? phv_data_70 : _GEN_1358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1360 = 8'h47 == local_offset_1 ? phv_data_71 : _GEN_1359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1361 = 8'h48 == local_offset_1 ? phv_data_72 : _GEN_1360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1362 = 8'h49 == local_offset_1 ? phv_data_73 : _GEN_1361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1363 = 8'h4a == local_offset_1 ? phv_data_74 : _GEN_1362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1364 = 8'h4b == local_offset_1 ? phv_data_75 : _GEN_1363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1365 = 8'h4c == local_offset_1 ? phv_data_76 : _GEN_1364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1366 = 8'h4d == local_offset_1 ? phv_data_77 : _GEN_1365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1367 = 8'h4e == local_offset_1 ? phv_data_78 : _GEN_1366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1368 = 8'h4f == local_offset_1 ? phv_data_79 : _GEN_1367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1369 = 8'h50 == local_offset_1 ? phv_data_80 : _GEN_1368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1370 = 8'h51 == local_offset_1 ? phv_data_81 : _GEN_1369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1371 = 8'h52 == local_offset_1 ? phv_data_82 : _GEN_1370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1372 = 8'h53 == local_offset_1 ? phv_data_83 : _GEN_1371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1373 = 8'h54 == local_offset_1 ? phv_data_84 : _GEN_1372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1374 = 8'h55 == local_offset_1 ? phv_data_85 : _GEN_1373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1375 = 8'h56 == local_offset_1 ? phv_data_86 : _GEN_1374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1376 = 8'h57 == local_offset_1 ? phv_data_87 : _GEN_1375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1377 = 8'h58 == local_offset_1 ? phv_data_88 : _GEN_1376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1378 = 8'h59 == local_offset_1 ? phv_data_89 : _GEN_1377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1379 = 8'h5a == local_offset_1 ? phv_data_90 : _GEN_1378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1380 = 8'h5b == local_offset_1 ? phv_data_91 : _GEN_1379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1381 = 8'h5c == local_offset_1 ? phv_data_92 : _GEN_1380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1382 = 8'h5d == local_offset_1 ? phv_data_93 : _GEN_1381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1383 = 8'h5e == local_offset_1 ? phv_data_94 : _GEN_1382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1384 = 8'h5f == local_offset_1 ? phv_data_95 : _GEN_1383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1385 = 8'h60 == local_offset_1 ? phv_data_96 : _GEN_1384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1386 = 8'h61 == local_offset_1 ? phv_data_97 : _GEN_1385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1387 = 8'h62 == local_offset_1 ? phv_data_98 : _GEN_1386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1388 = 8'h63 == local_offset_1 ? phv_data_99 : _GEN_1387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1389 = 8'h64 == local_offset_1 ? phv_data_100 : _GEN_1388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1390 = 8'h65 == local_offset_1 ? phv_data_101 : _GEN_1389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1391 = 8'h66 == local_offset_1 ? phv_data_102 : _GEN_1390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1392 = 8'h67 == local_offset_1 ? phv_data_103 : _GEN_1391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1393 = 8'h68 == local_offset_1 ? phv_data_104 : _GEN_1392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1394 = 8'h69 == local_offset_1 ? phv_data_105 : _GEN_1393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1395 = 8'h6a == local_offset_1 ? phv_data_106 : _GEN_1394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1396 = 8'h6b == local_offset_1 ? phv_data_107 : _GEN_1395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1397 = 8'h6c == local_offset_1 ? phv_data_108 : _GEN_1396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1398 = 8'h6d == local_offset_1 ? phv_data_109 : _GEN_1397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1399 = 8'h6e == local_offset_1 ? phv_data_110 : _GEN_1398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1400 = 8'h6f == local_offset_1 ? phv_data_111 : _GEN_1399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1401 = 8'h70 == local_offset_1 ? phv_data_112 : _GEN_1400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1402 = 8'h71 == local_offset_1 ? phv_data_113 : _GEN_1401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1403 = 8'h72 == local_offset_1 ? phv_data_114 : _GEN_1402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1404 = 8'h73 == local_offset_1 ? phv_data_115 : _GEN_1403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1405 = 8'h74 == local_offset_1 ? phv_data_116 : _GEN_1404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1406 = 8'h75 == local_offset_1 ? phv_data_117 : _GEN_1405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1407 = 8'h76 == local_offset_1 ? phv_data_118 : _GEN_1406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1408 = 8'h77 == local_offset_1 ? phv_data_119 : _GEN_1407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1409 = 8'h78 == local_offset_1 ? phv_data_120 : _GEN_1408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1410 = 8'h79 == local_offset_1 ? phv_data_121 : _GEN_1409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1411 = 8'h7a == local_offset_1 ? phv_data_122 : _GEN_1410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1412 = 8'h7b == local_offset_1 ? phv_data_123 : _GEN_1411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1413 = 8'h7c == local_offset_1 ? phv_data_124 : _GEN_1412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1414 = 8'h7d == local_offset_1 ? phv_data_125 : _GEN_1413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1415 = 8'h7e == local_offset_1 ? phv_data_126 : _GEN_1414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1416 = 8'h7f == local_offset_1 ? phv_data_127 : _GEN_1415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1417 = 8'h80 == local_offset_1 ? phv_data_128 : _GEN_1416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1418 = 8'h81 == local_offset_1 ? phv_data_129 : _GEN_1417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1419 = 8'h82 == local_offset_1 ? phv_data_130 : _GEN_1418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1420 = 8'h83 == local_offset_1 ? phv_data_131 : _GEN_1419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1421 = 8'h84 == local_offset_1 ? phv_data_132 : _GEN_1420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1422 = 8'h85 == local_offset_1 ? phv_data_133 : _GEN_1421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1423 = 8'h86 == local_offset_1 ? phv_data_134 : _GEN_1422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1424 = 8'h87 == local_offset_1 ? phv_data_135 : _GEN_1423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1425 = 8'h88 == local_offset_1 ? phv_data_136 : _GEN_1424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1426 = 8'h89 == local_offset_1 ? phv_data_137 : _GEN_1425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1427 = 8'h8a == local_offset_1 ? phv_data_138 : _GEN_1426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1428 = 8'h8b == local_offset_1 ? phv_data_139 : _GEN_1427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1429 = 8'h8c == local_offset_1 ? phv_data_140 : _GEN_1428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1430 = 8'h8d == local_offset_1 ? phv_data_141 : _GEN_1429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1431 = 8'h8e == local_offset_1 ? phv_data_142 : _GEN_1430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1432 = 8'h8f == local_offset_1 ? phv_data_143 : _GEN_1431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1433 = 8'h90 == local_offset_1 ? phv_data_144 : _GEN_1432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1434 = 8'h91 == local_offset_1 ? phv_data_145 : _GEN_1433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1435 = 8'h92 == local_offset_1 ? phv_data_146 : _GEN_1434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1436 = 8'h93 == local_offset_1 ? phv_data_147 : _GEN_1435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1437 = 8'h94 == local_offset_1 ? phv_data_148 : _GEN_1436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1438 = 8'h95 == local_offset_1 ? phv_data_149 : _GEN_1437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1439 = 8'h96 == local_offset_1 ? phv_data_150 : _GEN_1438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1440 = 8'h97 == local_offset_1 ? phv_data_151 : _GEN_1439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1441 = 8'h98 == local_offset_1 ? phv_data_152 : _GEN_1440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1442 = 8'h99 == local_offset_1 ? phv_data_153 : _GEN_1441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1443 = 8'h9a == local_offset_1 ? phv_data_154 : _GEN_1442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1444 = 8'h9b == local_offset_1 ? phv_data_155 : _GEN_1443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1445 = 8'h9c == local_offset_1 ? phv_data_156 : _GEN_1444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1446 = 8'h9d == local_offset_1 ? phv_data_157 : _GEN_1445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1447 = 8'h9e == local_offset_1 ? phv_data_158 : _GEN_1446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1448 = 8'h9f == local_offset_1 ? phv_data_159 : _GEN_1447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1449 = 8'ha0 == local_offset_1 ? phv_data_160 : _GEN_1448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1450 = 8'ha1 == local_offset_1 ? phv_data_161 : _GEN_1449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1451 = 8'ha2 == local_offset_1 ? phv_data_162 : _GEN_1450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1452 = 8'ha3 == local_offset_1 ? phv_data_163 : _GEN_1451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1453 = 8'ha4 == local_offset_1 ? phv_data_164 : _GEN_1452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1454 = 8'ha5 == local_offset_1 ? phv_data_165 : _GEN_1453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1455 = 8'ha6 == local_offset_1 ? phv_data_166 : _GEN_1454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1456 = 8'ha7 == local_offset_1 ? phv_data_167 : _GEN_1455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1457 = 8'ha8 == local_offset_1 ? phv_data_168 : _GEN_1456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1458 = 8'ha9 == local_offset_1 ? phv_data_169 : _GEN_1457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1459 = 8'haa == local_offset_1 ? phv_data_170 : _GEN_1458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1460 = 8'hab == local_offset_1 ? phv_data_171 : _GEN_1459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1461 = 8'hac == local_offset_1 ? phv_data_172 : _GEN_1460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1462 = 8'had == local_offset_1 ? phv_data_173 : _GEN_1461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1463 = 8'hae == local_offset_1 ? phv_data_174 : _GEN_1462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1464 = 8'haf == local_offset_1 ? phv_data_175 : _GEN_1463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1465 = 8'hb0 == local_offset_1 ? phv_data_176 : _GEN_1464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1466 = 8'hb1 == local_offset_1 ? phv_data_177 : _GEN_1465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1467 = 8'hb2 == local_offset_1 ? phv_data_178 : _GEN_1466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1468 = 8'hb3 == local_offset_1 ? phv_data_179 : _GEN_1467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1469 = 8'hb4 == local_offset_1 ? phv_data_180 : _GEN_1468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1470 = 8'hb5 == local_offset_1 ? phv_data_181 : _GEN_1469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1471 = 8'hb6 == local_offset_1 ? phv_data_182 : _GEN_1470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1472 = 8'hb7 == local_offset_1 ? phv_data_183 : _GEN_1471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1473 = 8'hb8 == local_offset_1 ? phv_data_184 : _GEN_1472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1474 = 8'hb9 == local_offset_1 ? phv_data_185 : _GEN_1473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1475 = 8'hba == local_offset_1 ? phv_data_186 : _GEN_1474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1476 = 8'hbb == local_offset_1 ? phv_data_187 : _GEN_1475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1477 = 8'hbc == local_offset_1 ? phv_data_188 : _GEN_1476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1478 = 8'hbd == local_offset_1 ? phv_data_189 : _GEN_1477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1479 = 8'hbe == local_offset_1 ? phv_data_190 : _GEN_1478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1480 = 8'hbf == local_offset_1 ? phv_data_191 : _GEN_1479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1481 = 8'hc0 == local_offset_1 ? phv_data_192 : _GEN_1480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1482 = 8'hc1 == local_offset_1 ? phv_data_193 : _GEN_1481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1483 = 8'hc2 == local_offset_1 ? phv_data_194 : _GEN_1482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1484 = 8'hc3 == local_offset_1 ? phv_data_195 : _GEN_1483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1485 = 8'hc4 == local_offset_1 ? phv_data_196 : _GEN_1484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1486 = 8'hc5 == local_offset_1 ? phv_data_197 : _GEN_1485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1487 = 8'hc6 == local_offset_1 ? phv_data_198 : _GEN_1486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1488 = 8'hc7 == local_offset_1 ? phv_data_199 : _GEN_1487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1489 = 8'hc8 == local_offset_1 ? phv_data_200 : _GEN_1488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1490 = 8'hc9 == local_offset_1 ? phv_data_201 : _GEN_1489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1491 = 8'hca == local_offset_1 ? phv_data_202 : _GEN_1490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1492 = 8'hcb == local_offset_1 ? phv_data_203 : _GEN_1491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1493 = 8'hcc == local_offset_1 ? phv_data_204 : _GEN_1492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1494 = 8'hcd == local_offset_1 ? phv_data_205 : _GEN_1493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1495 = 8'hce == local_offset_1 ? phv_data_206 : _GEN_1494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1496 = 8'hcf == local_offset_1 ? phv_data_207 : _GEN_1495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1497 = 8'hd0 == local_offset_1 ? phv_data_208 : _GEN_1496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1498 = 8'hd1 == local_offset_1 ? phv_data_209 : _GEN_1497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1499 = 8'hd2 == local_offset_1 ? phv_data_210 : _GEN_1498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1500 = 8'hd3 == local_offset_1 ? phv_data_211 : _GEN_1499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1501 = 8'hd4 == local_offset_1 ? phv_data_212 : _GEN_1500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1502 = 8'hd5 == local_offset_1 ? phv_data_213 : _GEN_1501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1503 = 8'hd6 == local_offset_1 ? phv_data_214 : _GEN_1502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1504 = 8'hd7 == local_offset_1 ? phv_data_215 : _GEN_1503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1505 = 8'hd8 == local_offset_1 ? phv_data_216 : _GEN_1504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1506 = 8'hd9 == local_offset_1 ? phv_data_217 : _GEN_1505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1507 = 8'hda == local_offset_1 ? phv_data_218 : _GEN_1506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1508 = 8'hdb == local_offset_1 ? phv_data_219 : _GEN_1507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1509 = 8'hdc == local_offset_1 ? phv_data_220 : _GEN_1508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1510 = 8'hdd == local_offset_1 ? phv_data_221 : _GEN_1509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1511 = 8'hde == local_offset_1 ? phv_data_222 : _GEN_1510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1512 = 8'hdf == local_offset_1 ? phv_data_223 : _GEN_1511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1513 = 8'he0 == local_offset_1 ? phv_data_224 : _GEN_1512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1514 = 8'he1 == local_offset_1 ? phv_data_225 : _GEN_1513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1515 = 8'he2 == local_offset_1 ? phv_data_226 : _GEN_1514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1516 = 8'he3 == local_offset_1 ? phv_data_227 : _GEN_1515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1517 = 8'he4 == local_offset_1 ? phv_data_228 : _GEN_1516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1518 = 8'he5 == local_offset_1 ? phv_data_229 : _GEN_1517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1519 = 8'he6 == local_offset_1 ? phv_data_230 : _GEN_1518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1520 = 8'he7 == local_offset_1 ? phv_data_231 : _GEN_1519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1521 = 8'he8 == local_offset_1 ? phv_data_232 : _GEN_1520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1522 = 8'he9 == local_offset_1 ? phv_data_233 : _GEN_1521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1523 = 8'hea == local_offset_1 ? phv_data_234 : _GEN_1522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1524 = 8'heb == local_offset_1 ? phv_data_235 : _GEN_1523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1525 = 8'hec == local_offset_1 ? phv_data_236 : _GEN_1524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1526 = 8'hed == local_offset_1 ? phv_data_237 : _GEN_1525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1527 = 8'hee == local_offset_1 ? phv_data_238 : _GEN_1526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1528 = 8'hef == local_offset_1 ? phv_data_239 : _GEN_1527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1529 = 8'hf0 == local_offset_1 ? phv_data_240 : _GEN_1528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1530 = 8'hf1 == local_offset_1 ? phv_data_241 : _GEN_1529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1531 = 8'hf2 == local_offset_1 ? phv_data_242 : _GEN_1530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1532 = 8'hf3 == local_offset_1 ? phv_data_243 : _GEN_1531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1533 = 8'hf4 == local_offset_1 ? phv_data_244 : _GEN_1532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1534 = 8'hf5 == local_offset_1 ? phv_data_245 : _GEN_1533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1535 = 8'hf6 == local_offset_1 ? phv_data_246 : _GEN_1534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1536 = 8'hf7 == local_offset_1 ? phv_data_247 : _GEN_1535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1537 = 8'hf8 == local_offset_1 ? phv_data_248 : _GEN_1536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1538 = 8'hf9 == local_offset_1 ? phv_data_249 : _GEN_1537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1539 = 8'hfa == local_offset_1 ? phv_data_250 : _GEN_1538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1540 = 8'hfb == local_offset_1 ? phv_data_251 : _GEN_1539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1541 = 8'hfc == local_offset_1 ? phv_data_252 : _GEN_1540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1542 = 8'hfd == local_offset_1 ? phv_data_253 : _GEN_1541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1543 = 8'hfe == local_offset_1 ? phv_data_254 : _GEN_1542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1544 = 8'hff == local_offset_1 ? phv_data_255 : _GEN_1543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1546 = 8'h1 == _match_key_qbytes_1_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1547 = 8'h2 == _match_key_qbytes_1_T ? phv_data_2 : _GEN_1546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1548 = 8'h3 == _match_key_qbytes_1_T ? phv_data_3 : _GEN_1547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1549 = 8'h4 == _match_key_qbytes_1_T ? phv_data_4 : _GEN_1548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1550 = 8'h5 == _match_key_qbytes_1_T ? phv_data_5 : _GEN_1549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1551 = 8'h6 == _match_key_qbytes_1_T ? phv_data_6 : _GEN_1550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1552 = 8'h7 == _match_key_qbytes_1_T ? phv_data_7 : _GEN_1551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1553 = 8'h8 == _match_key_qbytes_1_T ? phv_data_8 : _GEN_1552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1554 = 8'h9 == _match_key_qbytes_1_T ? phv_data_9 : _GEN_1553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1555 = 8'ha == _match_key_qbytes_1_T ? phv_data_10 : _GEN_1554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1556 = 8'hb == _match_key_qbytes_1_T ? phv_data_11 : _GEN_1555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1557 = 8'hc == _match_key_qbytes_1_T ? phv_data_12 : _GEN_1556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1558 = 8'hd == _match_key_qbytes_1_T ? phv_data_13 : _GEN_1557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1559 = 8'he == _match_key_qbytes_1_T ? phv_data_14 : _GEN_1558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1560 = 8'hf == _match_key_qbytes_1_T ? phv_data_15 : _GEN_1559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1561 = 8'h10 == _match_key_qbytes_1_T ? phv_data_16 : _GEN_1560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1562 = 8'h11 == _match_key_qbytes_1_T ? phv_data_17 : _GEN_1561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1563 = 8'h12 == _match_key_qbytes_1_T ? phv_data_18 : _GEN_1562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1564 = 8'h13 == _match_key_qbytes_1_T ? phv_data_19 : _GEN_1563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1565 = 8'h14 == _match_key_qbytes_1_T ? phv_data_20 : _GEN_1564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1566 = 8'h15 == _match_key_qbytes_1_T ? phv_data_21 : _GEN_1565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1567 = 8'h16 == _match_key_qbytes_1_T ? phv_data_22 : _GEN_1566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1568 = 8'h17 == _match_key_qbytes_1_T ? phv_data_23 : _GEN_1567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1569 = 8'h18 == _match_key_qbytes_1_T ? phv_data_24 : _GEN_1568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1570 = 8'h19 == _match_key_qbytes_1_T ? phv_data_25 : _GEN_1569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1571 = 8'h1a == _match_key_qbytes_1_T ? phv_data_26 : _GEN_1570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1572 = 8'h1b == _match_key_qbytes_1_T ? phv_data_27 : _GEN_1571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1573 = 8'h1c == _match_key_qbytes_1_T ? phv_data_28 : _GEN_1572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1574 = 8'h1d == _match_key_qbytes_1_T ? phv_data_29 : _GEN_1573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1575 = 8'h1e == _match_key_qbytes_1_T ? phv_data_30 : _GEN_1574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1576 = 8'h1f == _match_key_qbytes_1_T ? phv_data_31 : _GEN_1575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1577 = 8'h20 == _match_key_qbytes_1_T ? phv_data_32 : _GEN_1576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1578 = 8'h21 == _match_key_qbytes_1_T ? phv_data_33 : _GEN_1577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1579 = 8'h22 == _match_key_qbytes_1_T ? phv_data_34 : _GEN_1578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1580 = 8'h23 == _match_key_qbytes_1_T ? phv_data_35 : _GEN_1579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1581 = 8'h24 == _match_key_qbytes_1_T ? phv_data_36 : _GEN_1580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1582 = 8'h25 == _match_key_qbytes_1_T ? phv_data_37 : _GEN_1581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1583 = 8'h26 == _match_key_qbytes_1_T ? phv_data_38 : _GEN_1582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1584 = 8'h27 == _match_key_qbytes_1_T ? phv_data_39 : _GEN_1583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1585 = 8'h28 == _match_key_qbytes_1_T ? phv_data_40 : _GEN_1584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1586 = 8'h29 == _match_key_qbytes_1_T ? phv_data_41 : _GEN_1585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1587 = 8'h2a == _match_key_qbytes_1_T ? phv_data_42 : _GEN_1586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1588 = 8'h2b == _match_key_qbytes_1_T ? phv_data_43 : _GEN_1587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1589 = 8'h2c == _match_key_qbytes_1_T ? phv_data_44 : _GEN_1588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1590 = 8'h2d == _match_key_qbytes_1_T ? phv_data_45 : _GEN_1589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1591 = 8'h2e == _match_key_qbytes_1_T ? phv_data_46 : _GEN_1590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1592 = 8'h2f == _match_key_qbytes_1_T ? phv_data_47 : _GEN_1591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1593 = 8'h30 == _match_key_qbytes_1_T ? phv_data_48 : _GEN_1592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1594 = 8'h31 == _match_key_qbytes_1_T ? phv_data_49 : _GEN_1593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1595 = 8'h32 == _match_key_qbytes_1_T ? phv_data_50 : _GEN_1594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1596 = 8'h33 == _match_key_qbytes_1_T ? phv_data_51 : _GEN_1595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1597 = 8'h34 == _match_key_qbytes_1_T ? phv_data_52 : _GEN_1596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1598 = 8'h35 == _match_key_qbytes_1_T ? phv_data_53 : _GEN_1597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1599 = 8'h36 == _match_key_qbytes_1_T ? phv_data_54 : _GEN_1598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1600 = 8'h37 == _match_key_qbytes_1_T ? phv_data_55 : _GEN_1599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1601 = 8'h38 == _match_key_qbytes_1_T ? phv_data_56 : _GEN_1600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1602 = 8'h39 == _match_key_qbytes_1_T ? phv_data_57 : _GEN_1601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1603 = 8'h3a == _match_key_qbytes_1_T ? phv_data_58 : _GEN_1602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1604 = 8'h3b == _match_key_qbytes_1_T ? phv_data_59 : _GEN_1603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1605 = 8'h3c == _match_key_qbytes_1_T ? phv_data_60 : _GEN_1604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1606 = 8'h3d == _match_key_qbytes_1_T ? phv_data_61 : _GEN_1605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1607 = 8'h3e == _match_key_qbytes_1_T ? phv_data_62 : _GEN_1606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1608 = 8'h3f == _match_key_qbytes_1_T ? phv_data_63 : _GEN_1607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1609 = 8'h40 == _match_key_qbytes_1_T ? phv_data_64 : _GEN_1608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1610 = 8'h41 == _match_key_qbytes_1_T ? phv_data_65 : _GEN_1609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1611 = 8'h42 == _match_key_qbytes_1_T ? phv_data_66 : _GEN_1610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1612 = 8'h43 == _match_key_qbytes_1_T ? phv_data_67 : _GEN_1611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1613 = 8'h44 == _match_key_qbytes_1_T ? phv_data_68 : _GEN_1612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1614 = 8'h45 == _match_key_qbytes_1_T ? phv_data_69 : _GEN_1613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1615 = 8'h46 == _match_key_qbytes_1_T ? phv_data_70 : _GEN_1614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1616 = 8'h47 == _match_key_qbytes_1_T ? phv_data_71 : _GEN_1615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1617 = 8'h48 == _match_key_qbytes_1_T ? phv_data_72 : _GEN_1616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1618 = 8'h49 == _match_key_qbytes_1_T ? phv_data_73 : _GEN_1617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1619 = 8'h4a == _match_key_qbytes_1_T ? phv_data_74 : _GEN_1618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1620 = 8'h4b == _match_key_qbytes_1_T ? phv_data_75 : _GEN_1619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1621 = 8'h4c == _match_key_qbytes_1_T ? phv_data_76 : _GEN_1620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1622 = 8'h4d == _match_key_qbytes_1_T ? phv_data_77 : _GEN_1621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1623 = 8'h4e == _match_key_qbytes_1_T ? phv_data_78 : _GEN_1622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1624 = 8'h4f == _match_key_qbytes_1_T ? phv_data_79 : _GEN_1623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1625 = 8'h50 == _match_key_qbytes_1_T ? phv_data_80 : _GEN_1624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1626 = 8'h51 == _match_key_qbytes_1_T ? phv_data_81 : _GEN_1625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1627 = 8'h52 == _match_key_qbytes_1_T ? phv_data_82 : _GEN_1626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1628 = 8'h53 == _match_key_qbytes_1_T ? phv_data_83 : _GEN_1627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1629 = 8'h54 == _match_key_qbytes_1_T ? phv_data_84 : _GEN_1628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1630 = 8'h55 == _match_key_qbytes_1_T ? phv_data_85 : _GEN_1629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1631 = 8'h56 == _match_key_qbytes_1_T ? phv_data_86 : _GEN_1630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1632 = 8'h57 == _match_key_qbytes_1_T ? phv_data_87 : _GEN_1631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1633 = 8'h58 == _match_key_qbytes_1_T ? phv_data_88 : _GEN_1632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1634 = 8'h59 == _match_key_qbytes_1_T ? phv_data_89 : _GEN_1633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1635 = 8'h5a == _match_key_qbytes_1_T ? phv_data_90 : _GEN_1634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1636 = 8'h5b == _match_key_qbytes_1_T ? phv_data_91 : _GEN_1635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1637 = 8'h5c == _match_key_qbytes_1_T ? phv_data_92 : _GEN_1636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1638 = 8'h5d == _match_key_qbytes_1_T ? phv_data_93 : _GEN_1637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1639 = 8'h5e == _match_key_qbytes_1_T ? phv_data_94 : _GEN_1638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1640 = 8'h5f == _match_key_qbytes_1_T ? phv_data_95 : _GEN_1639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1641 = 8'h60 == _match_key_qbytes_1_T ? phv_data_96 : _GEN_1640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1642 = 8'h61 == _match_key_qbytes_1_T ? phv_data_97 : _GEN_1641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1643 = 8'h62 == _match_key_qbytes_1_T ? phv_data_98 : _GEN_1642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1644 = 8'h63 == _match_key_qbytes_1_T ? phv_data_99 : _GEN_1643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1645 = 8'h64 == _match_key_qbytes_1_T ? phv_data_100 : _GEN_1644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1646 = 8'h65 == _match_key_qbytes_1_T ? phv_data_101 : _GEN_1645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1647 = 8'h66 == _match_key_qbytes_1_T ? phv_data_102 : _GEN_1646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1648 = 8'h67 == _match_key_qbytes_1_T ? phv_data_103 : _GEN_1647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1649 = 8'h68 == _match_key_qbytes_1_T ? phv_data_104 : _GEN_1648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1650 = 8'h69 == _match_key_qbytes_1_T ? phv_data_105 : _GEN_1649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1651 = 8'h6a == _match_key_qbytes_1_T ? phv_data_106 : _GEN_1650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1652 = 8'h6b == _match_key_qbytes_1_T ? phv_data_107 : _GEN_1651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1653 = 8'h6c == _match_key_qbytes_1_T ? phv_data_108 : _GEN_1652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1654 = 8'h6d == _match_key_qbytes_1_T ? phv_data_109 : _GEN_1653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1655 = 8'h6e == _match_key_qbytes_1_T ? phv_data_110 : _GEN_1654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1656 = 8'h6f == _match_key_qbytes_1_T ? phv_data_111 : _GEN_1655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1657 = 8'h70 == _match_key_qbytes_1_T ? phv_data_112 : _GEN_1656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1658 = 8'h71 == _match_key_qbytes_1_T ? phv_data_113 : _GEN_1657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1659 = 8'h72 == _match_key_qbytes_1_T ? phv_data_114 : _GEN_1658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1660 = 8'h73 == _match_key_qbytes_1_T ? phv_data_115 : _GEN_1659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1661 = 8'h74 == _match_key_qbytes_1_T ? phv_data_116 : _GEN_1660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1662 = 8'h75 == _match_key_qbytes_1_T ? phv_data_117 : _GEN_1661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1663 = 8'h76 == _match_key_qbytes_1_T ? phv_data_118 : _GEN_1662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1664 = 8'h77 == _match_key_qbytes_1_T ? phv_data_119 : _GEN_1663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1665 = 8'h78 == _match_key_qbytes_1_T ? phv_data_120 : _GEN_1664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1666 = 8'h79 == _match_key_qbytes_1_T ? phv_data_121 : _GEN_1665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1667 = 8'h7a == _match_key_qbytes_1_T ? phv_data_122 : _GEN_1666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1668 = 8'h7b == _match_key_qbytes_1_T ? phv_data_123 : _GEN_1667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1669 = 8'h7c == _match_key_qbytes_1_T ? phv_data_124 : _GEN_1668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1670 = 8'h7d == _match_key_qbytes_1_T ? phv_data_125 : _GEN_1669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1671 = 8'h7e == _match_key_qbytes_1_T ? phv_data_126 : _GEN_1670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1672 = 8'h7f == _match_key_qbytes_1_T ? phv_data_127 : _GEN_1671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1673 = 8'h80 == _match_key_qbytes_1_T ? phv_data_128 : _GEN_1672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1674 = 8'h81 == _match_key_qbytes_1_T ? phv_data_129 : _GEN_1673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1675 = 8'h82 == _match_key_qbytes_1_T ? phv_data_130 : _GEN_1674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1676 = 8'h83 == _match_key_qbytes_1_T ? phv_data_131 : _GEN_1675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1677 = 8'h84 == _match_key_qbytes_1_T ? phv_data_132 : _GEN_1676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1678 = 8'h85 == _match_key_qbytes_1_T ? phv_data_133 : _GEN_1677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1679 = 8'h86 == _match_key_qbytes_1_T ? phv_data_134 : _GEN_1678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1680 = 8'h87 == _match_key_qbytes_1_T ? phv_data_135 : _GEN_1679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1681 = 8'h88 == _match_key_qbytes_1_T ? phv_data_136 : _GEN_1680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1682 = 8'h89 == _match_key_qbytes_1_T ? phv_data_137 : _GEN_1681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1683 = 8'h8a == _match_key_qbytes_1_T ? phv_data_138 : _GEN_1682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1684 = 8'h8b == _match_key_qbytes_1_T ? phv_data_139 : _GEN_1683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1685 = 8'h8c == _match_key_qbytes_1_T ? phv_data_140 : _GEN_1684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1686 = 8'h8d == _match_key_qbytes_1_T ? phv_data_141 : _GEN_1685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1687 = 8'h8e == _match_key_qbytes_1_T ? phv_data_142 : _GEN_1686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1688 = 8'h8f == _match_key_qbytes_1_T ? phv_data_143 : _GEN_1687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1689 = 8'h90 == _match_key_qbytes_1_T ? phv_data_144 : _GEN_1688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1690 = 8'h91 == _match_key_qbytes_1_T ? phv_data_145 : _GEN_1689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1691 = 8'h92 == _match_key_qbytes_1_T ? phv_data_146 : _GEN_1690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1692 = 8'h93 == _match_key_qbytes_1_T ? phv_data_147 : _GEN_1691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1693 = 8'h94 == _match_key_qbytes_1_T ? phv_data_148 : _GEN_1692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1694 = 8'h95 == _match_key_qbytes_1_T ? phv_data_149 : _GEN_1693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1695 = 8'h96 == _match_key_qbytes_1_T ? phv_data_150 : _GEN_1694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1696 = 8'h97 == _match_key_qbytes_1_T ? phv_data_151 : _GEN_1695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1697 = 8'h98 == _match_key_qbytes_1_T ? phv_data_152 : _GEN_1696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1698 = 8'h99 == _match_key_qbytes_1_T ? phv_data_153 : _GEN_1697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1699 = 8'h9a == _match_key_qbytes_1_T ? phv_data_154 : _GEN_1698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1700 = 8'h9b == _match_key_qbytes_1_T ? phv_data_155 : _GEN_1699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1701 = 8'h9c == _match_key_qbytes_1_T ? phv_data_156 : _GEN_1700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1702 = 8'h9d == _match_key_qbytes_1_T ? phv_data_157 : _GEN_1701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1703 = 8'h9e == _match_key_qbytes_1_T ? phv_data_158 : _GEN_1702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1704 = 8'h9f == _match_key_qbytes_1_T ? phv_data_159 : _GEN_1703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1705 = 8'ha0 == _match_key_qbytes_1_T ? phv_data_160 : _GEN_1704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1706 = 8'ha1 == _match_key_qbytes_1_T ? phv_data_161 : _GEN_1705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1707 = 8'ha2 == _match_key_qbytes_1_T ? phv_data_162 : _GEN_1706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1708 = 8'ha3 == _match_key_qbytes_1_T ? phv_data_163 : _GEN_1707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1709 = 8'ha4 == _match_key_qbytes_1_T ? phv_data_164 : _GEN_1708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1710 = 8'ha5 == _match_key_qbytes_1_T ? phv_data_165 : _GEN_1709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1711 = 8'ha6 == _match_key_qbytes_1_T ? phv_data_166 : _GEN_1710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1712 = 8'ha7 == _match_key_qbytes_1_T ? phv_data_167 : _GEN_1711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1713 = 8'ha8 == _match_key_qbytes_1_T ? phv_data_168 : _GEN_1712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1714 = 8'ha9 == _match_key_qbytes_1_T ? phv_data_169 : _GEN_1713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1715 = 8'haa == _match_key_qbytes_1_T ? phv_data_170 : _GEN_1714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1716 = 8'hab == _match_key_qbytes_1_T ? phv_data_171 : _GEN_1715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1717 = 8'hac == _match_key_qbytes_1_T ? phv_data_172 : _GEN_1716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1718 = 8'had == _match_key_qbytes_1_T ? phv_data_173 : _GEN_1717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1719 = 8'hae == _match_key_qbytes_1_T ? phv_data_174 : _GEN_1718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1720 = 8'haf == _match_key_qbytes_1_T ? phv_data_175 : _GEN_1719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1721 = 8'hb0 == _match_key_qbytes_1_T ? phv_data_176 : _GEN_1720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1722 = 8'hb1 == _match_key_qbytes_1_T ? phv_data_177 : _GEN_1721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1723 = 8'hb2 == _match_key_qbytes_1_T ? phv_data_178 : _GEN_1722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1724 = 8'hb3 == _match_key_qbytes_1_T ? phv_data_179 : _GEN_1723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1725 = 8'hb4 == _match_key_qbytes_1_T ? phv_data_180 : _GEN_1724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1726 = 8'hb5 == _match_key_qbytes_1_T ? phv_data_181 : _GEN_1725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1727 = 8'hb6 == _match_key_qbytes_1_T ? phv_data_182 : _GEN_1726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1728 = 8'hb7 == _match_key_qbytes_1_T ? phv_data_183 : _GEN_1727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1729 = 8'hb8 == _match_key_qbytes_1_T ? phv_data_184 : _GEN_1728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1730 = 8'hb9 == _match_key_qbytes_1_T ? phv_data_185 : _GEN_1729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1731 = 8'hba == _match_key_qbytes_1_T ? phv_data_186 : _GEN_1730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1732 = 8'hbb == _match_key_qbytes_1_T ? phv_data_187 : _GEN_1731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1733 = 8'hbc == _match_key_qbytes_1_T ? phv_data_188 : _GEN_1732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1734 = 8'hbd == _match_key_qbytes_1_T ? phv_data_189 : _GEN_1733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1735 = 8'hbe == _match_key_qbytes_1_T ? phv_data_190 : _GEN_1734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1736 = 8'hbf == _match_key_qbytes_1_T ? phv_data_191 : _GEN_1735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1737 = 8'hc0 == _match_key_qbytes_1_T ? phv_data_192 : _GEN_1736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1738 = 8'hc1 == _match_key_qbytes_1_T ? phv_data_193 : _GEN_1737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1739 = 8'hc2 == _match_key_qbytes_1_T ? phv_data_194 : _GEN_1738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1740 = 8'hc3 == _match_key_qbytes_1_T ? phv_data_195 : _GEN_1739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1741 = 8'hc4 == _match_key_qbytes_1_T ? phv_data_196 : _GEN_1740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1742 = 8'hc5 == _match_key_qbytes_1_T ? phv_data_197 : _GEN_1741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1743 = 8'hc6 == _match_key_qbytes_1_T ? phv_data_198 : _GEN_1742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1744 = 8'hc7 == _match_key_qbytes_1_T ? phv_data_199 : _GEN_1743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1745 = 8'hc8 == _match_key_qbytes_1_T ? phv_data_200 : _GEN_1744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1746 = 8'hc9 == _match_key_qbytes_1_T ? phv_data_201 : _GEN_1745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1747 = 8'hca == _match_key_qbytes_1_T ? phv_data_202 : _GEN_1746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1748 = 8'hcb == _match_key_qbytes_1_T ? phv_data_203 : _GEN_1747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1749 = 8'hcc == _match_key_qbytes_1_T ? phv_data_204 : _GEN_1748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1750 = 8'hcd == _match_key_qbytes_1_T ? phv_data_205 : _GEN_1749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1751 = 8'hce == _match_key_qbytes_1_T ? phv_data_206 : _GEN_1750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1752 = 8'hcf == _match_key_qbytes_1_T ? phv_data_207 : _GEN_1751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1753 = 8'hd0 == _match_key_qbytes_1_T ? phv_data_208 : _GEN_1752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1754 = 8'hd1 == _match_key_qbytes_1_T ? phv_data_209 : _GEN_1753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1755 = 8'hd2 == _match_key_qbytes_1_T ? phv_data_210 : _GEN_1754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1756 = 8'hd3 == _match_key_qbytes_1_T ? phv_data_211 : _GEN_1755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1757 = 8'hd4 == _match_key_qbytes_1_T ? phv_data_212 : _GEN_1756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1758 = 8'hd5 == _match_key_qbytes_1_T ? phv_data_213 : _GEN_1757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1759 = 8'hd6 == _match_key_qbytes_1_T ? phv_data_214 : _GEN_1758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1760 = 8'hd7 == _match_key_qbytes_1_T ? phv_data_215 : _GEN_1759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1761 = 8'hd8 == _match_key_qbytes_1_T ? phv_data_216 : _GEN_1760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1762 = 8'hd9 == _match_key_qbytes_1_T ? phv_data_217 : _GEN_1761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1763 = 8'hda == _match_key_qbytes_1_T ? phv_data_218 : _GEN_1762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1764 = 8'hdb == _match_key_qbytes_1_T ? phv_data_219 : _GEN_1763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1765 = 8'hdc == _match_key_qbytes_1_T ? phv_data_220 : _GEN_1764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1766 = 8'hdd == _match_key_qbytes_1_T ? phv_data_221 : _GEN_1765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1767 = 8'hde == _match_key_qbytes_1_T ? phv_data_222 : _GEN_1766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1768 = 8'hdf == _match_key_qbytes_1_T ? phv_data_223 : _GEN_1767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1769 = 8'he0 == _match_key_qbytes_1_T ? phv_data_224 : _GEN_1768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1770 = 8'he1 == _match_key_qbytes_1_T ? phv_data_225 : _GEN_1769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1771 = 8'he2 == _match_key_qbytes_1_T ? phv_data_226 : _GEN_1770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1772 = 8'he3 == _match_key_qbytes_1_T ? phv_data_227 : _GEN_1771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1773 = 8'he4 == _match_key_qbytes_1_T ? phv_data_228 : _GEN_1772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1774 = 8'he5 == _match_key_qbytes_1_T ? phv_data_229 : _GEN_1773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1775 = 8'he6 == _match_key_qbytes_1_T ? phv_data_230 : _GEN_1774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1776 = 8'he7 == _match_key_qbytes_1_T ? phv_data_231 : _GEN_1775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1777 = 8'he8 == _match_key_qbytes_1_T ? phv_data_232 : _GEN_1776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1778 = 8'he9 == _match_key_qbytes_1_T ? phv_data_233 : _GEN_1777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1779 = 8'hea == _match_key_qbytes_1_T ? phv_data_234 : _GEN_1778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1780 = 8'heb == _match_key_qbytes_1_T ? phv_data_235 : _GEN_1779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1781 = 8'hec == _match_key_qbytes_1_T ? phv_data_236 : _GEN_1780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1782 = 8'hed == _match_key_qbytes_1_T ? phv_data_237 : _GEN_1781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1783 = 8'hee == _match_key_qbytes_1_T ? phv_data_238 : _GEN_1782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1784 = 8'hef == _match_key_qbytes_1_T ? phv_data_239 : _GEN_1783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1785 = 8'hf0 == _match_key_qbytes_1_T ? phv_data_240 : _GEN_1784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1786 = 8'hf1 == _match_key_qbytes_1_T ? phv_data_241 : _GEN_1785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1787 = 8'hf2 == _match_key_qbytes_1_T ? phv_data_242 : _GEN_1786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1788 = 8'hf3 == _match_key_qbytes_1_T ? phv_data_243 : _GEN_1787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1789 = 8'hf4 == _match_key_qbytes_1_T ? phv_data_244 : _GEN_1788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1790 = 8'hf5 == _match_key_qbytes_1_T ? phv_data_245 : _GEN_1789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1791 = 8'hf6 == _match_key_qbytes_1_T ? phv_data_246 : _GEN_1790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1792 = 8'hf7 == _match_key_qbytes_1_T ? phv_data_247 : _GEN_1791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1793 = 8'hf8 == _match_key_qbytes_1_T ? phv_data_248 : _GEN_1792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1794 = 8'hf9 == _match_key_qbytes_1_T ? phv_data_249 : _GEN_1793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1795 = 8'hfa == _match_key_qbytes_1_T ? phv_data_250 : _GEN_1794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1796 = 8'hfb == _match_key_qbytes_1_T ? phv_data_251 : _GEN_1795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1797 = 8'hfc == _match_key_qbytes_1_T ? phv_data_252 : _GEN_1796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1798 = 8'hfd == _match_key_qbytes_1_T ? phv_data_253 : _GEN_1797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1799 = 8'hfe == _match_key_qbytes_1_T ? phv_data_254 : _GEN_1798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1800 = 8'hff == _match_key_qbytes_1_T ? phv_data_255 : _GEN_1799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1802 = 8'h1 == _match_key_qbytes_1_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1803 = 8'h2 == _match_key_qbytes_1_T_1 ? phv_data_2 : _GEN_1802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1804 = 8'h3 == _match_key_qbytes_1_T_1 ? phv_data_3 : _GEN_1803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1805 = 8'h4 == _match_key_qbytes_1_T_1 ? phv_data_4 : _GEN_1804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1806 = 8'h5 == _match_key_qbytes_1_T_1 ? phv_data_5 : _GEN_1805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1807 = 8'h6 == _match_key_qbytes_1_T_1 ? phv_data_6 : _GEN_1806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1808 = 8'h7 == _match_key_qbytes_1_T_1 ? phv_data_7 : _GEN_1807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1809 = 8'h8 == _match_key_qbytes_1_T_1 ? phv_data_8 : _GEN_1808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1810 = 8'h9 == _match_key_qbytes_1_T_1 ? phv_data_9 : _GEN_1809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1811 = 8'ha == _match_key_qbytes_1_T_1 ? phv_data_10 : _GEN_1810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1812 = 8'hb == _match_key_qbytes_1_T_1 ? phv_data_11 : _GEN_1811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1813 = 8'hc == _match_key_qbytes_1_T_1 ? phv_data_12 : _GEN_1812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1814 = 8'hd == _match_key_qbytes_1_T_1 ? phv_data_13 : _GEN_1813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1815 = 8'he == _match_key_qbytes_1_T_1 ? phv_data_14 : _GEN_1814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1816 = 8'hf == _match_key_qbytes_1_T_1 ? phv_data_15 : _GEN_1815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1817 = 8'h10 == _match_key_qbytes_1_T_1 ? phv_data_16 : _GEN_1816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1818 = 8'h11 == _match_key_qbytes_1_T_1 ? phv_data_17 : _GEN_1817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1819 = 8'h12 == _match_key_qbytes_1_T_1 ? phv_data_18 : _GEN_1818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1820 = 8'h13 == _match_key_qbytes_1_T_1 ? phv_data_19 : _GEN_1819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1821 = 8'h14 == _match_key_qbytes_1_T_1 ? phv_data_20 : _GEN_1820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1822 = 8'h15 == _match_key_qbytes_1_T_1 ? phv_data_21 : _GEN_1821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1823 = 8'h16 == _match_key_qbytes_1_T_1 ? phv_data_22 : _GEN_1822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1824 = 8'h17 == _match_key_qbytes_1_T_1 ? phv_data_23 : _GEN_1823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1825 = 8'h18 == _match_key_qbytes_1_T_1 ? phv_data_24 : _GEN_1824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1826 = 8'h19 == _match_key_qbytes_1_T_1 ? phv_data_25 : _GEN_1825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1827 = 8'h1a == _match_key_qbytes_1_T_1 ? phv_data_26 : _GEN_1826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1828 = 8'h1b == _match_key_qbytes_1_T_1 ? phv_data_27 : _GEN_1827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1829 = 8'h1c == _match_key_qbytes_1_T_1 ? phv_data_28 : _GEN_1828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1830 = 8'h1d == _match_key_qbytes_1_T_1 ? phv_data_29 : _GEN_1829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1831 = 8'h1e == _match_key_qbytes_1_T_1 ? phv_data_30 : _GEN_1830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1832 = 8'h1f == _match_key_qbytes_1_T_1 ? phv_data_31 : _GEN_1831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1833 = 8'h20 == _match_key_qbytes_1_T_1 ? phv_data_32 : _GEN_1832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1834 = 8'h21 == _match_key_qbytes_1_T_1 ? phv_data_33 : _GEN_1833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1835 = 8'h22 == _match_key_qbytes_1_T_1 ? phv_data_34 : _GEN_1834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1836 = 8'h23 == _match_key_qbytes_1_T_1 ? phv_data_35 : _GEN_1835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1837 = 8'h24 == _match_key_qbytes_1_T_1 ? phv_data_36 : _GEN_1836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1838 = 8'h25 == _match_key_qbytes_1_T_1 ? phv_data_37 : _GEN_1837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1839 = 8'h26 == _match_key_qbytes_1_T_1 ? phv_data_38 : _GEN_1838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1840 = 8'h27 == _match_key_qbytes_1_T_1 ? phv_data_39 : _GEN_1839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1841 = 8'h28 == _match_key_qbytes_1_T_1 ? phv_data_40 : _GEN_1840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1842 = 8'h29 == _match_key_qbytes_1_T_1 ? phv_data_41 : _GEN_1841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1843 = 8'h2a == _match_key_qbytes_1_T_1 ? phv_data_42 : _GEN_1842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1844 = 8'h2b == _match_key_qbytes_1_T_1 ? phv_data_43 : _GEN_1843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1845 = 8'h2c == _match_key_qbytes_1_T_1 ? phv_data_44 : _GEN_1844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1846 = 8'h2d == _match_key_qbytes_1_T_1 ? phv_data_45 : _GEN_1845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1847 = 8'h2e == _match_key_qbytes_1_T_1 ? phv_data_46 : _GEN_1846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1848 = 8'h2f == _match_key_qbytes_1_T_1 ? phv_data_47 : _GEN_1847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1849 = 8'h30 == _match_key_qbytes_1_T_1 ? phv_data_48 : _GEN_1848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1850 = 8'h31 == _match_key_qbytes_1_T_1 ? phv_data_49 : _GEN_1849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1851 = 8'h32 == _match_key_qbytes_1_T_1 ? phv_data_50 : _GEN_1850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1852 = 8'h33 == _match_key_qbytes_1_T_1 ? phv_data_51 : _GEN_1851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1853 = 8'h34 == _match_key_qbytes_1_T_1 ? phv_data_52 : _GEN_1852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1854 = 8'h35 == _match_key_qbytes_1_T_1 ? phv_data_53 : _GEN_1853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1855 = 8'h36 == _match_key_qbytes_1_T_1 ? phv_data_54 : _GEN_1854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1856 = 8'h37 == _match_key_qbytes_1_T_1 ? phv_data_55 : _GEN_1855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1857 = 8'h38 == _match_key_qbytes_1_T_1 ? phv_data_56 : _GEN_1856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1858 = 8'h39 == _match_key_qbytes_1_T_1 ? phv_data_57 : _GEN_1857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1859 = 8'h3a == _match_key_qbytes_1_T_1 ? phv_data_58 : _GEN_1858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1860 = 8'h3b == _match_key_qbytes_1_T_1 ? phv_data_59 : _GEN_1859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1861 = 8'h3c == _match_key_qbytes_1_T_1 ? phv_data_60 : _GEN_1860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1862 = 8'h3d == _match_key_qbytes_1_T_1 ? phv_data_61 : _GEN_1861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1863 = 8'h3e == _match_key_qbytes_1_T_1 ? phv_data_62 : _GEN_1862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1864 = 8'h3f == _match_key_qbytes_1_T_1 ? phv_data_63 : _GEN_1863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1865 = 8'h40 == _match_key_qbytes_1_T_1 ? phv_data_64 : _GEN_1864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1866 = 8'h41 == _match_key_qbytes_1_T_1 ? phv_data_65 : _GEN_1865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1867 = 8'h42 == _match_key_qbytes_1_T_1 ? phv_data_66 : _GEN_1866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1868 = 8'h43 == _match_key_qbytes_1_T_1 ? phv_data_67 : _GEN_1867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1869 = 8'h44 == _match_key_qbytes_1_T_1 ? phv_data_68 : _GEN_1868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1870 = 8'h45 == _match_key_qbytes_1_T_1 ? phv_data_69 : _GEN_1869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1871 = 8'h46 == _match_key_qbytes_1_T_1 ? phv_data_70 : _GEN_1870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1872 = 8'h47 == _match_key_qbytes_1_T_1 ? phv_data_71 : _GEN_1871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1873 = 8'h48 == _match_key_qbytes_1_T_1 ? phv_data_72 : _GEN_1872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1874 = 8'h49 == _match_key_qbytes_1_T_1 ? phv_data_73 : _GEN_1873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1875 = 8'h4a == _match_key_qbytes_1_T_1 ? phv_data_74 : _GEN_1874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1876 = 8'h4b == _match_key_qbytes_1_T_1 ? phv_data_75 : _GEN_1875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1877 = 8'h4c == _match_key_qbytes_1_T_1 ? phv_data_76 : _GEN_1876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1878 = 8'h4d == _match_key_qbytes_1_T_1 ? phv_data_77 : _GEN_1877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1879 = 8'h4e == _match_key_qbytes_1_T_1 ? phv_data_78 : _GEN_1878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1880 = 8'h4f == _match_key_qbytes_1_T_1 ? phv_data_79 : _GEN_1879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1881 = 8'h50 == _match_key_qbytes_1_T_1 ? phv_data_80 : _GEN_1880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1882 = 8'h51 == _match_key_qbytes_1_T_1 ? phv_data_81 : _GEN_1881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1883 = 8'h52 == _match_key_qbytes_1_T_1 ? phv_data_82 : _GEN_1882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1884 = 8'h53 == _match_key_qbytes_1_T_1 ? phv_data_83 : _GEN_1883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1885 = 8'h54 == _match_key_qbytes_1_T_1 ? phv_data_84 : _GEN_1884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1886 = 8'h55 == _match_key_qbytes_1_T_1 ? phv_data_85 : _GEN_1885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1887 = 8'h56 == _match_key_qbytes_1_T_1 ? phv_data_86 : _GEN_1886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1888 = 8'h57 == _match_key_qbytes_1_T_1 ? phv_data_87 : _GEN_1887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1889 = 8'h58 == _match_key_qbytes_1_T_1 ? phv_data_88 : _GEN_1888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1890 = 8'h59 == _match_key_qbytes_1_T_1 ? phv_data_89 : _GEN_1889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1891 = 8'h5a == _match_key_qbytes_1_T_1 ? phv_data_90 : _GEN_1890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1892 = 8'h5b == _match_key_qbytes_1_T_1 ? phv_data_91 : _GEN_1891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1893 = 8'h5c == _match_key_qbytes_1_T_1 ? phv_data_92 : _GEN_1892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1894 = 8'h5d == _match_key_qbytes_1_T_1 ? phv_data_93 : _GEN_1893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1895 = 8'h5e == _match_key_qbytes_1_T_1 ? phv_data_94 : _GEN_1894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1896 = 8'h5f == _match_key_qbytes_1_T_1 ? phv_data_95 : _GEN_1895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1897 = 8'h60 == _match_key_qbytes_1_T_1 ? phv_data_96 : _GEN_1896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1898 = 8'h61 == _match_key_qbytes_1_T_1 ? phv_data_97 : _GEN_1897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1899 = 8'h62 == _match_key_qbytes_1_T_1 ? phv_data_98 : _GEN_1898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1900 = 8'h63 == _match_key_qbytes_1_T_1 ? phv_data_99 : _GEN_1899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1901 = 8'h64 == _match_key_qbytes_1_T_1 ? phv_data_100 : _GEN_1900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1902 = 8'h65 == _match_key_qbytes_1_T_1 ? phv_data_101 : _GEN_1901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1903 = 8'h66 == _match_key_qbytes_1_T_1 ? phv_data_102 : _GEN_1902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1904 = 8'h67 == _match_key_qbytes_1_T_1 ? phv_data_103 : _GEN_1903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1905 = 8'h68 == _match_key_qbytes_1_T_1 ? phv_data_104 : _GEN_1904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1906 = 8'h69 == _match_key_qbytes_1_T_1 ? phv_data_105 : _GEN_1905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1907 = 8'h6a == _match_key_qbytes_1_T_1 ? phv_data_106 : _GEN_1906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1908 = 8'h6b == _match_key_qbytes_1_T_1 ? phv_data_107 : _GEN_1907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1909 = 8'h6c == _match_key_qbytes_1_T_1 ? phv_data_108 : _GEN_1908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1910 = 8'h6d == _match_key_qbytes_1_T_1 ? phv_data_109 : _GEN_1909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1911 = 8'h6e == _match_key_qbytes_1_T_1 ? phv_data_110 : _GEN_1910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1912 = 8'h6f == _match_key_qbytes_1_T_1 ? phv_data_111 : _GEN_1911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1913 = 8'h70 == _match_key_qbytes_1_T_1 ? phv_data_112 : _GEN_1912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1914 = 8'h71 == _match_key_qbytes_1_T_1 ? phv_data_113 : _GEN_1913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1915 = 8'h72 == _match_key_qbytes_1_T_1 ? phv_data_114 : _GEN_1914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1916 = 8'h73 == _match_key_qbytes_1_T_1 ? phv_data_115 : _GEN_1915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1917 = 8'h74 == _match_key_qbytes_1_T_1 ? phv_data_116 : _GEN_1916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1918 = 8'h75 == _match_key_qbytes_1_T_1 ? phv_data_117 : _GEN_1917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1919 = 8'h76 == _match_key_qbytes_1_T_1 ? phv_data_118 : _GEN_1918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1920 = 8'h77 == _match_key_qbytes_1_T_1 ? phv_data_119 : _GEN_1919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1921 = 8'h78 == _match_key_qbytes_1_T_1 ? phv_data_120 : _GEN_1920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1922 = 8'h79 == _match_key_qbytes_1_T_1 ? phv_data_121 : _GEN_1921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1923 = 8'h7a == _match_key_qbytes_1_T_1 ? phv_data_122 : _GEN_1922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1924 = 8'h7b == _match_key_qbytes_1_T_1 ? phv_data_123 : _GEN_1923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1925 = 8'h7c == _match_key_qbytes_1_T_1 ? phv_data_124 : _GEN_1924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1926 = 8'h7d == _match_key_qbytes_1_T_1 ? phv_data_125 : _GEN_1925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1927 = 8'h7e == _match_key_qbytes_1_T_1 ? phv_data_126 : _GEN_1926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1928 = 8'h7f == _match_key_qbytes_1_T_1 ? phv_data_127 : _GEN_1927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1929 = 8'h80 == _match_key_qbytes_1_T_1 ? phv_data_128 : _GEN_1928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1930 = 8'h81 == _match_key_qbytes_1_T_1 ? phv_data_129 : _GEN_1929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1931 = 8'h82 == _match_key_qbytes_1_T_1 ? phv_data_130 : _GEN_1930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1932 = 8'h83 == _match_key_qbytes_1_T_1 ? phv_data_131 : _GEN_1931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1933 = 8'h84 == _match_key_qbytes_1_T_1 ? phv_data_132 : _GEN_1932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1934 = 8'h85 == _match_key_qbytes_1_T_1 ? phv_data_133 : _GEN_1933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1935 = 8'h86 == _match_key_qbytes_1_T_1 ? phv_data_134 : _GEN_1934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1936 = 8'h87 == _match_key_qbytes_1_T_1 ? phv_data_135 : _GEN_1935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1937 = 8'h88 == _match_key_qbytes_1_T_1 ? phv_data_136 : _GEN_1936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1938 = 8'h89 == _match_key_qbytes_1_T_1 ? phv_data_137 : _GEN_1937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1939 = 8'h8a == _match_key_qbytes_1_T_1 ? phv_data_138 : _GEN_1938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1940 = 8'h8b == _match_key_qbytes_1_T_1 ? phv_data_139 : _GEN_1939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1941 = 8'h8c == _match_key_qbytes_1_T_1 ? phv_data_140 : _GEN_1940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1942 = 8'h8d == _match_key_qbytes_1_T_1 ? phv_data_141 : _GEN_1941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1943 = 8'h8e == _match_key_qbytes_1_T_1 ? phv_data_142 : _GEN_1942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1944 = 8'h8f == _match_key_qbytes_1_T_1 ? phv_data_143 : _GEN_1943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1945 = 8'h90 == _match_key_qbytes_1_T_1 ? phv_data_144 : _GEN_1944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1946 = 8'h91 == _match_key_qbytes_1_T_1 ? phv_data_145 : _GEN_1945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1947 = 8'h92 == _match_key_qbytes_1_T_1 ? phv_data_146 : _GEN_1946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1948 = 8'h93 == _match_key_qbytes_1_T_1 ? phv_data_147 : _GEN_1947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1949 = 8'h94 == _match_key_qbytes_1_T_1 ? phv_data_148 : _GEN_1948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1950 = 8'h95 == _match_key_qbytes_1_T_1 ? phv_data_149 : _GEN_1949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1951 = 8'h96 == _match_key_qbytes_1_T_1 ? phv_data_150 : _GEN_1950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1952 = 8'h97 == _match_key_qbytes_1_T_1 ? phv_data_151 : _GEN_1951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1953 = 8'h98 == _match_key_qbytes_1_T_1 ? phv_data_152 : _GEN_1952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1954 = 8'h99 == _match_key_qbytes_1_T_1 ? phv_data_153 : _GEN_1953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1955 = 8'h9a == _match_key_qbytes_1_T_1 ? phv_data_154 : _GEN_1954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1956 = 8'h9b == _match_key_qbytes_1_T_1 ? phv_data_155 : _GEN_1955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1957 = 8'h9c == _match_key_qbytes_1_T_1 ? phv_data_156 : _GEN_1956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1958 = 8'h9d == _match_key_qbytes_1_T_1 ? phv_data_157 : _GEN_1957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1959 = 8'h9e == _match_key_qbytes_1_T_1 ? phv_data_158 : _GEN_1958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1960 = 8'h9f == _match_key_qbytes_1_T_1 ? phv_data_159 : _GEN_1959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1961 = 8'ha0 == _match_key_qbytes_1_T_1 ? phv_data_160 : _GEN_1960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1962 = 8'ha1 == _match_key_qbytes_1_T_1 ? phv_data_161 : _GEN_1961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1963 = 8'ha2 == _match_key_qbytes_1_T_1 ? phv_data_162 : _GEN_1962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1964 = 8'ha3 == _match_key_qbytes_1_T_1 ? phv_data_163 : _GEN_1963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1965 = 8'ha4 == _match_key_qbytes_1_T_1 ? phv_data_164 : _GEN_1964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1966 = 8'ha5 == _match_key_qbytes_1_T_1 ? phv_data_165 : _GEN_1965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1967 = 8'ha6 == _match_key_qbytes_1_T_1 ? phv_data_166 : _GEN_1966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1968 = 8'ha7 == _match_key_qbytes_1_T_1 ? phv_data_167 : _GEN_1967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1969 = 8'ha8 == _match_key_qbytes_1_T_1 ? phv_data_168 : _GEN_1968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1970 = 8'ha9 == _match_key_qbytes_1_T_1 ? phv_data_169 : _GEN_1969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1971 = 8'haa == _match_key_qbytes_1_T_1 ? phv_data_170 : _GEN_1970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1972 = 8'hab == _match_key_qbytes_1_T_1 ? phv_data_171 : _GEN_1971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1973 = 8'hac == _match_key_qbytes_1_T_1 ? phv_data_172 : _GEN_1972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1974 = 8'had == _match_key_qbytes_1_T_1 ? phv_data_173 : _GEN_1973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1975 = 8'hae == _match_key_qbytes_1_T_1 ? phv_data_174 : _GEN_1974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1976 = 8'haf == _match_key_qbytes_1_T_1 ? phv_data_175 : _GEN_1975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1977 = 8'hb0 == _match_key_qbytes_1_T_1 ? phv_data_176 : _GEN_1976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1978 = 8'hb1 == _match_key_qbytes_1_T_1 ? phv_data_177 : _GEN_1977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1979 = 8'hb2 == _match_key_qbytes_1_T_1 ? phv_data_178 : _GEN_1978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1980 = 8'hb3 == _match_key_qbytes_1_T_1 ? phv_data_179 : _GEN_1979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1981 = 8'hb4 == _match_key_qbytes_1_T_1 ? phv_data_180 : _GEN_1980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1982 = 8'hb5 == _match_key_qbytes_1_T_1 ? phv_data_181 : _GEN_1981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1983 = 8'hb6 == _match_key_qbytes_1_T_1 ? phv_data_182 : _GEN_1982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1984 = 8'hb7 == _match_key_qbytes_1_T_1 ? phv_data_183 : _GEN_1983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1985 = 8'hb8 == _match_key_qbytes_1_T_1 ? phv_data_184 : _GEN_1984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1986 = 8'hb9 == _match_key_qbytes_1_T_1 ? phv_data_185 : _GEN_1985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1987 = 8'hba == _match_key_qbytes_1_T_1 ? phv_data_186 : _GEN_1986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1988 = 8'hbb == _match_key_qbytes_1_T_1 ? phv_data_187 : _GEN_1987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1989 = 8'hbc == _match_key_qbytes_1_T_1 ? phv_data_188 : _GEN_1988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1990 = 8'hbd == _match_key_qbytes_1_T_1 ? phv_data_189 : _GEN_1989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1991 = 8'hbe == _match_key_qbytes_1_T_1 ? phv_data_190 : _GEN_1990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1992 = 8'hbf == _match_key_qbytes_1_T_1 ? phv_data_191 : _GEN_1991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1993 = 8'hc0 == _match_key_qbytes_1_T_1 ? phv_data_192 : _GEN_1992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1994 = 8'hc1 == _match_key_qbytes_1_T_1 ? phv_data_193 : _GEN_1993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1995 = 8'hc2 == _match_key_qbytes_1_T_1 ? phv_data_194 : _GEN_1994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1996 = 8'hc3 == _match_key_qbytes_1_T_1 ? phv_data_195 : _GEN_1995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1997 = 8'hc4 == _match_key_qbytes_1_T_1 ? phv_data_196 : _GEN_1996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1998 = 8'hc5 == _match_key_qbytes_1_T_1 ? phv_data_197 : _GEN_1997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1999 = 8'hc6 == _match_key_qbytes_1_T_1 ? phv_data_198 : _GEN_1998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2000 = 8'hc7 == _match_key_qbytes_1_T_1 ? phv_data_199 : _GEN_1999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2001 = 8'hc8 == _match_key_qbytes_1_T_1 ? phv_data_200 : _GEN_2000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2002 = 8'hc9 == _match_key_qbytes_1_T_1 ? phv_data_201 : _GEN_2001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2003 = 8'hca == _match_key_qbytes_1_T_1 ? phv_data_202 : _GEN_2002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2004 = 8'hcb == _match_key_qbytes_1_T_1 ? phv_data_203 : _GEN_2003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2005 = 8'hcc == _match_key_qbytes_1_T_1 ? phv_data_204 : _GEN_2004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2006 = 8'hcd == _match_key_qbytes_1_T_1 ? phv_data_205 : _GEN_2005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2007 = 8'hce == _match_key_qbytes_1_T_1 ? phv_data_206 : _GEN_2006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2008 = 8'hcf == _match_key_qbytes_1_T_1 ? phv_data_207 : _GEN_2007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2009 = 8'hd0 == _match_key_qbytes_1_T_1 ? phv_data_208 : _GEN_2008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2010 = 8'hd1 == _match_key_qbytes_1_T_1 ? phv_data_209 : _GEN_2009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2011 = 8'hd2 == _match_key_qbytes_1_T_1 ? phv_data_210 : _GEN_2010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2012 = 8'hd3 == _match_key_qbytes_1_T_1 ? phv_data_211 : _GEN_2011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2013 = 8'hd4 == _match_key_qbytes_1_T_1 ? phv_data_212 : _GEN_2012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2014 = 8'hd5 == _match_key_qbytes_1_T_1 ? phv_data_213 : _GEN_2013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2015 = 8'hd6 == _match_key_qbytes_1_T_1 ? phv_data_214 : _GEN_2014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2016 = 8'hd7 == _match_key_qbytes_1_T_1 ? phv_data_215 : _GEN_2015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2017 = 8'hd8 == _match_key_qbytes_1_T_1 ? phv_data_216 : _GEN_2016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2018 = 8'hd9 == _match_key_qbytes_1_T_1 ? phv_data_217 : _GEN_2017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2019 = 8'hda == _match_key_qbytes_1_T_1 ? phv_data_218 : _GEN_2018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2020 = 8'hdb == _match_key_qbytes_1_T_1 ? phv_data_219 : _GEN_2019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2021 = 8'hdc == _match_key_qbytes_1_T_1 ? phv_data_220 : _GEN_2020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2022 = 8'hdd == _match_key_qbytes_1_T_1 ? phv_data_221 : _GEN_2021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2023 = 8'hde == _match_key_qbytes_1_T_1 ? phv_data_222 : _GEN_2022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2024 = 8'hdf == _match_key_qbytes_1_T_1 ? phv_data_223 : _GEN_2023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2025 = 8'he0 == _match_key_qbytes_1_T_1 ? phv_data_224 : _GEN_2024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2026 = 8'he1 == _match_key_qbytes_1_T_1 ? phv_data_225 : _GEN_2025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2027 = 8'he2 == _match_key_qbytes_1_T_1 ? phv_data_226 : _GEN_2026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2028 = 8'he3 == _match_key_qbytes_1_T_1 ? phv_data_227 : _GEN_2027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2029 = 8'he4 == _match_key_qbytes_1_T_1 ? phv_data_228 : _GEN_2028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2030 = 8'he5 == _match_key_qbytes_1_T_1 ? phv_data_229 : _GEN_2029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2031 = 8'he6 == _match_key_qbytes_1_T_1 ? phv_data_230 : _GEN_2030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2032 = 8'he7 == _match_key_qbytes_1_T_1 ? phv_data_231 : _GEN_2031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2033 = 8'he8 == _match_key_qbytes_1_T_1 ? phv_data_232 : _GEN_2032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2034 = 8'he9 == _match_key_qbytes_1_T_1 ? phv_data_233 : _GEN_2033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2035 = 8'hea == _match_key_qbytes_1_T_1 ? phv_data_234 : _GEN_2034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2036 = 8'heb == _match_key_qbytes_1_T_1 ? phv_data_235 : _GEN_2035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2037 = 8'hec == _match_key_qbytes_1_T_1 ? phv_data_236 : _GEN_2036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2038 = 8'hed == _match_key_qbytes_1_T_1 ? phv_data_237 : _GEN_2037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2039 = 8'hee == _match_key_qbytes_1_T_1 ? phv_data_238 : _GEN_2038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2040 = 8'hef == _match_key_qbytes_1_T_1 ? phv_data_239 : _GEN_2039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2041 = 8'hf0 == _match_key_qbytes_1_T_1 ? phv_data_240 : _GEN_2040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2042 = 8'hf1 == _match_key_qbytes_1_T_1 ? phv_data_241 : _GEN_2041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2043 = 8'hf2 == _match_key_qbytes_1_T_1 ? phv_data_242 : _GEN_2042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2044 = 8'hf3 == _match_key_qbytes_1_T_1 ? phv_data_243 : _GEN_2043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2045 = 8'hf4 == _match_key_qbytes_1_T_1 ? phv_data_244 : _GEN_2044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2046 = 8'hf5 == _match_key_qbytes_1_T_1 ? phv_data_245 : _GEN_2045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2047 = 8'hf6 == _match_key_qbytes_1_T_1 ? phv_data_246 : _GEN_2046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2048 = 8'hf7 == _match_key_qbytes_1_T_1 ? phv_data_247 : _GEN_2047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2049 = 8'hf8 == _match_key_qbytes_1_T_1 ? phv_data_248 : _GEN_2048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2050 = 8'hf9 == _match_key_qbytes_1_T_1 ? phv_data_249 : _GEN_2049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2051 = 8'hfa == _match_key_qbytes_1_T_1 ? phv_data_250 : _GEN_2050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2052 = 8'hfb == _match_key_qbytes_1_T_1 ? phv_data_251 : _GEN_2051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2053 = 8'hfc == _match_key_qbytes_1_T_1 ? phv_data_252 : _GEN_2052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2054 = 8'hfd == _match_key_qbytes_1_T_1 ? phv_data_253 : _GEN_2053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2055 = 8'hfe == _match_key_qbytes_1_T_1 ? phv_data_254 : _GEN_2054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2056 = 8'hff == _match_key_qbytes_1_T_1 ? phv_data_255 : _GEN_2055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_1_T_3 = {_GEN_1800,_GEN_2056,_GEN_1288,_GEN_1544}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_1 = local_offset_1 < end_offset ? _match_key_qbytes_1_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_2 = 8'h8 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_2_hi = local_offset_2[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_2_T = {match_key_qbytes_2_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_2_T_1 = {match_key_qbytes_2_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_2_T_2 = {match_key_qbytes_2_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2059 = 8'h1 == _match_key_qbytes_2_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2060 = 8'h2 == _match_key_qbytes_2_T_2 ? phv_data_2 : _GEN_2059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2061 = 8'h3 == _match_key_qbytes_2_T_2 ? phv_data_3 : _GEN_2060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2062 = 8'h4 == _match_key_qbytes_2_T_2 ? phv_data_4 : _GEN_2061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2063 = 8'h5 == _match_key_qbytes_2_T_2 ? phv_data_5 : _GEN_2062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2064 = 8'h6 == _match_key_qbytes_2_T_2 ? phv_data_6 : _GEN_2063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2065 = 8'h7 == _match_key_qbytes_2_T_2 ? phv_data_7 : _GEN_2064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2066 = 8'h8 == _match_key_qbytes_2_T_2 ? phv_data_8 : _GEN_2065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2067 = 8'h9 == _match_key_qbytes_2_T_2 ? phv_data_9 : _GEN_2066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2068 = 8'ha == _match_key_qbytes_2_T_2 ? phv_data_10 : _GEN_2067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2069 = 8'hb == _match_key_qbytes_2_T_2 ? phv_data_11 : _GEN_2068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2070 = 8'hc == _match_key_qbytes_2_T_2 ? phv_data_12 : _GEN_2069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2071 = 8'hd == _match_key_qbytes_2_T_2 ? phv_data_13 : _GEN_2070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2072 = 8'he == _match_key_qbytes_2_T_2 ? phv_data_14 : _GEN_2071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2073 = 8'hf == _match_key_qbytes_2_T_2 ? phv_data_15 : _GEN_2072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2074 = 8'h10 == _match_key_qbytes_2_T_2 ? phv_data_16 : _GEN_2073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2075 = 8'h11 == _match_key_qbytes_2_T_2 ? phv_data_17 : _GEN_2074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2076 = 8'h12 == _match_key_qbytes_2_T_2 ? phv_data_18 : _GEN_2075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2077 = 8'h13 == _match_key_qbytes_2_T_2 ? phv_data_19 : _GEN_2076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2078 = 8'h14 == _match_key_qbytes_2_T_2 ? phv_data_20 : _GEN_2077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2079 = 8'h15 == _match_key_qbytes_2_T_2 ? phv_data_21 : _GEN_2078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2080 = 8'h16 == _match_key_qbytes_2_T_2 ? phv_data_22 : _GEN_2079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2081 = 8'h17 == _match_key_qbytes_2_T_2 ? phv_data_23 : _GEN_2080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2082 = 8'h18 == _match_key_qbytes_2_T_2 ? phv_data_24 : _GEN_2081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2083 = 8'h19 == _match_key_qbytes_2_T_2 ? phv_data_25 : _GEN_2082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2084 = 8'h1a == _match_key_qbytes_2_T_2 ? phv_data_26 : _GEN_2083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2085 = 8'h1b == _match_key_qbytes_2_T_2 ? phv_data_27 : _GEN_2084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2086 = 8'h1c == _match_key_qbytes_2_T_2 ? phv_data_28 : _GEN_2085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2087 = 8'h1d == _match_key_qbytes_2_T_2 ? phv_data_29 : _GEN_2086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2088 = 8'h1e == _match_key_qbytes_2_T_2 ? phv_data_30 : _GEN_2087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2089 = 8'h1f == _match_key_qbytes_2_T_2 ? phv_data_31 : _GEN_2088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2090 = 8'h20 == _match_key_qbytes_2_T_2 ? phv_data_32 : _GEN_2089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2091 = 8'h21 == _match_key_qbytes_2_T_2 ? phv_data_33 : _GEN_2090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2092 = 8'h22 == _match_key_qbytes_2_T_2 ? phv_data_34 : _GEN_2091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2093 = 8'h23 == _match_key_qbytes_2_T_2 ? phv_data_35 : _GEN_2092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2094 = 8'h24 == _match_key_qbytes_2_T_2 ? phv_data_36 : _GEN_2093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2095 = 8'h25 == _match_key_qbytes_2_T_2 ? phv_data_37 : _GEN_2094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2096 = 8'h26 == _match_key_qbytes_2_T_2 ? phv_data_38 : _GEN_2095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2097 = 8'h27 == _match_key_qbytes_2_T_2 ? phv_data_39 : _GEN_2096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2098 = 8'h28 == _match_key_qbytes_2_T_2 ? phv_data_40 : _GEN_2097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2099 = 8'h29 == _match_key_qbytes_2_T_2 ? phv_data_41 : _GEN_2098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2100 = 8'h2a == _match_key_qbytes_2_T_2 ? phv_data_42 : _GEN_2099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2101 = 8'h2b == _match_key_qbytes_2_T_2 ? phv_data_43 : _GEN_2100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2102 = 8'h2c == _match_key_qbytes_2_T_2 ? phv_data_44 : _GEN_2101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2103 = 8'h2d == _match_key_qbytes_2_T_2 ? phv_data_45 : _GEN_2102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2104 = 8'h2e == _match_key_qbytes_2_T_2 ? phv_data_46 : _GEN_2103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2105 = 8'h2f == _match_key_qbytes_2_T_2 ? phv_data_47 : _GEN_2104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2106 = 8'h30 == _match_key_qbytes_2_T_2 ? phv_data_48 : _GEN_2105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2107 = 8'h31 == _match_key_qbytes_2_T_2 ? phv_data_49 : _GEN_2106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2108 = 8'h32 == _match_key_qbytes_2_T_2 ? phv_data_50 : _GEN_2107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2109 = 8'h33 == _match_key_qbytes_2_T_2 ? phv_data_51 : _GEN_2108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2110 = 8'h34 == _match_key_qbytes_2_T_2 ? phv_data_52 : _GEN_2109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2111 = 8'h35 == _match_key_qbytes_2_T_2 ? phv_data_53 : _GEN_2110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2112 = 8'h36 == _match_key_qbytes_2_T_2 ? phv_data_54 : _GEN_2111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2113 = 8'h37 == _match_key_qbytes_2_T_2 ? phv_data_55 : _GEN_2112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2114 = 8'h38 == _match_key_qbytes_2_T_2 ? phv_data_56 : _GEN_2113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2115 = 8'h39 == _match_key_qbytes_2_T_2 ? phv_data_57 : _GEN_2114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2116 = 8'h3a == _match_key_qbytes_2_T_2 ? phv_data_58 : _GEN_2115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2117 = 8'h3b == _match_key_qbytes_2_T_2 ? phv_data_59 : _GEN_2116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2118 = 8'h3c == _match_key_qbytes_2_T_2 ? phv_data_60 : _GEN_2117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2119 = 8'h3d == _match_key_qbytes_2_T_2 ? phv_data_61 : _GEN_2118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2120 = 8'h3e == _match_key_qbytes_2_T_2 ? phv_data_62 : _GEN_2119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2121 = 8'h3f == _match_key_qbytes_2_T_2 ? phv_data_63 : _GEN_2120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2122 = 8'h40 == _match_key_qbytes_2_T_2 ? phv_data_64 : _GEN_2121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2123 = 8'h41 == _match_key_qbytes_2_T_2 ? phv_data_65 : _GEN_2122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2124 = 8'h42 == _match_key_qbytes_2_T_2 ? phv_data_66 : _GEN_2123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2125 = 8'h43 == _match_key_qbytes_2_T_2 ? phv_data_67 : _GEN_2124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2126 = 8'h44 == _match_key_qbytes_2_T_2 ? phv_data_68 : _GEN_2125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2127 = 8'h45 == _match_key_qbytes_2_T_2 ? phv_data_69 : _GEN_2126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2128 = 8'h46 == _match_key_qbytes_2_T_2 ? phv_data_70 : _GEN_2127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2129 = 8'h47 == _match_key_qbytes_2_T_2 ? phv_data_71 : _GEN_2128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2130 = 8'h48 == _match_key_qbytes_2_T_2 ? phv_data_72 : _GEN_2129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2131 = 8'h49 == _match_key_qbytes_2_T_2 ? phv_data_73 : _GEN_2130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2132 = 8'h4a == _match_key_qbytes_2_T_2 ? phv_data_74 : _GEN_2131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2133 = 8'h4b == _match_key_qbytes_2_T_2 ? phv_data_75 : _GEN_2132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2134 = 8'h4c == _match_key_qbytes_2_T_2 ? phv_data_76 : _GEN_2133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2135 = 8'h4d == _match_key_qbytes_2_T_2 ? phv_data_77 : _GEN_2134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2136 = 8'h4e == _match_key_qbytes_2_T_2 ? phv_data_78 : _GEN_2135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2137 = 8'h4f == _match_key_qbytes_2_T_2 ? phv_data_79 : _GEN_2136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2138 = 8'h50 == _match_key_qbytes_2_T_2 ? phv_data_80 : _GEN_2137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2139 = 8'h51 == _match_key_qbytes_2_T_2 ? phv_data_81 : _GEN_2138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2140 = 8'h52 == _match_key_qbytes_2_T_2 ? phv_data_82 : _GEN_2139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2141 = 8'h53 == _match_key_qbytes_2_T_2 ? phv_data_83 : _GEN_2140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2142 = 8'h54 == _match_key_qbytes_2_T_2 ? phv_data_84 : _GEN_2141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2143 = 8'h55 == _match_key_qbytes_2_T_2 ? phv_data_85 : _GEN_2142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2144 = 8'h56 == _match_key_qbytes_2_T_2 ? phv_data_86 : _GEN_2143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2145 = 8'h57 == _match_key_qbytes_2_T_2 ? phv_data_87 : _GEN_2144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2146 = 8'h58 == _match_key_qbytes_2_T_2 ? phv_data_88 : _GEN_2145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2147 = 8'h59 == _match_key_qbytes_2_T_2 ? phv_data_89 : _GEN_2146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2148 = 8'h5a == _match_key_qbytes_2_T_2 ? phv_data_90 : _GEN_2147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2149 = 8'h5b == _match_key_qbytes_2_T_2 ? phv_data_91 : _GEN_2148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2150 = 8'h5c == _match_key_qbytes_2_T_2 ? phv_data_92 : _GEN_2149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2151 = 8'h5d == _match_key_qbytes_2_T_2 ? phv_data_93 : _GEN_2150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2152 = 8'h5e == _match_key_qbytes_2_T_2 ? phv_data_94 : _GEN_2151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2153 = 8'h5f == _match_key_qbytes_2_T_2 ? phv_data_95 : _GEN_2152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2154 = 8'h60 == _match_key_qbytes_2_T_2 ? phv_data_96 : _GEN_2153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2155 = 8'h61 == _match_key_qbytes_2_T_2 ? phv_data_97 : _GEN_2154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2156 = 8'h62 == _match_key_qbytes_2_T_2 ? phv_data_98 : _GEN_2155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2157 = 8'h63 == _match_key_qbytes_2_T_2 ? phv_data_99 : _GEN_2156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2158 = 8'h64 == _match_key_qbytes_2_T_2 ? phv_data_100 : _GEN_2157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2159 = 8'h65 == _match_key_qbytes_2_T_2 ? phv_data_101 : _GEN_2158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2160 = 8'h66 == _match_key_qbytes_2_T_2 ? phv_data_102 : _GEN_2159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2161 = 8'h67 == _match_key_qbytes_2_T_2 ? phv_data_103 : _GEN_2160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2162 = 8'h68 == _match_key_qbytes_2_T_2 ? phv_data_104 : _GEN_2161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2163 = 8'h69 == _match_key_qbytes_2_T_2 ? phv_data_105 : _GEN_2162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2164 = 8'h6a == _match_key_qbytes_2_T_2 ? phv_data_106 : _GEN_2163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2165 = 8'h6b == _match_key_qbytes_2_T_2 ? phv_data_107 : _GEN_2164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2166 = 8'h6c == _match_key_qbytes_2_T_2 ? phv_data_108 : _GEN_2165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2167 = 8'h6d == _match_key_qbytes_2_T_2 ? phv_data_109 : _GEN_2166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2168 = 8'h6e == _match_key_qbytes_2_T_2 ? phv_data_110 : _GEN_2167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2169 = 8'h6f == _match_key_qbytes_2_T_2 ? phv_data_111 : _GEN_2168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2170 = 8'h70 == _match_key_qbytes_2_T_2 ? phv_data_112 : _GEN_2169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2171 = 8'h71 == _match_key_qbytes_2_T_2 ? phv_data_113 : _GEN_2170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2172 = 8'h72 == _match_key_qbytes_2_T_2 ? phv_data_114 : _GEN_2171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2173 = 8'h73 == _match_key_qbytes_2_T_2 ? phv_data_115 : _GEN_2172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2174 = 8'h74 == _match_key_qbytes_2_T_2 ? phv_data_116 : _GEN_2173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2175 = 8'h75 == _match_key_qbytes_2_T_2 ? phv_data_117 : _GEN_2174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2176 = 8'h76 == _match_key_qbytes_2_T_2 ? phv_data_118 : _GEN_2175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2177 = 8'h77 == _match_key_qbytes_2_T_2 ? phv_data_119 : _GEN_2176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2178 = 8'h78 == _match_key_qbytes_2_T_2 ? phv_data_120 : _GEN_2177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2179 = 8'h79 == _match_key_qbytes_2_T_2 ? phv_data_121 : _GEN_2178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2180 = 8'h7a == _match_key_qbytes_2_T_2 ? phv_data_122 : _GEN_2179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2181 = 8'h7b == _match_key_qbytes_2_T_2 ? phv_data_123 : _GEN_2180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2182 = 8'h7c == _match_key_qbytes_2_T_2 ? phv_data_124 : _GEN_2181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2183 = 8'h7d == _match_key_qbytes_2_T_2 ? phv_data_125 : _GEN_2182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2184 = 8'h7e == _match_key_qbytes_2_T_2 ? phv_data_126 : _GEN_2183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2185 = 8'h7f == _match_key_qbytes_2_T_2 ? phv_data_127 : _GEN_2184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2186 = 8'h80 == _match_key_qbytes_2_T_2 ? phv_data_128 : _GEN_2185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2187 = 8'h81 == _match_key_qbytes_2_T_2 ? phv_data_129 : _GEN_2186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2188 = 8'h82 == _match_key_qbytes_2_T_2 ? phv_data_130 : _GEN_2187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2189 = 8'h83 == _match_key_qbytes_2_T_2 ? phv_data_131 : _GEN_2188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2190 = 8'h84 == _match_key_qbytes_2_T_2 ? phv_data_132 : _GEN_2189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2191 = 8'h85 == _match_key_qbytes_2_T_2 ? phv_data_133 : _GEN_2190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2192 = 8'h86 == _match_key_qbytes_2_T_2 ? phv_data_134 : _GEN_2191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2193 = 8'h87 == _match_key_qbytes_2_T_2 ? phv_data_135 : _GEN_2192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2194 = 8'h88 == _match_key_qbytes_2_T_2 ? phv_data_136 : _GEN_2193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2195 = 8'h89 == _match_key_qbytes_2_T_2 ? phv_data_137 : _GEN_2194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2196 = 8'h8a == _match_key_qbytes_2_T_2 ? phv_data_138 : _GEN_2195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2197 = 8'h8b == _match_key_qbytes_2_T_2 ? phv_data_139 : _GEN_2196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2198 = 8'h8c == _match_key_qbytes_2_T_2 ? phv_data_140 : _GEN_2197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2199 = 8'h8d == _match_key_qbytes_2_T_2 ? phv_data_141 : _GEN_2198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2200 = 8'h8e == _match_key_qbytes_2_T_2 ? phv_data_142 : _GEN_2199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2201 = 8'h8f == _match_key_qbytes_2_T_2 ? phv_data_143 : _GEN_2200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2202 = 8'h90 == _match_key_qbytes_2_T_2 ? phv_data_144 : _GEN_2201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2203 = 8'h91 == _match_key_qbytes_2_T_2 ? phv_data_145 : _GEN_2202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2204 = 8'h92 == _match_key_qbytes_2_T_2 ? phv_data_146 : _GEN_2203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2205 = 8'h93 == _match_key_qbytes_2_T_2 ? phv_data_147 : _GEN_2204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2206 = 8'h94 == _match_key_qbytes_2_T_2 ? phv_data_148 : _GEN_2205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2207 = 8'h95 == _match_key_qbytes_2_T_2 ? phv_data_149 : _GEN_2206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2208 = 8'h96 == _match_key_qbytes_2_T_2 ? phv_data_150 : _GEN_2207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2209 = 8'h97 == _match_key_qbytes_2_T_2 ? phv_data_151 : _GEN_2208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2210 = 8'h98 == _match_key_qbytes_2_T_2 ? phv_data_152 : _GEN_2209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2211 = 8'h99 == _match_key_qbytes_2_T_2 ? phv_data_153 : _GEN_2210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2212 = 8'h9a == _match_key_qbytes_2_T_2 ? phv_data_154 : _GEN_2211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2213 = 8'h9b == _match_key_qbytes_2_T_2 ? phv_data_155 : _GEN_2212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2214 = 8'h9c == _match_key_qbytes_2_T_2 ? phv_data_156 : _GEN_2213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2215 = 8'h9d == _match_key_qbytes_2_T_2 ? phv_data_157 : _GEN_2214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2216 = 8'h9e == _match_key_qbytes_2_T_2 ? phv_data_158 : _GEN_2215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2217 = 8'h9f == _match_key_qbytes_2_T_2 ? phv_data_159 : _GEN_2216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2218 = 8'ha0 == _match_key_qbytes_2_T_2 ? phv_data_160 : _GEN_2217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2219 = 8'ha1 == _match_key_qbytes_2_T_2 ? phv_data_161 : _GEN_2218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2220 = 8'ha2 == _match_key_qbytes_2_T_2 ? phv_data_162 : _GEN_2219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2221 = 8'ha3 == _match_key_qbytes_2_T_2 ? phv_data_163 : _GEN_2220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2222 = 8'ha4 == _match_key_qbytes_2_T_2 ? phv_data_164 : _GEN_2221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2223 = 8'ha5 == _match_key_qbytes_2_T_2 ? phv_data_165 : _GEN_2222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2224 = 8'ha6 == _match_key_qbytes_2_T_2 ? phv_data_166 : _GEN_2223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2225 = 8'ha7 == _match_key_qbytes_2_T_2 ? phv_data_167 : _GEN_2224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2226 = 8'ha8 == _match_key_qbytes_2_T_2 ? phv_data_168 : _GEN_2225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2227 = 8'ha9 == _match_key_qbytes_2_T_2 ? phv_data_169 : _GEN_2226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2228 = 8'haa == _match_key_qbytes_2_T_2 ? phv_data_170 : _GEN_2227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2229 = 8'hab == _match_key_qbytes_2_T_2 ? phv_data_171 : _GEN_2228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2230 = 8'hac == _match_key_qbytes_2_T_2 ? phv_data_172 : _GEN_2229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2231 = 8'had == _match_key_qbytes_2_T_2 ? phv_data_173 : _GEN_2230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2232 = 8'hae == _match_key_qbytes_2_T_2 ? phv_data_174 : _GEN_2231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2233 = 8'haf == _match_key_qbytes_2_T_2 ? phv_data_175 : _GEN_2232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2234 = 8'hb0 == _match_key_qbytes_2_T_2 ? phv_data_176 : _GEN_2233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2235 = 8'hb1 == _match_key_qbytes_2_T_2 ? phv_data_177 : _GEN_2234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2236 = 8'hb2 == _match_key_qbytes_2_T_2 ? phv_data_178 : _GEN_2235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2237 = 8'hb3 == _match_key_qbytes_2_T_2 ? phv_data_179 : _GEN_2236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2238 = 8'hb4 == _match_key_qbytes_2_T_2 ? phv_data_180 : _GEN_2237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2239 = 8'hb5 == _match_key_qbytes_2_T_2 ? phv_data_181 : _GEN_2238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2240 = 8'hb6 == _match_key_qbytes_2_T_2 ? phv_data_182 : _GEN_2239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2241 = 8'hb7 == _match_key_qbytes_2_T_2 ? phv_data_183 : _GEN_2240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2242 = 8'hb8 == _match_key_qbytes_2_T_2 ? phv_data_184 : _GEN_2241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2243 = 8'hb9 == _match_key_qbytes_2_T_2 ? phv_data_185 : _GEN_2242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2244 = 8'hba == _match_key_qbytes_2_T_2 ? phv_data_186 : _GEN_2243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2245 = 8'hbb == _match_key_qbytes_2_T_2 ? phv_data_187 : _GEN_2244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2246 = 8'hbc == _match_key_qbytes_2_T_2 ? phv_data_188 : _GEN_2245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2247 = 8'hbd == _match_key_qbytes_2_T_2 ? phv_data_189 : _GEN_2246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2248 = 8'hbe == _match_key_qbytes_2_T_2 ? phv_data_190 : _GEN_2247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2249 = 8'hbf == _match_key_qbytes_2_T_2 ? phv_data_191 : _GEN_2248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2250 = 8'hc0 == _match_key_qbytes_2_T_2 ? phv_data_192 : _GEN_2249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2251 = 8'hc1 == _match_key_qbytes_2_T_2 ? phv_data_193 : _GEN_2250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2252 = 8'hc2 == _match_key_qbytes_2_T_2 ? phv_data_194 : _GEN_2251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2253 = 8'hc3 == _match_key_qbytes_2_T_2 ? phv_data_195 : _GEN_2252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2254 = 8'hc4 == _match_key_qbytes_2_T_2 ? phv_data_196 : _GEN_2253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2255 = 8'hc5 == _match_key_qbytes_2_T_2 ? phv_data_197 : _GEN_2254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2256 = 8'hc6 == _match_key_qbytes_2_T_2 ? phv_data_198 : _GEN_2255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2257 = 8'hc7 == _match_key_qbytes_2_T_2 ? phv_data_199 : _GEN_2256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2258 = 8'hc8 == _match_key_qbytes_2_T_2 ? phv_data_200 : _GEN_2257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2259 = 8'hc9 == _match_key_qbytes_2_T_2 ? phv_data_201 : _GEN_2258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2260 = 8'hca == _match_key_qbytes_2_T_2 ? phv_data_202 : _GEN_2259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2261 = 8'hcb == _match_key_qbytes_2_T_2 ? phv_data_203 : _GEN_2260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2262 = 8'hcc == _match_key_qbytes_2_T_2 ? phv_data_204 : _GEN_2261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2263 = 8'hcd == _match_key_qbytes_2_T_2 ? phv_data_205 : _GEN_2262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2264 = 8'hce == _match_key_qbytes_2_T_2 ? phv_data_206 : _GEN_2263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2265 = 8'hcf == _match_key_qbytes_2_T_2 ? phv_data_207 : _GEN_2264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2266 = 8'hd0 == _match_key_qbytes_2_T_2 ? phv_data_208 : _GEN_2265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2267 = 8'hd1 == _match_key_qbytes_2_T_2 ? phv_data_209 : _GEN_2266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2268 = 8'hd2 == _match_key_qbytes_2_T_2 ? phv_data_210 : _GEN_2267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2269 = 8'hd3 == _match_key_qbytes_2_T_2 ? phv_data_211 : _GEN_2268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2270 = 8'hd4 == _match_key_qbytes_2_T_2 ? phv_data_212 : _GEN_2269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2271 = 8'hd5 == _match_key_qbytes_2_T_2 ? phv_data_213 : _GEN_2270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2272 = 8'hd6 == _match_key_qbytes_2_T_2 ? phv_data_214 : _GEN_2271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2273 = 8'hd7 == _match_key_qbytes_2_T_2 ? phv_data_215 : _GEN_2272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2274 = 8'hd8 == _match_key_qbytes_2_T_2 ? phv_data_216 : _GEN_2273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2275 = 8'hd9 == _match_key_qbytes_2_T_2 ? phv_data_217 : _GEN_2274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2276 = 8'hda == _match_key_qbytes_2_T_2 ? phv_data_218 : _GEN_2275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2277 = 8'hdb == _match_key_qbytes_2_T_2 ? phv_data_219 : _GEN_2276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2278 = 8'hdc == _match_key_qbytes_2_T_2 ? phv_data_220 : _GEN_2277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2279 = 8'hdd == _match_key_qbytes_2_T_2 ? phv_data_221 : _GEN_2278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2280 = 8'hde == _match_key_qbytes_2_T_2 ? phv_data_222 : _GEN_2279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2281 = 8'hdf == _match_key_qbytes_2_T_2 ? phv_data_223 : _GEN_2280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2282 = 8'he0 == _match_key_qbytes_2_T_2 ? phv_data_224 : _GEN_2281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2283 = 8'he1 == _match_key_qbytes_2_T_2 ? phv_data_225 : _GEN_2282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2284 = 8'he2 == _match_key_qbytes_2_T_2 ? phv_data_226 : _GEN_2283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2285 = 8'he3 == _match_key_qbytes_2_T_2 ? phv_data_227 : _GEN_2284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2286 = 8'he4 == _match_key_qbytes_2_T_2 ? phv_data_228 : _GEN_2285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2287 = 8'he5 == _match_key_qbytes_2_T_2 ? phv_data_229 : _GEN_2286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2288 = 8'he6 == _match_key_qbytes_2_T_2 ? phv_data_230 : _GEN_2287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2289 = 8'he7 == _match_key_qbytes_2_T_2 ? phv_data_231 : _GEN_2288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2290 = 8'he8 == _match_key_qbytes_2_T_2 ? phv_data_232 : _GEN_2289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2291 = 8'he9 == _match_key_qbytes_2_T_2 ? phv_data_233 : _GEN_2290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2292 = 8'hea == _match_key_qbytes_2_T_2 ? phv_data_234 : _GEN_2291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2293 = 8'heb == _match_key_qbytes_2_T_2 ? phv_data_235 : _GEN_2292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2294 = 8'hec == _match_key_qbytes_2_T_2 ? phv_data_236 : _GEN_2293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2295 = 8'hed == _match_key_qbytes_2_T_2 ? phv_data_237 : _GEN_2294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2296 = 8'hee == _match_key_qbytes_2_T_2 ? phv_data_238 : _GEN_2295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2297 = 8'hef == _match_key_qbytes_2_T_2 ? phv_data_239 : _GEN_2296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2298 = 8'hf0 == _match_key_qbytes_2_T_2 ? phv_data_240 : _GEN_2297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2299 = 8'hf1 == _match_key_qbytes_2_T_2 ? phv_data_241 : _GEN_2298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2300 = 8'hf2 == _match_key_qbytes_2_T_2 ? phv_data_242 : _GEN_2299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2301 = 8'hf3 == _match_key_qbytes_2_T_2 ? phv_data_243 : _GEN_2300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2302 = 8'hf4 == _match_key_qbytes_2_T_2 ? phv_data_244 : _GEN_2301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2303 = 8'hf5 == _match_key_qbytes_2_T_2 ? phv_data_245 : _GEN_2302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2304 = 8'hf6 == _match_key_qbytes_2_T_2 ? phv_data_246 : _GEN_2303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2305 = 8'hf7 == _match_key_qbytes_2_T_2 ? phv_data_247 : _GEN_2304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2306 = 8'hf8 == _match_key_qbytes_2_T_2 ? phv_data_248 : _GEN_2305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2307 = 8'hf9 == _match_key_qbytes_2_T_2 ? phv_data_249 : _GEN_2306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2308 = 8'hfa == _match_key_qbytes_2_T_2 ? phv_data_250 : _GEN_2307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2309 = 8'hfb == _match_key_qbytes_2_T_2 ? phv_data_251 : _GEN_2308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2310 = 8'hfc == _match_key_qbytes_2_T_2 ? phv_data_252 : _GEN_2309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2311 = 8'hfd == _match_key_qbytes_2_T_2 ? phv_data_253 : _GEN_2310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2312 = 8'hfe == _match_key_qbytes_2_T_2 ? phv_data_254 : _GEN_2311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2313 = 8'hff == _match_key_qbytes_2_T_2 ? phv_data_255 : _GEN_2312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2315 = 8'h1 == local_offset_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2316 = 8'h2 == local_offset_2 ? phv_data_2 : _GEN_2315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2317 = 8'h3 == local_offset_2 ? phv_data_3 : _GEN_2316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2318 = 8'h4 == local_offset_2 ? phv_data_4 : _GEN_2317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2319 = 8'h5 == local_offset_2 ? phv_data_5 : _GEN_2318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2320 = 8'h6 == local_offset_2 ? phv_data_6 : _GEN_2319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2321 = 8'h7 == local_offset_2 ? phv_data_7 : _GEN_2320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2322 = 8'h8 == local_offset_2 ? phv_data_8 : _GEN_2321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2323 = 8'h9 == local_offset_2 ? phv_data_9 : _GEN_2322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2324 = 8'ha == local_offset_2 ? phv_data_10 : _GEN_2323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2325 = 8'hb == local_offset_2 ? phv_data_11 : _GEN_2324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2326 = 8'hc == local_offset_2 ? phv_data_12 : _GEN_2325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2327 = 8'hd == local_offset_2 ? phv_data_13 : _GEN_2326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2328 = 8'he == local_offset_2 ? phv_data_14 : _GEN_2327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2329 = 8'hf == local_offset_2 ? phv_data_15 : _GEN_2328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2330 = 8'h10 == local_offset_2 ? phv_data_16 : _GEN_2329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2331 = 8'h11 == local_offset_2 ? phv_data_17 : _GEN_2330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2332 = 8'h12 == local_offset_2 ? phv_data_18 : _GEN_2331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2333 = 8'h13 == local_offset_2 ? phv_data_19 : _GEN_2332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2334 = 8'h14 == local_offset_2 ? phv_data_20 : _GEN_2333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2335 = 8'h15 == local_offset_2 ? phv_data_21 : _GEN_2334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2336 = 8'h16 == local_offset_2 ? phv_data_22 : _GEN_2335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2337 = 8'h17 == local_offset_2 ? phv_data_23 : _GEN_2336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2338 = 8'h18 == local_offset_2 ? phv_data_24 : _GEN_2337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2339 = 8'h19 == local_offset_2 ? phv_data_25 : _GEN_2338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2340 = 8'h1a == local_offset_2 ? phv_data_26 : _GEN_2339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2341 = 8'h1b == local_offset_2 ? phv_data_27 : _GEN_2340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2342 = 8'h1c == local_offset_2 ? phv_data_28 : _GEN_2341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2343 = 8'h1d == local_offset_2 ? phv_data_29 : _GEN_2342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2344 = 8'h1e == local_offset_2 ? phv_data_30 : _GEN_2343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2345 = 8'h1f == local_offset_2 ? phv_data_31 : _GEN_2344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2346 = 8'h20 == local_offset_2 ? phv_data_32 : _GEN_2345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2347 = 8'h21 == local_offset_2 ? phv_data_33 : _GEN_2346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2348 = 8'h22 == local_offset_2 ? phv_data_34 : _GEN_2347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2349 = 8'h23 == local_offset_2 ? phv_data_35 : _GEN_2348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2350 = 8'h24 == local_offset_2 ? phv_data_36 : _GEN_2349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2351 = 8'h25 == local_offset_2 ? phv_data_37 : _GEN_2350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2352 = 8'h26 == local_offset_2 ? phv_data_38 : _GEN_2351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2353 = 8'h27 == local_offset_2 ? phv_data_39 : _GEN_2352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2354 = 8'h28 == local_offset_2 ? phv_data_40 : _GEN_2353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2355 = 8'h29 == local_offset_2 ? phv_data_41 : _GEN_2354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2356 = 8'h2a == local_offset_2 ? phv_data_42 : _GEN_2355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2357 = 8'h2b == local_offset_2 ? phv_data_43 : _GEN_2356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2358 = 8'h2c == local_offset_2 ? phv_data_44 : _GEN_2357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2359 = 8'h2d == local_offset_2 ? phv_data_45 : _GEN_2358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2360 = 8'h2e == local_offset_2 ? phv_data_46 : _GEN_2359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2361 = 8'h2f == local_offset_2 ? phv_data_47 : _GEN_2360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2362 = 8'h30 == local_offset_2 ? phv_data_48 : _GEN_2361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2363 = 8'h31 == local_offset_2 ? phv_data_49 : _GEN_2362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2364 = 8'h32 == local_offset_2 ? phv_data_50 : _GEN_2363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2365 = 8'h33 == local_offset_2 ? phv_data_51 : _GEN_2364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2366 = 8'h34 == local_offset_2 ? phv_data_52 : _GEN_2365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2367 = 8'h35 == local_offset_2 ? phv_data_53 : _GEN_2366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2368 = 8'h36 == local_offset_2 ? phv_data_54 : _GEN_2367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2369 = 8'h37 == local_offset_2 ? phv_data_55 : _GEN_2368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2370 = 8'h38 == local_offset_2 ? phv_data_56 : _GEN_2369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2371 = 8'h39 == local_offset_2 ? phv_data_57 : _GEN_2370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2372 = 8'h3a == local_offset_2 ? phv_data_58 : _GEN_2371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2373 = 8'h3b == local_offset_2 ? phv_data_59 : _GEN_2372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2374 = 8'h3c == local_offset_2 ? phv_data_60 : _GEN_2373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2375 = 8'h3d == local_offset_2 ? phv_data_61 : _GEN_2374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2376 = 8'h3e == local_offset_2 ? phv_data_62 : _GEN_2375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2377 = 8'h3f == local_offset_2 ? phv_data_63 : _GEN_2376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2378 = 8'h40 == local_offset_2 ? phv_data_64 : _GEN_2377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2379 = 8'h41 == local_offset_2 ? phv_data_65 : _GEN_2378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2380 = 8'h42 == local_offset_2 ? phv_data_66 : _GEN_2379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2381 = 8'h43 == local_offset_2 ? phv_data_67 : _GEN_2380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2382 = 8'h44 == local_offset_2 ? phv_data_68 : _GEN_2381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2383 = 8'h45 == local_offset_2 ? phv_data_69 : _GEN_2382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2384 = 8'h46 == local_offset_2 ? phv_data_70 : _GEN_2383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2385 = 8'h47 == local_offset_2 ? phv_data_71 : _GEN_2384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2386 = 8'h48 == local_offset_2 ? phv_data_72 : _GEN_2385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2387 = 8'h49 == local_offset_2 ? phv_data_73 : _GEN_2386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2388 = 8'h4a == local_offset_2 ? phv_data_74 : _GEN_2387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2389 = 8'h4b == local_offset_2 ? phv_data_75 : _GEN_2388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2390 = 8'h4c == local_offset_2 ? phv_data_76 : _GEN_2389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2391 = 8'h4d == local_offset_2 ? phv_data_77 : _GEN_2390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2392 = 8'h4e == local_offset_2 ? phv_data_78 : _GEN_2391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2393 = 8'h4f == local_offset_2 ? phv_data_79 : _GEN_2392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2394 = 8'h50 == local_offset_2 ? phv_data_80 : _GEN_2393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2395 = 8'h51 == local_offset_2 ? phv_data_81 : _GEN_2394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2396 = 8'h52 == local_offset_2 ? phv_data_82 : _GEN_2395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2397 = 8'h53 == local_offset_2 ? phv_data_83 : _GEN_2396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2398 = 8'h54 == local_offset_2 ? phv_data_84 : _GEN_2397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2399 = 8'h55 == local_offset_2 ? phv_data_85 : _GEN_2398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2400 = 8'h56 == local_offset_2 ? phv_data_86 : _GEN_2399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2401 = 8'h57 == local_offset_2 ? phv_data_87 : _GEN_2400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2402 = 8'h58 == local_offset_2 ? phv_data_88 : _GEN_2401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2403 = 8'h59 == local_offset_2 ? phv_data_89 : _GEN_2402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2404 = 8'h5a == local_offset_2 ? phv_data_90 : _GEN_2403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2405 = 8'h5b == local_offset_2 ? phv_data_91 : _GEN_2404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2406 = 8'h5c == local_offset_2 ? phv_data_92 : _GEN_2405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2407 = 8'h5d == local_offset_2 ? phv_data_93 : _GEN_2406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2408 = 8'h5e == local_offset_2 ? phv_data_94 : _GEN_2407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2409 = 8'h5f == local_offset_2 ? phv_data_95 : _GEN_2408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2410 = 8'h60 == local_offset_2 ? phv_data_96 : _GEN_2409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2411 = 8'h61 == local_offset_2 ? phv_data_97 : _GEN_2410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2412 = 8'h62 == local_offset_2 ? phv_data_98 : _GEN_2411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2413 = 8'h63 == local_offset_2 ? phv_data_99 : _GEN_2412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2414 = 8'h64 == local_offset_2 ? phv_data_100 : _GEN_2413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2415 = 8'h65 == local_offset_2 ? phv_data_101 : _GEN_2414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2416 = 8'h66 == local_offset_2 ? phv_data_102 : _GEN_2415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2417 = 8'h67 == local_offset_2 ? phv_data_103 : _GEN_2416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2418 = 8'h68 == local_offset_2 ? phv_data_104 : _GEN_2417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2419 = 8'h69 == local_offset_2 ? phv_data_105 : _GEN_2418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2420 = 8'h6a == local_offset_2 ? phv_data_106 : _GEN_2419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2421 = 8'h6b == local_offset_2 ? phv_data_107 : _GEN_2420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2422 = 8'h6c == local_offset_2 ? phv_data_108 : _GEN_2421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2423 = 8'h6d == local_offset_2 ? phv_data_109 : _GEN_2422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2424 = 8'h6e == local_offset_2 ? phv_data_110 : _GEN_2423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2425 = 8'h6f == local_offset_2 ? phv_data_111 : _GEN_2424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2426 = 8'h70 == local_offset_2 ? phv_data_112 : _GEN_2425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2427 = 8'h71 == local_offset_2 ? phv_data_113 : _GEN_2426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2428 = 8'h72 == local_offset_2 ? phv_data_114 : _GEN_2427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2429 = 8'h73 == local_offset_2 ? phv_data_115 : _GEN_2428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2430 = 8'h74 == local_offset_2 ? phv_data_116 : _GEN_2429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2431 = 8'h75 == local_offset_2 ? phv_data_117 : _GEN_2430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2432 = 8'h76 == local_offset_2 ? phv_data_118 : _GEN_2431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2433 = 8'h77 == local_offset_2 ? phv_data_119 : _GEN_2432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2434 = 8'h78 == local_offset_2 ? phv_data_120 : _GEN_2433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2435 = 8'h79 == local_offset_2 ? phv_data_121 : _GEN_2434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2436 = 8'h7a == local_offset_2 ? phv_data_122 : _GEN_2435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2437 = 8'h7b == local_offset_2 ? phv_data_123 : _GEN_2436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2438 = 8'h7c == local_offset_2 ? phv_data_124 : _GEN_2437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2439 = 8'h7d == local_offset_2 ? phv_data_125 : _GEN_2438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2440 = 8'h7e == local_offset_2 ? phv_data_126 : _GEN_2439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2441 = 8'h7f == local_offset_2 ? phv_data_127 : _GEN_2440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2442 = 8'h80 == local_offset_2 ? phv_data_128 : _GEN_2441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2443 = 8'h81 == local_offset_2 ? phv_data_129 : _GEN_2442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2444 = 8'h82 == local_offset_2 ? phv_data_130 : _GEN_2443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2445 = 8'h83 == local_offset_2 ? phv_data_131 : _GEN_2444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2446 = 8'h84 == local_offset_2 ? phv_data_132 : _GEN_2445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2447 = 8'h85 == local_offset_2 ? phv_data_133 : _GEN_2446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2448 = 8'h86 == local_offset_2 ? phv_data_134 : _GEN_2447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2449 = 8'h87 == local_offset_2 ? phv_data_135 : _GEN_2448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2450 = 8'h88 == local_offset_2 ? phv_data_136 : _GEN_2449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2451 = 8'h89 == local_offset_2 ? phv_data_137 : _GEN_2450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2452 = 8'h8a == local_offset_2 ? phv_data_138 : _GEN_2451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2453 = 8'h8b == local_offset_2 ? phv_data_139 : _GEN_2452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2454 = 8'h8c == local_offset_2 ? phv_data_140 : _GEN_2453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2455 = 8'h8d == local_offset_2 ? phv_data_141 : _GEN_2454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2456 = 8'h8e == local_offset_2 ? phv_data_142 : _GEN_2455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2457 = 8'h8f == local_offset_2 ? phv_data_143 : _GEN_2456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2458 = 8'h90 == local_offset_2 ? phv_data_144 : _GEN_2457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2459 = 8'h91 == local_offset_2 ? phv_data_145 : _GEN_2458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2460 = 8'h92 == local_offset_2 ? phv_data_146 : _GEN_2459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2461 = 8'h93 == local_offset_2 ? phv_data_147 : _GEN_2460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2462 = 8'h94 == local_offset_2 ? phv_data_148 : _GEN_2461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2463 = 8'h95 == local_offset_2 ? phv_data_149 : _GEN_2462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2464 = 8'h96 == local_offset_2 ? phv_data_150 : _GEN_2463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2465 = 8'h97 == local_offset_2 ? phv_data_151 : _GEN_2464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2466 = 8'h98 == local_offset_2 ? phv_data_152 : _GEN_2465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2467 = 8'h99 == local_offset_2 ? phv_data_153 : _GEN_2466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2468 = 8'h9a == local_offset_2 ? phv_data_154 : _GEN_2467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2469 = 8'h9b == local_offset_2 ? phv_data_155 : _GEN_2468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2470 = 8'h9c == local_offset_2 ? phv_data_156 : _GEN_2469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2471 = 8'h9d == local_offset_2 ? phv_data_157 : _GEN_2470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2472 = 8'h9e == local_offset_2 ? phv_data_158 : _GEN_2471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2473 = 8'h9f == local_offset_2 ? phv_data_159 : _GEN_2472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2474 = 8'ha0 == local_offset_2 ? phv_data_160 : _GEN_2473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2475 = 8'ha1 == local_offset_2 ? phv_data_161 : _GEN_2474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2476 = 8'ha2 == local_offset_2 ? phv_data_162 : _GEN_2475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2477 = 8'ha3 == local_offset_2 ? phv_data_163 : _GEN_2476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2478 = 8'ha4 == local_offset_2 ? phv_data_164 : _GEN_2477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2479 = 8'ha5 == local_offset_2 ? phv_data_165 : _GEN_2478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2480 = 8'ha6 == local_offset_2 ? phv_data_166 : _GEN_2479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2481 = 8'ha7 == local_offset_2 ? phv_data_167 : _GEN_2480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2482 = 8'ha8 == local_offset_2 ? phv_data_168 : _GEN_2481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2483 = 8'ha9 == local_offset_2 ? phv_data_169 : _GEN_2482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2484 = 8'haa == local_offset_2 ? phv_data_170 : _GEN_2483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2485 = 8'hab == local_offset_2 ? phv_data_171 : _GEN_2484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2486 = 8'hac == local_offset_2 ? phv_data_172 : _GEN_2485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2487 = 8'had == local_offset_2 ? phv_data_173 : _GEN_2486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2488 = 8'hae == local_offset_2 ? phv_data_174 : _GEN_2487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2489 = 8'haf == local_offset_2 ? phv_data_175 : _GEN_2488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2490 = 8'hb0 == local_offset_2 ? phv_data_176 : _GEN_2489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2491 = 8'hb1 == local_offset_2 ? phv_data_177 : _GEN_2490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2492 = 8'hb2 == local_offset_2 ? phv_data_178 : _GEN_2491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2493 = 8'hb3 == local_offset_2 ? phv_data_179 : _GEN_2492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2494 = 8'hb4 == local_offset_2 ? phv_data_180 : _GEN_2493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2495 = 8'hb5 == local_offset_2 ? phv_data_181 : _GEN_2494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2496 = 8'hb6 == local_offset_2 ? phv_data_182 : _GEN_2495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2497 = 8'hb7 == local_offset_2 ? phv_data_183 : _GEN_2496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2498 = 8'hb8 == local_offset_2 ? phv_data_184 : _GEN_2497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2499 = 8'hb9 == local_offset_2 ? phv_data_185 : _GEN_2498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2500 = 8'hba == local_offset_2 ? phv_data_186 : _GEN_2499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2501 = 8'hbb == local_offset_2 ? phv_data_187 : _GEN_2500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2502 = 8'hbc == local_offset_2 ? phv_data_188 : _GEN_2501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2503 = 8'hbd == local_offset_2 ? phv_data_189 : _GEN_2502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2504 = 8'hbe == local_offset_2 ? phv_data_190 : _GEN_2503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2505 = 8'hbf == local_offset_2 ? phv_data_191 : _GEN_2504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2506 = 8'hc0 == local_offset_2 ? phv_data_192 : _GEN_2505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2507 = 8'hc1 == local_offset_2 ? phv_data_193 : _GEN_2506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2508 = 8'hc2 == local_offset_2 ? phv_data_194 : _GEN_2507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2509 = 8'hc3 == local_offset_2 ? phv_data_195 : _GEN_2508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2510 = 8'hc4 == local_offset_2 ? phv_data_196 : _GEN_2509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2511 = 8'hc5 == local_offset_2 ? phv_data_197 : _GEN_2510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2512 = 8'hc6 == local_offset_2 ? phv_data_198 : _GEN_2511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2513 = 8'hc7 == local_offset_2 ? phv_data_199 : _GEN_2512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2514 = 8'hc8 == local_offset_2 ? phv_data_200 : _GEN_2513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2515 = 8'hc9 == local_offset_2 ? phv_data_201 : _GEN_2514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2516 = 8'hca == local_offset_2 ? phv_data_202 : _GEN_2515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2517 = 8'hcb == local_offset_2 ? phv_data_203 : _GEN_2516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2518 = 8'hcc == local_offset_2 ? phv_data_204 : _GEN_2517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2519 = 8'hcd == local_offset_2 ? phv_data_205 : _GEN_2518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2520 = 8'hce == local_offset_2 ? phv_data_206 : _GEN_2519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2521 = 8'hcf == local_offset_2 ? phv_data_207 : _GEN_2520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2522 = 8'hd0 == local_offset_2 ? phv_data_208 : _GEN_2521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2523 = 8'hd1 == local_offset_2 ? phv_data_209 : _GEN_2522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2524 = 8'hd2 == local_offset_2 ? phv_data_210 : _GEN_2523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2525 = 8'hd3 == local_offset_2 ? phv_data_211 : _GEN_2524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2526 = 8'hd4 == local_offset_2 ? phv_data_212 : _GEN_2525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2527 = 8'hd5 == local_offset_2 ? phv_data_213 : _GEN_2526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2528 = 8'hd6 == local_offset_2 ? phv_data_214 : _GEN_2527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2529 = 8'hd7 == local_offset_2 ? phv_data_215 : _GEN_2528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2530 = 8'hd8 == local_offset_2 ? phv_data_216 : _GEN_2529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2531 = 8'hd9 == local_offset_2 ? phv_data_217 : _GEN_2530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2532 = 8'hda == local_offset_2 ? phv_data_218 : _GEN_2531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2533 = 8'hdb == local_offset_2 ? phv_data_219 : _GEN_2532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2534 = 8'hdc == local_offset_2 ? phv_data_220 : _GEN_2533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2535 = 8'hdd == local_offset_2 ? phv_data_221 : _GEN_2534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2536 = 8'hde == local_offset_2 ? phv_data_222 : _GEN_2535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2537 = 8'hdf == local_offset_2 ? phv_data_223 : _GEN_2536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2538 = 8'he0 == local_offset_2 ? phv_data_224 : _GEN_2537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2539 = 8'he1 == local_offset_2 ? phv_data_225 : _GEN_2538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2540 = 8'he2 == local_offset_2 ? phv_data_226 : _GEN_2539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2541 = 8'he3 == local_offset_2 ? phv_data_227 : _GEN_2540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2542 = 8'he4 == local_offset_2 ? phv_data_228 : _GEN_2541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2543 = 8'he5 == local_offset_2 ? phv_data_229 : _GEN_2542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2544 = 8'he6 == local_offset_2 ? phv_data_230 : _GEN_2543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2545 = 8'he7 == local_offset_2 ? phv_data_231 : _GEN_2544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2546 = 8'he8 == local_offset_2 ? phv_data_232 : _GEN_2545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2547 = 8'he9 == local_offset_2 ? phv_data_233 : _GEN_2546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2548 = 8'hea == local_offset_2 ? phv_data_234 : _GEN_2547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2549 = 8'heb == local_offset_2 ? phv_data_235 : _GEN_2548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2550 = 8'hec == local_offset_2 ? phv_data_236 : _GEN_2549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2551 = 8'hed == local_offset_2 ? phv_data_237 : _GEN_2550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2552 = 8'hee == local_offset_2 ? phv_data_238 : _GEN_2551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2553 = 8'hef == local_offset_2 ? phv_data_239 : _GEN_2552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2554 = 8'hf0 == local_offset_2 ? phv_data_240 : _GEN_2553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2555 = 8'hf1 == local_offset_2 ? phv_data_241 : _GEN_2554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2556 = 8'hf2 == local_offset_2 ? phv_data_242 : _GEN_2555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2557 = 8'hf3 == local_offset_2 ? phv_data_243 : _GEN_2556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2558 = 8'hf4 == local_offset_2 ? phv_data_244 : _GEN_2557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2559 = 8'hf5 == local_offset_2 ? phv_data_245 : _GEN_2558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2560 = 8'hf6 == local_offset_2 ? phv_data_246 : _GEN_2559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2561 = 8'hf7 == local_offset_2 ? phv_data_247 : _GEN_2560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2562 = 8'hf8 == local_offset_2 ? phv_data_248 : _GEN_2561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2563 = 8'hf9 == local_offset_2 ? phv_data_249 : _GEN_2562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2564 = 8'hfa == local_offset_2 ? phv_data_250 : _GEN_2563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2565 = 8'hfb == local_offset_2 ? phv_data_251 : _GEN_2564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2566 = 8'hfc == local_offset_2 ? phv_data_252 : _GEN_2565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2567 = 8'hfd == local_offset_2 ? phv_data_253 : _GEN_2566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2568 = 8'hfe == local_offset_2 ? phv_data_254 : _GEN_2567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2569 = 8'hff == local_offset_2 ? phv_data_255 : _GEN_2568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2571 = 8'h1 == _match_key_qbytes_2_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2572 = 8'h2 == _match_key_qbytes_2_T ? phv_data_2 : _GEN_2571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2573 = 8'h3 == _match_key_qbytes_2_T ? phv_data_3 : _GEN_2572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2574 = 8'h4 == _match_key_qbytes_2_T ? phv_data_4 : _GEN_2573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2575 = 8'h5 == _match_key_qbytes_2_T ? phv_data_5 : _GEN_2574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2576 = 8'h6 == _match_key_qbytes_2_T ? phv_data_6 : _GEN_2575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2577 = 8'h7 == _match_key_qbytes_2_T ? phv_data_7 : _GEN_2576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2578 = 8'h8 == _match_key_qbytes_2_T ? phv_data_8 : _GEN_2577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2579 = 8'h9 == _match_key_qbytes_2_T ? phv_data_9 : _GEN_2578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2580 = 8'ha == _match_key_qbytes_2_T ? phv_data_10 : _GEN_2579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2581 = 8'hb == _match_key_qbytes_2_T ? phv_data_11 : _GEN_2580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2582 = 8'hc == _match_key_qbytes_2_T ? phv_data_12 : _GEN_2581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2583 = 8'hd == _match_key_qbytes_2_T ? phv_data_13 : _GEN_2582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2584 = 8'he == _match_key_qbytes_2_T ? phv_data_14 : _GEN_2583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2585 = 8'hf == _match_key_qbytes_2_T ? phv_data_15 : _GEN_2584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2586 = 8'h10 == _match_key_qbytes_2_T ? phv_data_16 : _GEN_2585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2587 = 8'h11 == _match_key_qbytes_2_T ? phv_data_17 : _GEN_2586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2588 = 8'h12 == _match_key_qbytes_2_T ? phv_data_18 : _GEN_2587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2589 = 8'h13 == _match_key_qbytes_2_T ? phv_data_19 : _GEN_2588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2590 = 8'h14 == _match_key_qbytes_2_T ? phv_data_20 : _GEN_2589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2591 = 8'h15 == _match_key_qbytes_2_T ? phv_data_21 : _GEN_2590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2592 = 8'h16 == _match_key_qbytes_2_T ? phv_data_22 : _GEN_2591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2593 = 8'h17 == _match_key_qbytes_2_T ? phv_data_23 : _GEN_2592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2594 = 8'h18 == _match_key_qbytes_2_T ? phv_data_24 : _GEN_2593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2595 = 8'h19 == _match_key_qbytes_2_T ? phv_data_25 : _GEN_2594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2596 = 8'h1a == _match_key_qbytes_2_T ? phv_data_26 : _GEN_2595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2597 = 8'h1b == _match_key_qbytes_2_T ? phv_data_27 : _GEN_2596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2598 = 8'h1c == _match_key_qbytes_2_T ? phv_data_28 : _GEN_2597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2599 = 8'h1d == _match_key_qbytes_2_T ? phv_data_29 : _GEN_2598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2600 = 8'h1e == _match_key_qbytes_2_T ? phv_data_30 : _GEN_2599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2601 = 8'h1f == _match_key_qbytes_2_T ? phv_data_31 : _GEN_2600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2602 = 8'h20 == _match_key_qbytes_2_T ? phv_data_32 : _GEN_2601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2603 = 8'h21 == _match_key_qbytes_2_T ? phv_data_33 : _GEN_2602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2604 = 8'h22 == _match_key_qbytes_2_T ? phv_data_34 : _GEN_2603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2605 = 8'h23 == _match_key_qbytes_2_T ? phv_data_35 : _GEN_2604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2606 = 8'h24 == _match_key_qbytes_2_T ? phv_data_36 : _GEN_2605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2607 = 8'h25 == _match_key_qbytes_2_T ? phv_data_37 : _GEN_2606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2608 = 8'h26 == _match_key_qbytes_2_T ? phv_data_38 : _GEN_2607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2609 = 8'h27 == _match_key_qbytes_2_T ? phv_data_39 : _GEN_2608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2610 = 8'h28 == _match_key_qbytes_2_T ? phv_data_40 : _GEN_2609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2611 = 8'h29 == _match_key_qbytes_2_T ? phv_data_41 : _GEN_2610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2612 = 8'h2a == _match_key_qbytes_2_T ? phv_data_42 : _GEN_2611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2613 = 8'h2b == _match_key_qbytes_2_T ? phv_data_43 : _GEN_2612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2614 = 8'h2c == _match_key_qbytes_2_T ? phv_data_44 : _GEN_2613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2615 = 8'h2d == _match_key_qbytes_2_T ? phv_data_45 : _GEN_2614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2616 = 8'h2e == _match_key_qbytes_2_T ? phv_data_46 : _GEN_2615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2617 = 8'h2f == _match_key_qbytes_2_T ? phv_data_47 : _GEN_2616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2618 = 8'h30 == _match_key_qbytes_2_T ? phv_data_48 : _GEN_2617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2619 = 8'h31 == _match_key_qbytes_2_T ? phv_data_49 : _GEN_2618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2620 = 8'h32 == _match_key_qbytes_2_T ? phv_data_50 : _GEN_2619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2621 = 8'h33 == _match_key_qbytes_2_T ? phv_data_51 : _GEN_2620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2622 = 8'h34 == _match_key_qbytes_2_T ? phv_data_52 : _GEN_2621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2623 = 8'h35 == _match_key_qbytes_2_T ? phv_data_53 : _GEN_2622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2624 = 8'h36 == _match_key_qbytes_2_T ? phv_data_54 : _GEN_2623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2625 = 8'h37 == _match_key_qbytes_2_T ? phv_data_55 : _GEN_2624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2626 = 8'h38 == _match_key_qbytes_2_T ? phv_data_56 : _GEN_2625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2627 = 8'h39 == _match_key_qbytes_2_T ? phv_data_57 : _GEN_2626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2628 = 8'h3a == _match_key_qbytes_2_T ? phv_data_58 : _GEN_2627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2629 = 8'h3b == _match_key_qbytes_2_T ? phv_data_59 : _GEN_2628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2630 = 8'h3c == _match_key_qbytes_2_T ? phv_data_60 : _GEN_2629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2631 = 8'h3d == _match_key_qbytes_2_T ? phv_data_61 : _GEN_2630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2632 = 8'h3e == _match_key_qbytes_2_T ? phv_data_62 : _GEN_2631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2633 = 8'h3f == _match_key_qbytes_2_T ? phv_data_63 : _GEN_2632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2634 = 8'h40 == _match_key_qbytes_2_T ? phv_data_64 : _GEN_2633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2635 = 8'h41 == _match_key_qbytes_2_T ? phv_data_65 : _GEN_2634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2636 = 8'h42 == _match_key_qbytes_2_T ? phv_data_66 : _GEN_2635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2637 = 8'h43 == _match_key_qbytes_2_T ? phv_data_67 : _GEN_2636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2638 = 8'h44 == _match_key_qbytes_2_T ? phv_data_68 : _GEN_2637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2639 = 8'h45 == _match_key_qbytes_2_T ? phv_data_69 : _GEN_2638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2640 = 8'h46 == _match_key_qbytes_2_T ? phv_data_70 : _GEN_2639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2641 = 8'h47 == _match_key_qbytes_2_T ? phv_data_71 : _GEN_2640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2642 = 8'h48 == _match_key_qbytes_2_T ? phv_data_72 : _GEN_2641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2643 = 8'h49 == _match_key_qbytes_2_T ? phv_data_73 : _GEN_2642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2644 = 8'h4a == _match_key_qbytes_2_T ? phv_data_74 : _GEN_2643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2645 = 8'h4b == _match_key_qbytes_2_T ? phv_data_75 : _GEN_2644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2646 = 8'h4c == _match_key_qbytes_2_T ? phv_data_76 : _GEN_2645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2647 = 8'h4d == _match_key_qbytes_2_T ? phv_data_77 : _GEN_2646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2648 = 8'h4e == _match_key_qbytes_2_T ? phv_data_78 : _GEN_2647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2649 = 8'h4f == _match_key_qbytes_2_T ? phv_data_79 : _GEN_2648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2650 = 8'h50 == _match_key_qbytes_2_T ? phv_data_80 : _GEN_2649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2651 = 8'h51 == _match_key_qbytes_2_T ? phv_data_81 : _GEN_2650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2652 = 8'h52 == _match_key_qbytes_2_T ? phv_data_82 : _GEN_2651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2653 = 8'h53 == _match_key_qbytes_2_T ? phv_data_83 : _GEN_2652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2654 = 8'h54 == _match_key_qbytes_2_T ? phv_data_84 : _GEN_2653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2655 = 8'h55 == _match_key_qbytes_2_T ? phv_data_85 : _GEN_2654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2656 = 8'h56 == _match_key_qbytes_2_T ? phv_data_86 : _GEN_2655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2657 = 8'h57 == _match_key_qbytes_2_T ? phv_data_87 : _GEN_2656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2658 = 8'h58 == _match_key_qbytes_2_T ? phv_data_88 : _GEN_2657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2659 = 8'h59 == _match_key_qbytes_2_T ? phv_data_89 : _GEN_2658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2660 = 8'h5a == _match_key_qbytes_2_T ? phv_data_90 : _GEN_2659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2661 = 8'h5b == _match_key_qbytes_2_T ? phv_data_91 : _GEN_2660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2662 = 8'h5c == _match_key_qbytes_2_T ? phv_data_92 : _GEN_2661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2663 = 8'h5d == _match_key_qbytes_2_T ? phv_data_93 : _GEN_2662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2664 = 8'h5e == _match_key_qbytes_2_T ? phv_data_94 : _GEN_2663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2665 = 8'h5f == _match_key_qbytes_2_T ? phv_data_95 : _GEN_2664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2666 = 8'h60 == _match_key_qbytes_2_T ? phv_data_96 : _GEN_2665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2667 = 8'h61 == _match_key_qbytes_2_T ? phv_data_97 : _GEN_2666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2668 = 8'h62 == _match_key_qbytes_2_T ? phv_data_98 : _GEN_2667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2669 = 8'h63 == _match_key_qbytes_2_T ? phv_data_99 : _GEN_2668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2670 = 8'h64 == _match_key_qbytes_2_T ? phv_data_100 : _GEN_2669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2671 = 8'h65 == _match_key_qbytes_2_T ? phv_data_101 : _GEN_2670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2672 = 8'h66 == _match_key_qbytes_2_T ? phv_data_102 : _GEN_2671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2673 = 8'h67 == _match_key_qbytes_2_T ? phv_data_103 : _GEN_2672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2674 = 8'h68 == _match_key_qbytes_2_T ? phv_data_104 : _GEN_2673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2675 = 8'h69 == _match_key_qbytes_2_T ? phv_data_105 : _GEN_2674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2676 = 8'h6a == _match_key_qbytes_2_T ? phv_data_106 : _GEN_2675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2677 = 8'h6b == _match_key_qbytes_2_T ? phv_data_107 : _GEN_2676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2678 = 8'h6c == _match_key_qbytes_2_T ? phv_data_108 : _GEN_2677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2679 = 8'h6d == _match_key_qbytes_2_T ? phv_data_109 : _GEN_2678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2680 = 8'h6e == _match_key_qbytes_2_T ? phv_data_110 : _GEN_2679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2681 = 8'h6f == _match_key_qbytes_2_T ? phv_data_111 : _GEN_2680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2682 = 8'h70 == _match_key_qbytes_2_T ? phv_data_112 : _GEN_2681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2683 = 8'h71 == _match_key_qbytes_2_T ? phv_data_113 : _GEN_2682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2684 = 8'h72 == _match_key_qbytes_2_T ? phv_data_114 : _GEN_2683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2685 = 8'h73 == _match_key_qbytes_2_T ? phv_data_115 : _GEN_2684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2686 = 8'h74 == _match_key_qbytes_2_T ? phv_data_116 : _GEN_2685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2687 = 8'h75 == _match_key_qbytes_2_T ? phv_data_117 : _GEN_2686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2688 = 8'h76 == _match_key_qbytes_2_T ? phv_data_118 : _GEN_2687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2689 = 8'h77 == _match_key_qbytes_2_T ? phv_data_119 : _GEN_2688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2690 = 8'h78 == _match_key_qbytes_2_T ? phv_data_120 : _GEN_2689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2691 = 8'h79 == _match_key_qbytes_2_T ? phv_data_121 : _GEN_2690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2692 = 8'h7a == _match_key_qbytes_2_T ? phv_data_122 : _GEN_2691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2693 = 8'h7b == _match_key_qbytes_2_T ? phv_data_123 : _GEN_2692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2694 = 8'h7c == _match_key_qbytes_2_T ? phv_data_124 : _GEN_2693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2695 = 8'h7d == _match_key_qbytes_2_T ? phv_data_125 : _GEN_2694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2696 = 8'h7e == _match_key_qbytes_2_T ? phv_data_126 : _GEN_2695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2697 = 8'h7f == _match_key_qbytes_2_T ? phv_data_127 : _GEN_2696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2698 = 8'h80 == _match_key_qbytes_2_T ? phv_data_128 : _GEN_2697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2699 = 8'h81 == _match_key_qbytes_2_T ? phv_data_129 : _GEN_2698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2700 = 8'h82 == _match_key_qbytes_2_T ? phv_data_130 : _GEN_2699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2701 = 8'h83 == _match_key_qbytes_2_T ? phv_data_131 : _GEN_2700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2702 = 8'h84 == _match_key_qbytes_2_T ? phv_data_132 : _GEN_2701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2703 = 8'h85 == _match_key_qbytes_2_T ? phv_data_133 : _GEN_2702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2704 = 8'h86 == _match_key_qbytes_2_T ? phv_data_134 : _GEN_2703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2705 = 8'h87 == _match_key_qbytes_2_T ? phv_data_135 : _GEN_2704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2706 = 8'h88 == _match_key_qbytes_2_T ? phv_data_136 : _GEN_2705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2707 = 8'h89 == _match_key_qbytes_2_T ? phv_data_137 : _GEN_2706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2708 = 8'h8a == _match_key_qbytes_2_T ? phv_data_138 : _GEN_2707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2709 = 8'h8b == _match_key_qbytes_2_T ? phv_data_139 : _GEN_2708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2710 = 8'h8c == _match_key_qbytes_2_T ? phv_data_140 : _GEN_2709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2711 = 8'h8d == _match_key_qbytes_2_T ? phv_data_141 : _GEN_2710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2712 = 8'h8e == _match_key_qbytes_2_T ? phv_data_142 : _GEN_2711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2713 = 8'h8f == _match_key_qbytes_2_T ? phv_data_143 : _GEN_2712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2714 = 8'h90 == _match_key_qbytes_2_T ? phv_data_144 : _GEN_2713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2715 = 8'h91 == _match_key_qbytes_2_T ? phv_data_145 : _GEN_2714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2716 = 8'h92 == _match_key_qbytes_2_T ? phv_data_146 : _GEN_2715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2717 = 8'h93 == _match_key_qbytes_2_T ? phv_data_147 : _GEN_2716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2718 = 8'h94 == _match_key_qbytes_2_T ? phv_data_148 : _GEN_2717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2719 = 8'h95 == _match_key_qbytes_2_T ? phv_data_149 : _GEN_2718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2720 = 8'h96 == _match_key_qbytes_2_T ? phv_data_150 : _GEN_2719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2721 = 8'h97 == _match_key_qbytes_2_T ? phv_data_151 : _GEN_2720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2722 = 8'h98 == _match_key_qbytes_2_T ? phv_data_152 : _GEN_2721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2723 = 8'h99 == _match_key_qbytes_2_T ? phv_data_153 : _GEN_2722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2724 = 8'h9a == _match_key_qbytes_2_T ? phv_data_154 : _GEN_2723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2725 = 8'h9b == _match_key_qbytes_2_T ? phv_data_155 : _GEN_2724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2726 = 8'h9c == _match_key_qbytes_2_T ? phv_data_156 : _GEN_2725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2727 = 8'h9d == _match_key_qbytes_2_T ? phv_data_157 : _GEN_2726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2728 = 8'h9e == _match_key_qbytes_2_T ? phv_data_158 : _GEN_2727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2729 = 8'h9f == _match_key_qbytes_2_T ? phv_data_159 : _GEN_2728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2730 = 8'ha0 == _match_key_qbytes_2_T ? phv_data_160 : _GEN_2729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2731 = 8'ha1 == _match_key_qbytes_2_T ? phv_data_161 : _GEN_2730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2732 = 8'ha2 == _match_key_qbytes_2_T ? phv_data_162 : _GEN_2731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2733 = 8'ha3 == _match_key_qbytes_2_T ? phv_data_163 : _GEN_2732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2734 = 8'ha4 == _match_key_qbytes_2_T ? phv_data_164 : _GEN_2733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2735 = 8'ha5 == _match_key_qbytes_2_T ? phv_data_165 : _GEN_2734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2736 = 8'ha6 == _match_key_qbytes_2_T ? phv_data_166 : _GEN_2735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2737 = 8'ha7 == _match_key_qbytes_2_T ? phv_data_167 : _GEN_2736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2738 = 8'ha8 == _match_key_qbytes_2_T ? phv_data_168 : _GEN_2737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2739 = 8'ha9 == _match_key_qbytes_2_T ? phv_data_169 : _GEN_2738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2740 = 8'haa == _match_key_qbytes_2_T ? phv_data_170 : _GEN_2739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2741 = 8'hab == _match_key_qbytes_2_T ? phv_data_171 : _GEN_2740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2742 = 8'hac == _match_key_qbytes_2_T ? phv_data_172 : _GEN_2741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2743 = 8'had == _match_key_qbytes_2_T ? phv_data_173 : _GEN_2742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2744 = 8'hae == _match_key_qbytes_2_T ? phv_data_174 : _GEN_2743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2745 = 8'haf == _match_key_qbytes_2_T ? phv_data_175 : _GEN_2744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2746 = 8'hb0 == _match_key_qbytes_2_T ? phv_data_176 : _GEN_2745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2747 = 8'hb1 == _match_key_qbytes_2_T ? phv_data_177 : _GEN_2746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2748 = 8'hb2 == _match_key_qbytes_2_T ? phv_data_178 : _GEN_2747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2749 = 8'hb3 == _match_key_qbytes_2_T ? phv_data_179 : _GEN_2748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2750 = 8'hb4 == _match_key_qbytes_2_T ? phv_data_180 : _GEN_2749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2751 = 8'hb5 == _match_key_qbytes_2_T ? phv_data_181 : _GEN_2750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2752 = 8'hb6 == _match_key_qbytes_2_T ? phv_data_182 : _GEN_2751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2753 = 8'hb7 == _match_key_qbytes_2_T ? phv_data_183 : _GEN_2752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2754 = 8'hb8 == _match_key_qbytes_2_T ? phv_data_184 : _GEN_2753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2755 = 8'hb9 == _match_key_qbytes_2_T ? phv_data_185 : _GEN_2754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2756 = 8'hba == _match_key_qbytes_2_T ? phv_data_186 : _GEN_2755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2757 = 8'hbb == _match_key_qbytes_2_T ? phv_data_187 : _GEN_2756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2758 = 8'hbc == _match_key_qbytes_2_T ? phv_data_188 : _GEN_2757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2759 = 8'hbd == _match_key_qbytes_2_T ? phv_data_189 : _GEN_2758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2760 = 8'hbe == _match_key_qbytes_2_T ? phv_data_190 : _GEN_2759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2761 = 8'hbf == _match_key_qbytes_2_T ? phv_data_191 : _GEN_2760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2762 = 8'hc0 == _match_key_qbytes_2_T ? phv_data_192 : _GEN_2761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2763 = 8'hc1 == _match_key_qbytes_2_T ? phv_data_193 : _GEN_2762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2764 = 8'hc2 == _match_key_qbytes_2_T ? phv_data_194 : _GEN_2763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2765 = 8'hc3 == _match_key_qbytes_2_T ? phv_data_195 : _GEN_2764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2766 = 8'hc4 == _match_key_qbytes_2_T ? phv_data_196 : _GEN_2765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2767 = 8'hc5 == _match_key_qbytes_2_T ? phv_data_197 : _GEN_2766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2768 = 8'hc6 == _match_key_qbytes_2_T ? phv_data_198 : _GEN_2767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2769 = 8'hc7 == _match_key_qbytes_2_T ? phv_data_199 : _GEN_2768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2770 = 8'hc8 == _match_key_qbytes_2_T ? phv_data_200 : _GEN_2769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2771 = 8'hc9 == _match_key_qbytes_2_T ? phv_data_201 : _GEN_2770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2772 = 8'hca == _match_key_qbytes_2_T ? phv_data_202 : _GEN_2771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2773 = 8'hcb == _match_key_qbytes_2_T ? phv_data_203 : _GEN_2772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2774 = 8'hcc == _match_key_qbytes_2_T ? phv_data_204 : _GEN_2773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2775 = 8'hcd == _match_key_qbytes_2_T ? phv_data_205 : _GEN_2774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2776 = 8'hce == _match_key_qbytes_2_T ? phv_data_206 : _GEN_2775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2777 = 8'hcf == _match_key_qbytes_2_T ? phv_data_207 : _GEN_2776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2778 = 8'hd0 == _match_key_qbytes_2_T ? phv_data_208 : _GEN_2777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2779 = 8'hd1 == _match_key_qbytes_2_T ? phv_data_209 : _GEN_2778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2780 = 8'hd2 == _match_key_qbytes_2_T ? phv_data_210 : _GEN_2779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2781 = 8'hd3 == _match_key_qbytes_2_T ? phv_data_211 : _GEN_2780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2782 = 8'hd4 == _match_key_qbytes_2_T ? phv_data_212 : _GEN_2781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2783 = 8'hd5 == _match_key_qbytes_2_T ? phv_data_213 : _GEN_2782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2784 = 8'hd6 == _match_key_qbytes_2_T ? phv_data_214 : _GEN_2783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2785 = 8'hd7 == _match_key_qbytes_2_T ? phv_data_215 : _GEN_2784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2786 = 8'hd8 == _match_key_qbytes_2_T ? phv_data_216 : _GEN_2785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2787 = 8'hd9 == _match_key_qbytes_2_T ? phv_data_217 : _GEN_2786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2788 = 8'hda == _match_key_qbytes_2_T ? phv_data_218 : _GEN_2787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2789 = 8'hdb == _match_key_qbytes_2_T ? phv_data_219 : _GEN_2788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2790 = 8'hdc == _match_key_qbytes_2_T ? phv_data_220 : _GEN_2789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2791 = 8'hdd == _match_key_qbytes_2_T ? phv_data_221 : _GEN_2790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2792 = 8'hde == _match_key_qbytes_2_T ? phv_data_222 : _GEN_2791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2793 = 8'hdf == _match_key_qbytes_2_T ? phv_data_223 : _GEN_2792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2794 = 8'he0 == _match_key_qbytes_2_T ? phv_data_224 : _GEN_2793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2795 = 8'he1 == _match_key_qbytes_2_T ? phv_data_225 : _GEN_2794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2796 = 8'he2 == _match_key_qbytes_2_T ? phv_data_226 : _GEN_2795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2797 = 8'he3 == _match_key_qbytes_2_T ? phv_data_227 : _GEN_2796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2798 = 8'he4 == _match_key_qbytes_2_T ? phv_data_228 : _GEN_2797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2799 = 8'he5 == _match_key_qbytes_2_T ? phv_data_229 : _GEN_2798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2800 = 8'he6 == _match_key_qbytes_2_T ? phv_data_230 : _GEN_2799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2801 = 8'he7 == _match_key_qbytes_2_T ? phv_data_231 : _GEN_2800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2802 = 8'he8 == _match_key_qbytes_2_T ? phv_data_232 : _GEN_2801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2803 = 8'he9 == _match_key_qbytes_2_T ? phv_data_233 : _GEN_2802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2804 = 8'hea == _match_key_qbytes_2_T ? phv_data_234 : _GEN_2803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2805 = 8'heb == _match_key_qbytes_2_T ? phv_data_235 : _GEN_2804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2806 = 8'hec == _match_key_qbytes_2_T ? phv_data_236 : _GEN_2805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2807 = 8'hed == _match_key_qbytes_2_T ? phv_data_237 : _GEN_2806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2808 = 8'hee == _match_key_qbytes_2_T ? phv_data_238 : _GEN_2807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2809 = 8'hef == _match_key_qbytes_2_T ? phv_data_239 : _GEN_2808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2810 = 8'hf0 == _match_key_qbytes_2_T ? phv_data_240 : _GEN_2809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2811 = 8'hf1 == _match_key_qbytes_2_T ? phv_data_241 : _GEN_2810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2812 = 8'hf2 == _match_key_qbytes_2_T ? phv_data_242 : _GEN_2811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2813 = 8'hf3 == _match_key_qbytes_2_T ? phv_data_243 : _GEN_2812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2814 = 8'hf4 == _match_key_qbytes_2_T ? phv_data_244 : _GEN_2813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2815 = 8'hf5 == _match_key_qbytes_2_T ? phv_data_245 : _GEN_2814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2816 = 8'hf6 == _match_key_qbytes_2_T ? phv_data_246 : _GEN_2815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2817 = 8'hf7 == _match_key_qbytes_2_T ? phv_data_247 : _GEN_2816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2818 = 8'hf8 == _match_key_qbytes_2_T ? phv_data_248 : _GEN_2817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2819 = 8'hf9 == _match_key_qbytes_2_T ? phv_data_249 : _GEN_2818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2820 = 8'hfa == _match_key_qbytes_2_T ? phv_data_250 : _GEN_2819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2821 = 8'hfb == _match_key_qbytes_2_T ? phv_data_251 : _GEN_2820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2822 = 8'hfc == _match_key_qbytes_2_T ? phv_data_252 : _GEN_2821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2823 = 8'hfd == _match_key_qbytes_2_T ? phv_data_253 : _GEN_2822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2824 = 8'hfe == _match_key_qbytes_2_T ? phv_data_254 : _GEN_2823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2825 = 8'hff == _match_key_qbytes_2_T ? phv_data_255 : _GEN_2824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2827 = 8'h1 == _match_key_qbytes_2_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2828 = 8'h2 == _match_key_qbytes_2_T_1 ? phv_data_2 : _GEN_2827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2829 = 8'h3 == _match_key_qbytes_2_T_1 ? phv_data_3 : _GEN_2828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2830 = 8'h4 == _match_key_qbytes_2_T_1 ? phv_data_4 : _GEN_2829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2831 = 8'h5 == _match_key_qbytes_2_T_1 ? phv_data_5 : _GEN_2830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2832 = 8'h6 == _match_key_qbytes_2_T_1 ? phv_data_6 : _GEN_2831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2833 = 8'h7 == _match_key_qbytes_2_T_1 ? phv_data_7 : _GEN_2832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2834 = 8'h8 == _match_key_qbytes_2_T_1 ? phv_data_8 : _GEN_2833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2835 = 8'h9 == _match_key_qbytes_2_T_1 ? phv_data_9 : _GEN_2834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2836 = 8'ha == _match_key_qbytes_2_T_1 ? phv_data_10 : _GEN_2835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2837 = 8'hb == _match_key_qbytes_2_T_1 ? phv_data_11 : _GEN_2836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2838 = 8'hc == _match_key_qbytes_2_T_1 ? phv_data_12 : _GEN_2837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2839 = 8'hd == _match_key_qbytes_2_T_1 ? phv_data_13 : _GEN_2838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2840 = 8'he == _match_key_qbytes_2_T_1 ? phv_data_14 : _GEN_2839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2841 = 8'hf == _match_key_qbytes_2_T_1 ? phv_data_15 : _GEN_2840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2842 = 8'h10 == _match_key_qbytes_2_T_1 ? phv_data_16 : _GEN_2841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2843 = 8'h11 == _match_key_qbytes_2_T_1 ? phv_data_17 : _GEN_2842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2844 = 8'h12 == _match_key_qbytes_2_T_1 ? phv_data_18 : _GEN_2843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2845 = 8'h13 == _match_key_qbytes_2_T_1 ? phv_data_19 : _GEN_2844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2846 = 8'h14 == _match_key_qbytes_2_T_1 ? phv_data_20 : _GEN_2845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2847 = 8'h15 == _match_key_qbytes_2_T_1 ? phv_data_21 : _GEN_2846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2848 = 8'h16 == _match_key_qbytes_2_T_1 ? phv_data_22 : _GEN_2847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2849 = 8'h17 == _match_key_qbytes_2_T_1 ? phv_data_23 : _GEN_2848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2850 = 8'h18 == _match_key_qbytes_2_T_1 ? phv_data_24 : _GEN_2849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2851 = 8'h19 == _match_key_qbytes_2_T_1 ? phv_data_25 : _GEN_2850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2852 = 8'h1a == _match_key_qbytes_2_T_1 ? phv_data_26 : _GEN_2851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2853 = 8'h1b == _match_key_qbytes_2_T_1 ? phv_data_27 : _GEN_2852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2854 = 8'h1c == _match_key_qbytes_2_T_1 ? phv_data_28 : _GEN_2853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2855 = 8'h1d == _match_key_qbytes_2_T_1 ? phv_data_29 : _GEN_2854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2856 = 8'h1e == _match_key_qbytes_2_T_1 ? phv_data_30 : _GEN_2855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2857 = 8'h1f == _match_key_qbytes_2_T_1 ? phv_data_31 : _GEN_2856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2858 = 8'h20 == _match_key_qbytes_2_T_1 ? phv_data_32 : _GEN_2857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2859 = 8'h21 == _match_key_qbytes_2_T_1 ? phv_data_33 : _GEN_2858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2860 = 8'h22 == _match_key_qbytes_2_T_1 ? phv_data_34 : _GEN_2859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2861 = 8'h23 == _match_key_qbytes_2_T_1 ? phv_data_35 : _GEN_2860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2862 = 8'h24 == _match_key_qbytes_2_T_1 ? phv_data_36 : _GEN_2861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2863 = 8'h25 == _match_key_qbytes_2_T_1 ? phv_data_37 : _GEN_2862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2864 = 8'h26 == _match_key_qbytes_2_T_1 ? phv_data_38 : _GEN_2863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2865 = 8'h27 == _match_key_qbytes_2_T_1 ? phv_data_39 : _GEN_2864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2866 = 8'h28 == _match_key_qbytes_2_T_1 ? phv_data_40 : _GEN_2865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2867 = 8'h29 == _match_key_qbytes_2_T_1 ? phv_data_41 : _GEN_2866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2868 = 8'h2a == _match_key_qbytes_2_T_1 ? phv_data_42 : _GEN_2867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2869 = 8'h2b == _match_key_qbytes_2_T_1 ? phv_data_43 : _GEN_2868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2870 = 8'h2c == _match_key_qbytes_2_T_1 ? phv_data_44 : _GEN_2869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2871 = 8'h2d == _match_key_qbytes_2_T_1 ? phv_data_45 : _GEN_2870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2872 = 8'h2e == _match_key_qbytes_2_T_1 ? phv_data_46 : _GEN_2871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2873 = 8'h2f == _match_key_qbytes_2_T_1 ? phv_data_47 : _GEN_2872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2874 = 8'h30 == _match_key_qbytes_2_T_1 ? phv_data_48 : _GEN_2873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2875 = 8'h31 == _match_key_qbytes_2_T_1 ? phv_data_49 : _GEN_2874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2876 = 8'h32 == _match_key_qbytes_2_T_1 ? phv_data_50 : _GEN_2875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2877 = 8'h33 == _match_key_qbytes_2_T_1 ? phv_data_51 : _GEN_2876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2878 = 8'h34 == _match_key_qbytes_2_T_1 ? phv_data_52 : _GEN_2877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2879 = 8'h35 == _match_key_qbytes_2_T_1 ? phv_data_53 : _GEN_2878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2880 = 8'h36 == _match_key_qbytes_2_T_1 ? phv_data_54 : _GEN_2879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2881 = 8'h37 == _match_key_qbytes_2_T_1 ? phv_data_55 : _GEN_2880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2882 = 8'h38 == _match_key_qbytes_2_T_1 ? phv_data_56 : _GEN_2881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2883 = 8'h39 == _match_key_qbytes_2_T_1 ? phv_data_57 : _GEN_2882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2884 = 8'h3a == _match_key_qbytes_2_T_1 ? phv_data_58 : _GEN_2883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2885 = 8'h3b == _match_key_qbytes_2_T_1 ? phv_data_59 : _GEN_2884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2886 = 8'h3c == _match_key_qbytes_2_T_1 ? phv_data_60 : _GEN_2885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2887 = 8'h3d == _match_key_qbytes_2_T_1 ? phv_data_61 : _GEN_2886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2888 = 8'h3e == _match_key_qbytes_2_T_1 ? phv_data_62 : _GEN_2887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2889 = 8'h3f == _match_key_qbytes_2_T_1 ? phv_data_63 : _GEN_2888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2890 = 8'h40 == _match_key_qbytes_2_T_1 ? phv_data_64 : _GEN_2889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2891 = 8'h41 == _match_key_qbytes_2_T_1 ? phv_data_65 : _GEN_2890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2892 = 8'h42 == _match_key_qbytes_2_T_1 ? phv_data_66 : _GEN_2891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2893 = 8'h43 == _match_key_qbytes_2_T_1 ? phv_data_67 : _GEN_2892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2894 = 8'h44 == _match_key_qbytes_2_T_1 ? phv_data_68 : _GEN_2893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2895 = 8'h45 == _match_key_qbytes_2_T_1 ? phv_data_69 : _GEN_2894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2896 = 8'h46 == _match_key_qbytes_2_T_1 ? phv_data_70 : _GEN_2895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2897 = 8'h47 == _match_key_qbytes_2_T_1 ? phv_data_71 : _GEN_2896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2898 = 8'h48 == _match_key_qbytes_2_T_1 ? phv_data_72 : _GEN_2897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2899 = 8'h49 == _match_key_qbytes_2_T_1 ? phv_data_73 : _GEN_2898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2900 = 8'h4a == _match_key_qbytes_2_T_1 ? phv_data_74 : _GEN_2899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2901 = 8'h4b == _match_key_qbytes_2_T_1 ? phv_data_75 : _GEN_2900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2902 = 8'h4c == _match_key_qbytes_2_T_1 ? phv_data_76 : _GEN_2901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2903 = 8'h4d == _match_key_qbytes_2_T_1 ? phv_data_77 : _GEN_2902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2904 = 8'h4e == _match_key_qbytes_2_T_1 ? phv_data_78 : _GEN_2903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2905 = 8'h4f == _match_key_qbytes_2_T_1 ? phv_data_79 : _GEN_2904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2906 = 8'h50 == _match_key_qbytes_2_T_1 ? phv_data_80 : _GEN_2905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2907 = 8'h51 == _match_key_qbytes_2_T_1 ? phv_data_81 : _GEN_2906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2908 = 8'h52 == _match_key_qbytes_2_T_1 ? phv_data_82 : _GEN_2907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2909 = 8'h53 == _match_key_qbytes_2_T_1 ? phv_data_83 : _GEN_2908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2910 = 8'h54 == _match_key_qbytes_2_T_1 ? phv_data_84 : _GEN_2909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2911 = 8'h55 == _match_key_qbytes_2_T_1 ? phv_data_85 : _GEN_2910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2912 = 8'h56 == _match_key_qbytes_2_T_1 ? phv_data_86 : _GEN_2911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2913 = 8'h57 == _match_key_qbytes_2_T_1 ? phv_data_87 : _GEN_2912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2914 = 8'h58 == _match_key_qbytes_2_T_1 ? phv_data_88 : _GEN_2913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2915 = 8'h59 == _match_key_qbytes_2_T_1 ? phv_data_89 : _GEN_2914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2916 = 8'h5a == _match_key_qbytes_2_T_1 ? phv_data_90 : _GEN_2915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2917 = 8'h5b == _match_key_qbytes_2_T_1 ? phv_data_91 : _GEN_2916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2918 = 8'h5c == _match_key_qbytes_2_T_1 ? phv_data_92 : _GEN_2917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2919 = 8'h5d == _match_key_qbytes_2_T_1 ? phv_data_93 : _GEN_2918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2920 = 8'h5e == _match_key_qbytes_2_T_1 ? phv_data_94 : _GEN_2919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2921 = 8'h5f == _match_key_qbytes_2_T_1 ? phv_data_95 : _GEN_2920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2922 = 8'h60 == _match_key_qbytes_2_T_1 ? phv_data_96 : _GEN_2921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2923 = 8'h61 == _match_key_qbytes_2_T_1 ? phv_data_97 : _GEN_2922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2924 = 8'h62 == _match_key_qbytes_2_T_1 ? phv_data_98 : _GEN_2923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2925 = 8'h63 == _match_key_qbytes_2_T_1 ? phv_data_99 : _GEN_2924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2926 = 8'h64 == _match_key_qbytes_2_T_1 ? phv_data_100 : _GEN_2925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2927 = 8'h65 == _match_key_qbytes_2_T_1 ? phv_data_101 : _GEN_2926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2928 = 8'h66 == _match_key_qbytes_2_T_1 ? phv_data_102 : _GEN_2927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2929 = 8'h67 == _match_key_qbytes_2_T_1 ? phv_data_103 : _GEN_2928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2930 = 8'h68 == _match_key_qbytes_2_T_1 ? phv_data_104 : _GEN_2929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2931 = 8'h69 == _match_key_qbytes_2_T_1 ? phv_data_105 : _GEN_2930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2932 = 8'h6a == _match_key_qbytes_2_T_1 ? phv_data_106 : _GEN_2931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2933 = 8'h6b == _match_key_qbytes_2_T_1 ? phv_data_107 : _GEN_2932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2934 = 8'h6c == _match_key_qbytes_2_T_1 ? phv_data_108 : _GEN_2933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2935 = 8'h6d == _match_key_qbytes_2_T_1 ? phv_data_109 : _GEN_2934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2936 = 8'h6e == _match_key_qbytes_2_T_1 ? phv_data_110 : _GEN_2935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2937 = 8'h6f == _match_key_qbytes_2_T_1 ? phv_data_111 : _GEN_2936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2938 = 8'h70 == _match_key_qbytes_2_T_1 ? phv_data_112 : _GEN_2937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2939 = 8'h71 == _match_key_qbytes_2_T_1 ? phv_data_113 : _GEN_2938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2940 = 8'h72 == _match_key_qbytes_2_T_1 ? phv_data_114 : _GEN_2939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2941 = 8'h73 == _match_key_qbytes_2_T_1 ? phv_data_115 : _GEN_2940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2942 = 8'h74 == _match_key_qbytes_2_T_1 ? phv_data_116 : _GEN_2941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2943 = 8'h75 == _match_key_qbytes_2_T_1 ? phv_data_117 : _GEN_2942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2944 = 8'h76 == _match_key_qbytes_2_T_1 ? phv_data_118 : _GEN_2943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2945 = 8'h77 == _match_key_qbytes_2_T_1 ? phv_data_119 : _GEN_2944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2946 = 8'h78 == _match_key_qbytes_2_T_1 ? phv_data_120 : _GEN_2945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2947 = 8'h79 == _match_key_qbytes_2_T_1 ? phv_data_121 : _GEN_2946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2948 = 8'h7a == _match_key_qbytes_2_T_1 ? phv_data_122 : _GEN_2947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2949 = 8'h7b == _match_key_qbytes_2_T_1 ? phv_data_123 : _GEN_2948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2950 = 8'h7c == _match_key_qbytes_2_T_1 ? phv_data_124 : _GEN_2949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2951 = 8'h7d == _match_key_qbytes_2_T_1 ? phv_data_125 : _GEN_2950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2952 = 8'h7e == _match_key_qbytes_2_T_1 ? phv_data_126 : _GEN_2951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2953 = 8'h7f == _match_key_qbytes_2_T_1 ? phv_data_127 : _GEN_2952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2954 = 8'h80 == _match_key_qbytes_2_T_1 ? phv_data_128 : _GEN_2953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2955 = 8'h81 == _match_key_qbytes_2_T_1 ? phv_data_129 : _GEN_2954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2956 = 8'h82 == _match_key_qbytes_2_T_1 ? phv_data_130 : _GEN_2955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2957 = 8'h83 == _match_key_qbytes_2_T_1 ? phv_data_131 : _GEN_2956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2958 = 8'h84 == _match_key_qbytes_2_T_1 ? phv_data_132 : _GEN_2957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2959 = 8'h85 == _match_key_qbytes_2_T_1 ? phv_data_133 : _GEN_2958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2960 = 8'h86 == _match_key_qbytes_2_T_1 ? phv_data_134 : _GEN_2959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2961 = 8'h87 == _match_key_qbytes_2_T_1 ? phv_data_135 : _GEN_2960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2962 = 8'h88 == _match_key_qbytes_2_T_1 ? phv_data_136 : _GEN_2961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2963 = 8'h89 == _match_key_qbytes_2_T_1 ? phv_data_137 : _GEN_2962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2964 = 8'h8a == _match_key_qbytes_2_T_1 ? phv_data_138 : _GEN_2963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2965 = 8'h8b == _match_key_qbytes_2_T_1 ? phv_data_139 : _GEN_2964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2966 = 8'h8c == _match_key_qbytes_2_T_1 ? phv_data_140 : _GEN_2965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2967 = 8'h8d == _match_key_qbytes_2_T_1 ? phv_data_141 : _GEN_2966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2968 = 8'h8e == _match_key_qbytes_2_T_1 ? phv_data_142 : _GEN_2967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2969 = 8'h8f == _match_key_qbytes_2_T_1 ? phv_data_143 : _GEN_2968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2970 = 8'h90 == _match_key_qbytes_2_T_1 ? phv_data_144 : _GEN_2969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2971 = 8'h91 == _match_key_qbytes_2_T_1 ? phv_data_145 : _GEN_2970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2972 = 8'h92 == _match_key_qbytes_2_T_1 ? phv_data_146 : _GEN_2971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2973 = 8'h93 == _match_key_qbytes_2_T_1 ? phv_data_147 : _GEN_2972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2974 = 8'h94 == _match_key_qbytes_2_T_1 ? phv_data_148 : _GEN_2973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2975 = 8'h95 == _match_key_qbytes_2_T_1 ? phv_data_149 : _GEN_2974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2976 = 8'h96 == _match_key_qbytes_2_T_1 ? phv_data_150 : _GEN_2975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2977 = 8'h97 == _match_key_qbytes_2_T_1 ? phv_data_151 : _GEN_2976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2978 = 8'h98 == _match_key_qbytes_2_T_1 ? phv_data_152 : _GEN_2977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2979 = 8'h99 == _match_key_qbytes_2_T_1 ? phv_data_153 : _GEN_2978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2980 = 8'h9a == _match_key_qbytes_2_T_1 ? phv_data_154 : _GEN_2979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2981 = 8'h9b == _match_key_qbytes_2_T_1 ? phv_data_155 : _GEN_2980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2982 = 8'h9c == _match_key_qbytes_2_T_1 ? phv_data_156 : _GEN_2981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2983 = 8'h9d == _match_key_qbytes_2_T_1 ? phv_data_157 : _GEN_2982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2984 = 8'h9e == _match_key_qbytes_2_T_1 ? phv_data_158 : _GEN_2983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2985 = 8'h9f == _match_key_qbytes_2_T_1 ? phv_data_159 : _GEN_2984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2986 = 8'ha0 == _match_key_qbytes_2_T_1 ? phv_data_160 : _GEN_2985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2987 = 8'ha1 == _match_key_qbytes_2_T_1 ? phv_data_161 : _GEN_2986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2988 = 8'ha2 == _match_key_qbytes_2_T_1 ? phv_data_162 : _GEN_2987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2989 = 8'ha3 == _match_key_qbytes_2_T_1 ? phv_data_163 : _GEN_2988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2990 = 8'ha4 == _match_key_qbytes_2_T_1 ? phv_data_164 : _GEN_2989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2991 = 8'ha5 == _match_key_qbytes_2_T_1 ? phv_data_165 : _GEN_2990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2992 = 8'ha6 == _match_key_qbytes_2_T_1 ? phv_data_166 : _GEN_2991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2993 = 8'ha7 == _match_key_qbytes_2_T_1 ? phv_data_167 : _GEN_2992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2994 = 8'ha8 == _match_key_qbytes_2_T_1 ? phv_data_168 : _GEN_2993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2995 = 8'ha9 == _match_key_qbytes_2_T_1 ? phv_data_169 : _GEN_2994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2996 = 8'haa == _match_key_qbytes_2_T_1 ? phv_data_170 : _GEN_2995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2997 = 8'hab == _match_key_qbytes_2_T_1 ? phv_data_171 : _GEN_2996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2998 = 8'hac == _match_key_qbytes_2_T_1 ? phv_data_172 : _GEN_2997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2999 = 8'had == _match_key_qbytes_2_T_1 ? phv_data_173 : _GEN_2998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3000 = 8'hae == _match_key_qbytes_2_T_1 ? phv_data_174 : _GEN_2999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3001 = 8'haf == _match_key_qbytes_2_T_1 ? phv_data_175 : _GEN_3000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3002 = 8'hb0 == _match_key_qbytes_2_T_1 ? phv_data_176 : _GEN_3001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3003 = 8'hb1 == _match_key_qbytes_2_T_1 ? phv_data_177 : _GEN_3002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3004 = 8'hb2 == _match_key_qbytes_2_T_1 ? phv_data_178 : _GEN_3003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3005 = 8'hb3 == _match_key_qbytes_2_T_1 ? phv_data_179 : _GEN_3004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3006 = 8'hb4 == _match_key_qbytes_2_T_1 ? phv_data_180 : _GEN_3005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3007 = 8'hb5 == _match_key_qbytes_2_T_1 ? phv_data_181 : _GEN_3006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3008 = 8'hb6 == _match_key_qbytes_2_T_1 ? phv_data_182 : _GEN_3007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3009 = 8'hb7 == _match_key_qbytes_2_T_1 ? phv_data_183 : _GEN_3008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3010 = 8'hb8 == _match_key_qbytes_2_T_1 ? phv_data_184 : _GEN_3009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3011 = 8'hb9 == _match_key_qbytes_2_T_1 ? phv_data_185 : _GEN_3010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3012 = 8'hba == _match_key_qbytes_2_T_1 ? phv_data_186 : _GEN_3011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3013 = 8'hbb == _match_key_qbytes_2_T_1 ? phv_data_187 : _GEN_3012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3014 = 8'hbc == _match_key_qbytes_2_T_1 ? phv_data_188 : _GEN_3013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3015 = 8'hbd == _match_key_qbytes_2_T_1 ? phv_data_189 : _GEN_3014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3016 = 8'hbe == _match_key_qbytes_2_T_1 ? phv_data_190 : _GEN_3015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3017 = 8'hbf == _match_key_qbytes_2_T_1 ? phv_data_191 : _GEN_3016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3018 = 8'hc0 == _match_key_qbytes_2_T_1 ? phv_data_192 : _GEN_3017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3019 = 8'hc1 == _match_key_qbytes_2_T_1 ? phv_data_193 : _GEN_3018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3020 = 8'hc2 == _match_key_qbytes_2_T_1 ? phv_data_194 : _GEN_3019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3021 = 8'hc3 == _match_key_qbytes_2_T_1 ? phv_data_195 : _GEN_3020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3022 = 8'hc4 == _match_key_qbytes_2_T_1 ? phv_data_196 : _GEN_3021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3023 = 8'hc5 == _match_key_qbytes_2_T_1 ? phv_data_197 : _GEN_3022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3024 = 8'hc6 == _match_key_qbytes_2_T_1 ? phv_data_198 : _GEN_3023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3025 = 8'hc7 == _match_key_qbytes_2_T_1 ? phv_data_199 : _GEN_3024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3026 = 8'hc8 == _match_key_qbytes_2_T_1 ? phv_data_200 : _GEN_3025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3027 = 8'hc9 == _match_key_qbytes_2_T_1 ? phv_data_201 : _GEN_3026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3028 = 8'hca == _match_key_qbytes_2_T_1 ? phv_data_202 : _GEN_3027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3029 = 8'hcb == _match_key_qbytes_2_T_1 ? phv_data_203 : _GEN_3028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3030 = 8'hcc == _match_key_qbytes_2_T_1 ? phv_data_204 : _GEN_3029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3031 = 8'hcd == _match_key_qbytes_2_T_1 ? phv_data_205 : _GEN_3030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3032 = 8'hce == _match_key_qbytes_2_T_1 ? phv_data_206 : _GEN_3031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3033 = 8'hcf == _match_key_qbytes_2_T_1 ? phv_data_207 : _GEN_3032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3034 = 8'hd0 == _match_key_qbytes_2_T_1 ? phv_data_208 : _GEN_3033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3035 = 8'hd1 == _match_key_qbytes_2_T_1 ? phv_data_209 : _GEN_3034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3036 = 8'hd2 == _match_key_qbytes_2_T_1 ? phv_data_210 : _GEN_3035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3037 = 8'hd3 == _match_key_qbytes_2_T_1 ? phv_data_211 : _GEN_3036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3038 = 8'hd4 == _match_key_qbytes_2_T_1 ? phv_data_212 : _GEN_3037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3039 = 8'hd5 == _match_key_qbytes_2_T_1 ? phv_data_213 : _GEN_3038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3040 = 8'hd6 == _match_key_qbytes_2_T_1 ? phv_data_214 : _GEN_3039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3041 = 8'hd7 == _match_key_qbytes_2_T_1 ? phv_data_215 : _GEN_3040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3042 = 8'hd8 == _match_key_qbytes_2_T_1 ? phv_data_216 : _GEN_3041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3043 = 8'hd9 == _match_key_qbytes_2_T_1 ? phv_data_217 : _GEN_3042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3044 = 8'hda == _match_key_qbytes_2_T_1 ? phv_data_218 : _GEN_3043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3045 = 8'hdb == _match_key_qbytes_2_T_1 ? phv_data_219 : _GEN_3044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3046 = 8'hdc == _match_key_qbytes_2_T_1 ? phv_data_220 : _GEN_3045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3047 = 8'hdd == _match_key_qbytes_2_T_1 ? phv_data_221 : _GEN_3046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3048 = 8'hde == _match_key_qbytes_2_T_1 ? phv_data_222 : _GEN_3047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3049 = 8'hdf == _match_key_qbytes_2_T_1 ? phv_data_223 : _GEN_3048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3050 = 8'he0 == _match_key_qbytes_2_T_1 ? phv_data_224 : _GEN_3049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3051 = 8'he1 == _match_key_qbytes_2_T_1 ? phv_data_225 : _GEN_3050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3052 = 8'he2 == _match_key_qbytes_2_T_1 ? phv_data_226 : _GEN_3051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3053 = 8'he3 == _match_key_qbytes_2_T_1 ? phv_data_227 : _GEN_3052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3054 = 8'he4 == _match_key_qbytes_2_T_1 ? phv_data_228 : _GEN_3053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3055 = 8'he5 == _match_key_qbytes_2_T_1 ? phv_data_229 : _GEN_3054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3056 = 8'he6 == _match_key_qbytes_2_T_1 ? phv_data_230 : _GEN_3055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3057 = 8'he7 == _match_key_qbytes_2_T_1 ? phv_data_231 : _GEN_3056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3058 = 8'he8 == _match_key_qbytes_2_T_1 ? phv_data_232 : _GEN_3057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3059 = 8'he9 == _match_key_qbytes_2_T_1 ? phv_data_233 : _GEN_3058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3060 = 8'hea == _match_key_qbytes_2_T_1 ? phv_data_234 : _GEN_3059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3061 = 8'heb == _match_key_qbytes_2_T_1 ? phv_data_235 : _GEN_3060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3062 = 8'hec == _match_key_qbytes_2_T_1 ? phv_data_236 : _GEN_3061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3063 = 8'hed == _match_key_qbytes_2_T_1 ? phv_data_237 : _GEN_3062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3064 = 8'hee == _match_key_qbytes_2_T_1 ? phv_data_238 : _GEN_3063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3065 = 8'hef == _match_key_qbytes_2_T_1 ? phv_data_239 : _GEN_3064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3066 = 8'hf0 == _match_key_qbytes_2_T_1 ? phv_data_240 : _GEN_3065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3067 = 8'hf1 == _match_key_qbytes_2_T_1 ? phv_data_241 : _GEN_3066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3068 = 8'hf2 == _match_key_qbytes_2_T_1 ? phv_data_242 : _GEN_3067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3069 = 8'hf3 == _match_key_qbytes_2_T_1 ? phv_data_243 : _GEN_3068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3070 = 8'hf4 == _match_key_qbytes_2_T_1 ? phv_data_244 : _GEN_3069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3071 = 8'hf5 == _match_key_qbytes_2_T_1 ? phv_data_245 : _GEN_3070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3072 = 8'hf6 == _match_key_qbytes_2_T_1 ? phv_data_246 : _GEN_3071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3073 = 8'hf7 == _match_key_qbytes_2_T_1 ? phv_data_247 : _GEN_3072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3074 = 8'hf8 == _match_key_qbytes_2_T_1 ? phv_data_248 : _GEN_3073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3075 = 8'hf9 == _match_key_qbytes_2_T_1 ? phv_data_249 : _GEN_3074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3076 = 8'hfa == _match_key_qbytes_2_T_1 ? phv_data_250 : _GEN_3075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3077 = 8'hfb == _match_key_qbytes_2_T_1 ? phv_data_251 : _GEN_3076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3078 = 8'hfc == _match_key_qbytes_2_T_1 ? phv_data_252 : _GEN_3077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3079 = 8'hfd == _match_key_qbytes_2_T_1 ? phv_data_253 : _GEN_3078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3080 = 8'hfe == _match_key_qbytes_2_T_1 ? phv_data_254 : _GEN_3079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3081 = 8'hff == _match_key_qbytes_2_T_1 ? phv_data_255 : _GEN_3080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_2_T_3 = {_GEN_2825,_GEN_3081,_GEN_2313,_GEN_2569}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_2 = local_offset_2 < end_offset ? _match_key_qbytes_2_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_3 = 8'hc + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_3_hi = local_offset_3[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_3_T = {match_key_qbytes_3_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_3_T_1 = {match_key_qbytes_3_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_3_T_2 = {match_key_qbytes_3_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_3084 = 8'h1 == _match_key_qbytes_3_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3085 = 8'h2 == _match_key_qbytes_3_T_2 ? phv_data_2 : _GEN_3084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3086 = 8'h3 == _match_key_qbytes_3_T_2 ? phv_data_3 : _GEN_3085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3087 = 8'h4 == _match_key_qbytes_3_T_2 ? phv_data_4 : _GEN_3086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3088 = 8'h5 == _match_key_qbytes_3_T_2 ? phv_data_5 : _GEN_3087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3089 = 8'h6 == _match_key_qbytes_3_T_2 ? phv_data_6 : _GEN_3088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3090 = 8'h7 == _match_key_qbytes_3_T_2 ? phv_data_7 : _GEN_3089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3091 = 8'h8 == _match_key_qbytes_3_T_2 ? phv_data_8 : _GEN_3090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3092 = 8'h9 == _match_key_qbytes_3_T_2 ? phv_data_9 : _GEN_3091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3093 = 8'ha == _match_key_qbytes_3_T_2 ? phv_data_10 : _GEN_3092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3094 = 8'hb == _match_key_qbytes_3_T_2 ? phv_data_11 : _GEN_3093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3095 = 8'hc == _match_key_qbytes_3_T_2 ? phv_data_12 : _GEN_3094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3096 = 8'hd == _match_key_qbytes_3_T_2 ? phv_data_13 : _GEN_3095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3097 = 8'he == _match_key_qbytes_3_T_2 ? phv_data_14 : _GEN_3096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3098 = 8'hf == _match_key_qbytes_3_T_2 ? phv_data_15 : _GEN_3097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3099 = 8'h10 == _match_key_qbytes_3_T_2 ? phv_data_16 : _GEN_3098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3100 = 8'h11 == _match_key_qbytes_3_T_2 ? phv_data_17 : _GEN_3099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3101 = 8'h12 == _match_key_qbytes_3_T_2 ? phv_data_18 : _GEN_3100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3102 = 8'h13 == _match_key_qbytes_3_T_2 ? phv_data_19 : _GEN_3101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3103 = 8'h14 == _match_key_qbytes_3_T_2 ? phv_data_20 : _GEN_3102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3104 = 8'h15 == _match_key_qbytes_3_T_2 ? phv_data_21 : _GEN_3103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3105 = 8'h16 == _match_key_qbytes_3_T_2 ? phv_data_22 : _GEN_3104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3106 = 8'h17 == _match_key_qbytes_3_T_2 ? phv_data_23 : _GEN_3105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3107 = 8'h18 == _match_key_qbytes_3_T_2 ? phv_data_24 : _GEN_3106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3108 = 8'h19 == _match_key_qbytes_3_T_2 ? phv_data_25 : _GEN_3107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3109 = 8'h1a == _match_key_qbytes_3_T_2 ? phv_data_26 : _GEN_3108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3110 = 8'h1b == _match_key_qbytes_3_T_2 ? phv_data_27 : _GEN_3109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3111 = 8'h1c == _match_key_qbytes_3_T_2 ? phv_data_28 : _GEN_3110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3112 = 8'h1d == _match_key_qbytes_3_T_2 ? phv_data_29 : _GEN_3111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3113 = 8'h1e == _match_key_qbytes_3_T_2 ? phv_data_30 : _GEN_3112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3114 = 8'h1f == _match_key_qbytes_3_T_2 ? phv_data_31 : _GEN_3113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3115 = 8'h20 == _match_key_qbytes_3_T_2 ? phv_data_32 : _GEN_3114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3116 = 8'h21 == _match_key_qbytes_3_T_2 ? phv_data_33 : _GEN_3115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3117 = 8'h22 == _match_key_qbytes_3_T_2 ? phv_data_34 : _GEN_3116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3118 = 8'h23 == _match_key_qbytes_3_T_2 ? phv_data_35 : _GEN_3117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3119 = 8'h24 == _match_key_qbytes_3_T_2 ? phv_data_36 : _GEN_3118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3120 = 8'h25 == _match_key_qbytes_3_T_2 ? phv_data_37 : _GEN_3119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3121 = 8'h26 == _match_key_qbytes_3_T_2 ? phv_data_38 : _GEN_3120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3122 = 8'h27 == _match_key_qbytes_3_T_2 ? phv_data_39 : _GEN_3121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3123 = 8'h28 == _match_key_qbytes_3_T_2 ? phv_data_40 : _GEN_3122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3124 = 8'h29 == _match_key_qbytes_3_T_2 ? phv_data_41 : _GEN_3123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3125 = 8'h2a == _match_key_qbytes_3_T_2 ? phv_data_42 : _GEN_3124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3126 = 8'h2b == _match_key_qbytes_3_T_2 ? phv_data_43 : _GEN_3125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3127 = 8'h2c == _match_key_qbytes_3_T_2 ? phv_data_44 : _GEN_3126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3128 = 8'h2d == _match_key_qbytes_3_T_2 ? phv_data_45 : _GEN_3127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3129 = 8'h2e == _match_key_qbytes_3_T_2 ? phv_data_46 : _GEN_3128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3130 = 8'h2f == _match_key_qbytes_3_T_2 ? phv_data_47 : _GEN_3129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3131 = 8'h30 == _match_key_qbytes_3_T_2 ? phv_data_48 : _GEN_3130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3132 = 8'h31 == _match_key_qbytes_3_T_2 ? phv_data_49 : _GEN_3131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3133 = 8'h32 == _match_key_qbytes_3_T_2 ? phv_data_50 : _GEN_3132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3134 = 8'h33 == _match_key_qbytes_3_T_2 ? phv_data_51 : _GEN_3133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3135 = 8'h34 == _match_key_qbytes_3_T_2 ? phv_data_52 : _GEN_3134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3136 = 8'h35 == _match_key_qbytes_3_T_2 ? phv_data_53 : _GEN_3135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3137 = 8'h36 == _match_key_qbytes_3_T_2 ? phv_data_54 : _GEN_3136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3138 = 8'h37 == _match_key_qbytes_3_T_2 ? phv_data_55 : _GEN_3137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3139 = 8'h38 == _match_key_qbytes_3_T_2 ? phv_data_56 : _GEN_3138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3140 = 8'h39 == _match_key_qbytes_3_T_2 ? phv_data_57 : _GEN_3139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3141 = 8'h3a == _match_key_qbytes_3_T_2 ? phv_data_58 : _GEN_3140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3142 = 8'h3b == _match_key_qbytes_3_T_2 ? phv_data_59 : _GEN_3141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3143 = 8'h3c == _match_key_qbytes_3_T_2 ? phv_data_60 : _GEN_3142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3144 = 8'h3d == _match_key_qbytes_3_T_2 ? phv_data_61 : _GEN_3143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3145 = 8'h3e == _match_key_qbytes_3_T_2 ? phv_data_62 : _GEN_3144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3146 = 8'h3f == _match_key_qbytes_3_T_2 ? phv_data_63 : _GEN_3145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3147 = 8'h40 == _match_key_qbytes_3_T_2 ? phv_data_64 : _GEN_3146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3148 = 8'h41 == _match_key_qbytes_3_T_2 ? phv_data_65 : _GEN_3147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3149 = 8'h42 == _match_key_qbytes_3_T_2 ? phv_data_66 : _GEN_3148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3150 = 8'h43 == _match_key_qbytes_3_T_2 ? phv_data_67 : _GEN_3149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3151 = 8'h44 == _match_key_qbytes_3_T_2 ? phv_data_68 : _GEN_3150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3152 = 8'h45 == _match_key_qbytes_3_T_2 ? phv_data_69 : _GEN_3151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3153 = 8'h46 == _match_key_qbytes_3_T_2 ? phv_data_70 : _GEN_3152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3154 = 8'h47 == _match_key_qbytes_3_T_2 ? phv_data_71 : _GEN_3153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3155 = 8'h48 == _match_key_qbytes_3_T_2 ? phv_data_72 : _GEN_3154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3156 = 8'h49 == _match_key_qbytes_3_T_2 ? phv_data_73 : _GEN_3155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3157 = 8'h4a == _match_key_qbytes_3_T_2 ? phv_data_74 : _GEN_3156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3158 = 8'h4b == _match_key_qbytes_3_T_2 ? phv_data_75 : _GEN_3157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3159 = 8'h4c == _match_key_qbytes_3_T_2 ? phv_data_76 : _GEN_3158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3160 = 8'h4d == _match_key_qbytes_3_T_2 ? phv_data_77 : _GEN_3159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3161 = 8'h4e == _match_key_qbytes_3_T_2 ? phv_data_78 : _GEN_3160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3162 = 8'h4f == _match_key_qbytes_3_T_2 ? phv_data_79 : _GEN_3161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3163 = 8'h50 == _match_key_qbytes_3_T_2 ? phv_data_80 : _GEN_3162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3164 = 8'h51 == _match_key_qbytes_3_T_2 ? phv_data_81 : _GEN_3163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3165 = 8'h52 == _match_key_qbytes_3_T_2 ? phv_data_82 : _GEN_3164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3166 = 8'h53 == _match_key_qbytes_3_T_2 ? phv_data_83 : _GEN_3165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3167 = 8'h54 == _match_key_qbytes_3_T_2 ? phv_data_84 : _GEN_3166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3168 = 8'h55 == _match_key_qbytes_3_T_2 ? phv_data_85 : _GEN_3167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3169 = 8'h56 == _match_key_qbytes_3_T_2 ? phv_data_86 : _GEN_3168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3170 = 8'h57 == _match_key_qbytes_3_T_2 ? phv_data_87 : _GEN_3169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3171 = 8'h58 == _match_key_qbytes_3_T_2 ? phv_data_88 : _GEN_3170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3172 = 8'h59 == _match_key_qbytes_3_T_2 ? phv_data_89 : _GEN_3171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3173 = 8'h5a == _match_key_qbytes_3_T_2 ? phv_data_90 : _GEN_3172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3174 = 8'h5b == _match_key_qbytes_3_T_2 ? phv_data_91 : _GEN_3173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3175 = 8'h5c == _match_key_qbytes_3_T_2 ? phv_data_92 : _GEN_3174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3176 = 8'h5d == _match_key_qbytes_3_T_2 ? phv_data_93 : _GEN_3175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3177 = 8'h5e == _match_key_qbytes_3_T_2 ? phv_data_94 : _GEN_3176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3178 = 8'h5f == _match_key_qbytes_3_T_2 ? phv_data_95 : _GEN_3177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3179 = 8'h60 == _match_key_qbytes_3_T_2 ? phv_data_96 : _GEN_3178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3180 = 8'h61 == _match_key_qbytes_3_T_2 ? phv_data_97 : _GEN_3179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3181 = 8'h62 == _match_key_qbytes_3_T_2 ? phv_data_98 : _GEN_3180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3182 = 8'h63 == _match_key_qbytes_3_T_2 ? phv_data_99 : _GEN_3181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3183 = 8'h64 == _match_key_qbytes_3_T_2 ? phv_data_100 : _GEN_3182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3184 = 8'h65 == _match_key_qbytes_3_T_2 ? phv_data_101 : _GEN_3183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3185 = 8'h66 == _match_key_qbytes_3_T_2 ? phv_data_102 : _GEN_3184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3186 = 8'h67 == _match_key_qbytes_3_T_2 ? phv_data_103 : _GEN_3185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3187 = 8'h68 == _match_key_qbytes_3_T_2 ? phv_data_104 : _GEN_3186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3188 = 8'h69 == _match_key_qbytes_3_T_2 ? phv_data_105 : _GEN_3187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3189 = 8'h6a == _match_key_qbytes_3_T_2 ? phv_data_106 : _GEN_3188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3190 = 8'h6b == _match_key_qbytes_3_T_2 ? phv_data_107 : _GEN_3189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3191 = 8'h6c == _match_key_qbytes_3_T_2 ? phv_data_108 : _GEN_3190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3192 = 8'h6d == _match_key_qbytes_3_T_2 ? phv_data_109 : _GEN_3191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3193 = 8'h6e == _match_key_qbytes_3_T_2 ? phv_data_110 : _GEN_3192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3194 = 8'h6f == _match_key_qbytes_3_T_2 ? phv_data_111 : _GEN_3193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3195 = 8'h70 == _match_key_qbytes_3_T_2 ? phv_data_112 : _GEN_3194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3196 = 8'h71 == _match_key_qbytes_3_T_2 ? phv_data_113 : _GEN_3195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3197 = 8'h72 == _match_key_qbytes_3_T_2 ? phv_data_114 : _GEN_3196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3198 = 8'h73 == _match_key_qbytes_3_T_2 ? phv_data_115 : _GEN_3197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3199 = 8'h74 == _match_key_qbytes_3_T_2 ? phv_data_116 : _GEN_3198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3200 = 8'h75 == _match_key_qbytes_3_T_2 ? phv_data_117 : _GEN_3199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3201 = 8'h76 == _match_key_qbytes_3_T_2 ? phv_data_118 : _GEN_3200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3202 = 8'h77 == _match_key_qbytes_3_T_2 ? phv_data_119 : _GEN_3201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3203 = 8'h78 == _match_key_qbytes_3_T_2 ? phv_data_120 : _GEN_3202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3204 = 8'h79 == _match_key_qbytes_3_T_2 ? phv_data_121 : _GEN_3203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3205 = 8'h7a == _match_key_qbytes_3_T_2 ? phv_data_122 : _GEN_3204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3206 = 8'h7b == _match_key_qbytes_3_T_2 ? phv_data_123 : _GEN_3205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3207 = 8'h7c == _match_key_qbytes_3_T_2 ? phv_data_124 : _GEN_3206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3208 = 8'h7d == _match_key_qbytes_3_T_2 ? phv_data_125 : _GEN_3207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3209 = 8'h7e == _match_key_qbytes_3_T_2 ? phv_data_126 : _GEN_3208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3210 = 8'h7f == _match_key_qbytes_3_T_2 ? phv_data_127 : _GEN_3209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3211 = 8'h80 == _match_key_qbytes_3_T_2 ? phv_data_128 : _GEN_3210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3212 = 8'h81 == _match_key_qbytes_3_T_2 ? phv_data_129 : _GEN_3211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3213 = 8'h82 == _match_key_qbytes_3_T_2 ? phv_data_130 : _GEN_3212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3214 = 8'h83 == _match_key_qbytes_3_T_2 ? phv_data_131 : _GEN_3213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3215 = 8'h84 == _match_key_qbytes_3_T_2 ? phv_data_132 : _GEN_3214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3216 = 8'h85 == _match_key_qbytes_3_T_2 ? phv_data_133 : _GEN_3215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3217 = 8'h86 == _match_key_qbytes_3_T_2 ? phv_data_134 : _GEN_3216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3218 = 8'h87 == _match_key_qbytes_3_T_2 ? phv_data_135 : _GEN_3217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3219 = 8'h88 == _match_key_qbytes_3_T_2 ? phv_data_136 : _GEN_3218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3220 = 8'h89 == _match_key_qbytes_3_T_2 ? phv_data_137 : _GEN_3219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3221 = 8'h8a == _match_key_qbytes_3_T_2 ? phv_data_138 : _GEN_3220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3222 = 8'h8b == _match_key_qbytes_3_T_2 ? phv_data_139 : _GEN_3221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3223 = 8'h8c == _match_key_qbytes_3_T_2 ? phv_data_140 : _GEN_3222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3224 = 8'h8d == _match_key_qbytes_3_T_2 ? phv_data_141 : _GEN_3223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3225 = 8'h8e == _match_key_qbytes_3_T_2 ? phv_data_142 : _GEN_3224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3226 = 8'h8f == _match_key_qbytes_3_T_2 ? phv_data_143 : _GEN_3225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3227 = 8'h90 == _match_key_qbytes_3_T_2 ? phv_data_144 : _GEN_3226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3228 = 8'h91 == _match_key_qbytes_3_T_2 ? phv_data_145 : _GEN_3227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3229 = 8'h92 == _match_key_qbytes_3_T_2 ? phv_data_146 : _GEN_3228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3230 = 8'h93 == _match_key_qbytes_3_T_2 ? phv_data_147 : _GEN_3229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3231 = 8'h94 == _match_key_qbytes_3_T_2 ? phv_data_148 : _GEN_3230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3232 = 8'h95 == _match_key_qbytes_3_T_2 ? phv_data_149 : _GEN_3231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3233 = 8'h96 == _match_key_qbytes_3_T_2 ? phv_data_150 : _GEN_3232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3234 = 8'h97 == _match_key_qbytes_3_T_2 ? phv_data_151 : _GEN_3233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3235 = 8'h98 == _match_key_qbytes_3_T_2 ? phv_data_152 : _GEN_3234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3236 = 8'h99 == _match_key_qbytes_3_T_2 ? phv_data_153 : _GEN_3235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3237 = 8'h9a == _match_key_qbytes_3_T_2 ? phv_data_154 : _GEN_3236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3238 = 8'h9b == _match_key_qbytes_3_T_2 ? phv_data_155 : _GEN_3237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3239 = 8'h9c == _match_key_qbytes_3_T_2 ? phv_data_156 : _GEN_3238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3240 = 8'h9d == _match_key_qbytes_3_T_2 ? phv_data_157 : _GEN_3239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3241 = 8'h9e == _match_key_qbytes_3_T_2 ? phv_data_158 : _GEN_3240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3242 = 8'h9f == _match_key_qbytes_3_T_2 ? phv_data_159 : _GEN_3241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3243 = 8'ha0 == _match_key_qbytes_3_T_2 ? phv_data_160 : _GEN_3242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3244 = 8'ha1 == _match_key_qbytes_3_T_2 ? phv_data_161 : _GEN_3243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3245 = 8'ha2 == _match_key_qbytes_3_T_2 ? phv_data_162 : _GEN_3244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3246 = 8'ha3 == _match_key_qbytes_3_T_2 ? phv_data_163 : _GEN_3245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3247 = 8'ha4 == _match_key_qbytes_3_T_2 ? phv_data_164 : _GEN_3246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3248 = 8'ha5 == _match_key_qbytes_3_T_2 ? phv_data_165 : _GEN_3247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3249 = 8'ha6 == _match_key_qbytes_3_T_2 ? phv_data_166 : _GEN_3248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3250 = 8'ha7 == _match_key_qbytes_3_T_2 ? phv_data_167 : _GEN_3249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3251 = 8'ha8 == _match_key_qbytes_3_T_2 ? phv_data_168 : _GEN_3250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3252 = 8'ha9 == _match_key_qbytes_3_T_2 ? phv_data_169 : _GEN_3251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3253 = 8'haa == _match_key_qbytes_3_T_2 ? phv_data_170 : _GEN_3252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3254 = 8'hab == _match_key_qbytes_3_T_2 ? phv_data_171 : _GEN_3253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3255 = 8'hac == _match_key_qbytes_3_T_2 ? phv_data_172 : _GEN_3254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3256 = 8'had == _match_key_qbytes_3_T_2 ? phv_data_173 : _GEN_3255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3257 = 8'hae == _match_key_qbytes_3_T_2 ? phv_data_174 : _GEN_3256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3258 = 8'haf == _match_key_qbytes_3_T_2 ? phv_data_175 : _GEN_3257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3259 = 8'hb0 == _match_key_qbytes_3_T_2 ? phv_data_176 : _GEN_3258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3260 = 8'hb1 == _match_key_qbytes_3_T_2 ? phv_data_177 : _GEN_3259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3261 = 8'hb2 == _match_key_qbytes_3_T_2 ? phv_data_178 : _GEN_3260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3262 = 8'hb3 == _match_key_qbytes_3_T_2 ? phv_data_179 : _GEN_3261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3263 = 8'hb4 == _match_key_qbytes_3_T_2 ? phv_data_180 : _GEN_3262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3264 = 8'hb5 == _match_key_qbytes_3_T_2 ? phv_data_181 : _GEN_3263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3265 = 8'hb6 == _match_key_qbytes_3_T_2 ? phv_data_182 : _GEN_3264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3266 = 8'hb7 == _match_key_qbytes_3_T_2 ? phv_data_183 : _GEN_3265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3267 = 8'hb8 == _match_key_qbytes_3_T_2 ? phv_data_184 : _GEN_3266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3268 = 8'hb9 == _match_key_qbytes_3_T_2 ? phv_data_185 : _GEN_3267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3269 = 8'hba == _match_key_qbytes_3_T_2 ? phv_data_186 : _GEN_3268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3270 = 8'hbb == _match_key_qbytes_3_T_2 ? phv_data_187 : _GEN_3269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3271 = 8'hbc == _match_key_qbytes_3_T_2 ? phv_data_188 : _GEN_3270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3272 = 8'hbd == _match_key_qbytes_3_T_2 ? phv_data_189 : _GEN_3271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3273 = 8'hbe == _match_key_qbytes_3_T_2 ? phv_data_190 : _GEN_3272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3274 = 8'hbf == _match_key_qbytes_3_T_2 ? phv_data_191 : _GEN_3273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3275 = 8'hc0 == _match_key_qbytes_3_T_2 ? phv_data_192 : _GEN_3274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3276 = 8'hc1 == _match_key_qbytes_3_T_2 ? phv_data_193 : _GEN_3275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3277 = 8'hc2 == _match_key_qbytes_3_T_2 ? phv_data_194 : _GEN_3276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3278 = 8'hc3 == _match_key_qbytes_3_T_2 ? phv_data_195 : _GEN_3277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3279 = 8'hc4 == _match_key_qbytes_3_T_2 ? phv_data_196 : _GEN_3278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3280 = 8'hc5 == _match_key_qbytes_3_T_2 ? phv_data_197 : _GEN_3279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3281 = 8'hc6 == _match_key_qbytes_3_T_2 ? phv_data_198 : _GEN_3280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3282 = 8'hc7 == _match_key_qbytes_3_T_2 ? phv_data_199 : _GEN_3281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3283 = 8'hc8 == _match_key_qbytes_3_T_2 ? phv_data_200 : _GEN_3282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3284 = 8'hc9 == _match_key_qbytes_3_T_2 ? phv_data_201 : _GEN_3283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3285 = 8'hca == _match_key_qbytes_3_T_2 ? phv_data_202 : _GEN_3284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3286 = 8'hcb == _match_key_qbytes_3_T_2 ? phv_data_203 : _GEN_3285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3287 = 8'hcc == _match_key_qbytes_3_T_2 ? phv_data_204 : _GEN_3286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3288 = 8'hcd == _match_key_qbytes_3_T_2 ? phv_data_205 : _GEN_3287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3289 = 8'hce == _match_key_qbytes_3_T_2 ? phv_data_206 : _GEN_3288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3290 = 8'hcf == _match_key_qbytes_3_T_2 ? phv_data_207 : _GEN_3289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3291 = 8'hd0 == _match_key_qbytes_3_T_2 ? phv_data_208 : _GEN_3290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3292 = 8'hd1 == _match_key_qbytes_3_T_2 ? phv_data_209 : _GEN_3291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3293 = 8'hd2 == _match_key_qbytes_3_T_2 ? phv_data_210 : _GEN_3292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3294 = 8'hd3 == _match_key_qbytes_3_T_2 ? phv_data_211 : _GEN_3293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3295 = 8'hd4 == _match_key_qbytes_3_T_2 ? phv_data_212 : _GEN_3294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3296 = 8'hd5 == _match_key_qbytes_3_T_2 ? phv_data_213 : _GEN_3295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3297 = 8'hd6 == _match_key_qbytes_3_T_2 ? phv_data_214 : _GEN_3296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3298 = 8'hd7 == _match_key_qbytes_3_T_2 ? phv_data_215 : _GEN_3297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3299 = 8'hd8 == _match_key_qbytes_3_T_2 ? phv_data_216 : _GEN_3298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3300 = 8'hd9 == _match_key_qbytes_3_T_2 ? phv_data_217 : _GEN_3299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3301 = 8'hda == _match_key_qbytes_3_T_2 ? phv_data_218 : _GEN_3300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3302 = 8'hdb == _match_key_qbytes_3_T_2 ? phv_data_219 : _GEN_3301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3303 = 8'hdc == _match_key_qbytes_3_T_2 ? phv_data_220 : _GEN_3302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3304 = 8'hdd == _match_key_qbytes_3_T_2 ? phv_data_221 : _GEN_3303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3305 = 8'hde == _match_key_qbytes_3_T_2 ? phv_data_222 : _GEN_3304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3306 = 8'hdf == _match_key_qbytes_3_T_2 ? phv_data_223 : _GEN_3305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3307 = 8'he0 == _match_key_qbytes_3_T_2 ? phv_data_224 : _GEN_3306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3308 = 8'he1 == _match_key_qbytes_3_T_2 ? phv_data_225 : _GEN_3307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3309 = 8'he2 == _match_key_qbytes_3_T_2 ? phv_data_226 : _GEN_3308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3310 = 8'he3 == _match_key_qbytes_3_T_2 ? phv_data_227 : _GEN_3309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3311 = 8'he4 == _match_key_qbytes_3_T_2 ? phv_data_228 : _GEN_3310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3312 = 8'he5 == _match_key_qbytes_3_T_2 ? phv_data_229 : _GEN_3311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3313 = 8'he6 == _match_key_qbytes_3_T_2 ? phv_data_230 : _GEN_3312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3314 = 8'he7 == _match_key_qbytes_3_T_2 ? phv_data_231 : _GEN_3313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3315 = 8'he8 == _match_key_qbytes_3_T_2 ? phv_data_232 : _GEN_3314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3316 = 8'he9 == _match_key_qbytes_3_T_2 ? phv_data_233 : _GEN_3315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3317 = 8'hea == _match_key_qbytes_3_T_2 ? phv_data_234 : _GEN_3316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3318 = 8'heb == _match_key_qbytes_3_T_2 ? phv_data_235 : _GEN_3317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3319 = 8'hec == _match_key_qbytes_3_T_2 ? phv_data_236 : _GEN_3318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3320 = 8'hed == _match_key_qbytes_3_T_2 ? phv_data_237 : _GEN_3319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3321 = 8'hee == _match_key_qbytes_3_T_2 ? phv_data_238 : _GEN_3320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3322 = 8'hef == _match_key_qbytes_3_T_2 ? phv_data_239 : _GEN_3321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3323 = 8'hf0 == _match_key_qbytes_3_T_2 ? phv_data_240 : _GEN_3322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3324 = 8'hf1 == _match_key_qbytes_3_T_2 ? phv_data_241 : _GEN_3323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3325 = 8'hf2 == _match_key_qbytes_3_T_2 ? phv_data_242 : _GEN_3324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3326 = 8'hf3 == _match_key_qbytes_3_T_2 ? phv_data_243 : _GEN_3325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3327 = 8'hf4 == _match_key_qbytes_3_T_2 ? phv_data_244 : _GEN_3326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3328 = 8'hf5 == _match_key_qbytes_3_T_2 ? phv_data_245 : _GEN_3327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3329 = 8'hf6 == _match_key_qbytes_3_T_2 ? phv_data_246 : _GEN_3328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3330 = 8'hf7 == _match_key_qbytes_3_T_2 ? phv_data_247 : _GEN_3329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3331 = 8'hf8 == _match_key_qbytes_3_T_2 ? phv_data_248 : _GEN_3330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3332 = 8'hf9 == _match_key_qbytes_3_T_2 ? phv_data_249 : _GEN_3331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3333 = 8'hfa == _match_key_qbytes_3_T_2 ? phv_data_250 : _GEN_3332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3334 = 8'hfb == _match_key_qbytes_3_T_2 ? phv_data_251 : _GEN_3333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3335 = 8'hfc == _match_key_qbytes_3_T_2 ? phv_data_252 : _GEN_3334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3336 = 8'hfd == _match_key_qbytes_3_T_2 ? phv_data_253 : _GEN_3335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3337 = 8'hfe == _match_key_qbytes_3_T_2 ? phv_data_254 : _GEN_3336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3338 = 8'hff == _match_key_qbytes_3_T_2 ? phv_data_255 : _GEN_3337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3340 = 8'h1 == local_offset_3 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3341 = 8'h2 == local_offset_3 ? phv_data_2 : _GEN_3340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3342 = 8'h3 == local_offset_3 ? phv_data_3 : _GEN_3341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3343 = 8'h4 == local_offset_3 ? phv_data_4 : _GEN_3342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3344 = 8'h5 == local_offset_3 ? phv_data_5 : _GEN_3343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3345 = 8'h6 == local_offset_3 ? phv_data_6 : _GEN_3344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3346 = 8'h7 == local_offset_3 ? phv_data_7 : _GEN_3345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3347 = 8'h8 == local_offset_3 ? phv_data_8 : _GEN_3346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3348 = 8'h9 == local_offset_3 ? phv_data_9 : _GEN_3347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3349 = 8'ha == local_offset_3 ? phv_data_10 : _GEN_3348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3350 = 8'hb == local_offset_3 ? phv_data_11 : _GEN_3349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3351 = 8'hc == local_offset_3 ? phv_data_12 : _GEN_3350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3352 = 8'hd == local_offset_3 ? phv_data_13 : _GEN_3351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3353 = 8'he == local_offset_3 ? phv_data_14 : _GEN_3352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3354 = 8'hf == local_offset_3 ? phv_data_15 : _GEN_3353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3355 = 8'h10 == local_offset_3 ? phv_data_16 : _GEN_3354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3356 = 8'h11 == local_offset_3 ? phv_data_17 : _GEN_3355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3357 = 8'h12 == local_offset_3 ? phv_data_18 : _GEN_3356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3358 = 8'h13 == local_offset_3 ? phv_data_19 : _GEN_3357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3359 = 8'h14 == local_offset_3 ? phv_data_20 : _GEN_3358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3360 = 8'h15 == local_offset_3 ? phv_data_21 : _GEN_3359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3361 = 8'h16 == local_offset_3 ? phv_data_22 : _GEN_3360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3362 = 8'h17 == local_offset_3 ? phv_data_23 : _GEN_3361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3363 = 8'h18 == local_offset_3 ? phv_data_24 : _GEN_3362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3364 = 8'h19 == local_offset_3 ? phv_data_25 : _GEN_3363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3365 = 8'h1a == local_offset_3 ? phv_data_26 : _GEN_3364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3366 = 8'h1b == local_offset_3 ? phv_data_27 : _GEN_3365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3367 = 8'h1c == local_offset_3 ? phv_data_28 : _GEN_3366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3368 = 8'h1d == local_offset_3 ? phv_data_29 : _GEN_3367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3369 = 8'h1e == local_offset_3 ? phv_data_30 : _GEN_3368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3370 = 8'h1f == local_offset_3 ? phv_data_31 : _GEN_3369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3371 = 8'h20 == local_offset_3 ? phv_data_32 : _GEN_3370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3372 = 8'h21 == local_offset_3 ? phv_data_33 : _GEN_3371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3373 = 8'h22 == local_offset_3 ? phv_data_34 : _GEN_3372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3374 = 8'h23 == local_offset_3 ? phv_data_35 : _GEN_3373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3375 = 8'h24 == local_offset_3 ? phv_data_36 : _GEN_3374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3376 = 8'h25 == local_offset_3 ? phv_data_37 : _GEN_3375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3377 = 8'h26 == local_offset_3 ? phv_data_38 : _GEN_3376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3378 = 8'h27 == local_offset_3 ? phv_data_39 : _GEN_3377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3379 = 8'h28 == local_offset_3 ? phv_data_40 : _GEN_3378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3380 = 8'h29 == local_offset_3 ? phv_data_41 : _GEN_3379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3381 = 8'h2a == local_offset_3 ? phv_data_42 : _GEN_3380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3382 = 8'h2b == local_offset_3 ? phv_data_43 : _GEN_3381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3383 = 8'h2c == local_offset_3 ? phv_data_44 : _GEN_3382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3384 = 8'h2d == local_offset_3 ? phv_data_45 : _GEN_3383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3385 = 8'h2e == local_offset_3 ? phv_data_46 : _GEN_3384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3386 = 8'h2f == local_offset_3 ? phv_data_47 : _GEN_3385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3387 = 8'h30 == local_offset_3 ? phv_data_48 : _GEN_3386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3388 = 8'h31 == local_offset_3 ? phv_data_49 : _GEN_3387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3389 = 8'h32 == local_offset_3 ? phv_data_50 : _GEN_3388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3390 = 8'h33 == local_offset_3 ? phv_data_51 : _GEN_3389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3391 = 8'h34 == local_offset_3 ? phv_data_52 : _GEN_3390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3392 = 8'h35 == local_offset_3 ? phv_data_53 : _GEN_3391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3393 = 8'h36 == local_offset_3 ? phv_data_54 : _GEN_3392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3394 = 8'h37 == local_offset_3 ? phv_data_55 : _GEN_3393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3395 = 8'h38 == local_offset_3 ? phv_data_56 : _GEN_3394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3396 = 8'h39 == local_offset_3 ? phv_data_57 : _GEN_3395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3397 = 8'h3a == local_offset_3 ? phv_data_58 : _GEN_3396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3398 = 8'h3b == local_offset_3 ? phv_data_59 : _GEN_3397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3399 = 8'h3c == local_offset_3 ? phv_data_60 : _GEN_3398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3400 = 8'h3d == local_offset_3 ? phv_data_61 : _GEN_3399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3401 = 8'h3e == local_offset_3 ? phv_data_62 : _GEN_3400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3402 = 8'h3f == local_offset_3 ? phv_data_63 : _GEN_3401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3403 = 8'h40 == local_offset_3 ? phv_data_64 : _GEN_3402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3404 = 8'h41 == local_offset_3 ? phv_data_65 : _GEN_3403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3405 = 8'h42 == local_offset_3 ? phv_data_66 : _GEN_3404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3406 = 8'h43 == local_offset_3 ? phv_data_67 : _GEN_3405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3407 = 8'h44 == local_offset_3 ? phv_data_68 : _GEN_3406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3408 = 8'h45 == local_offset_3 ? phv_data_69 : _GEN_3407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3409 = 8'h46 == local_offset_3 ? phv_data_70 : _GEN_3408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3410 = 8'h47 == local_offset_3 ? phv_data_71 : _GEN_3409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3411 = 8'h48 == local_offset_3 ? phv_data_72 : _GEN_3410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3412 = 8'h49 == local_offset_3 ? phv_data_73 : _GEN_3411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3413 = 8'h4a == local_offset_3 ? phv_data_74 : _GEN_3412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3414 = 8'h4b == local_offset_3 ? phv_data_75 : _GEN_3413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3415 = 8'h4c == local_offset_3 ? phv_data_76 : _GEN_3414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3416 = 8'h4d == local_offset_3 ? phv_data_77 : _GEN_3415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3417 = 8'h4e == local_offset_3 ? phv_data_78 : _GEN_3416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3418 = 8'h4f == local_offset_3 ? phv_data_79 : _GEN_3417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3419 = 8'h50 == local_offset_3 ? phv_data_80 : _GEN_3418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3420 = 8'h51 == local_offset_3 ? phv_data_81 : _GEN_3419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3421 = 8'h52 == local_offset_3 ? phv_data_82 : _GEN_3420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3422 = 8'h53 == local_offset_3 ? phv_data_83 : _GEN_3421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3423 = 8'h54 == local_offset_3 ? phv_data_84 : _GEN_3422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3424 = 8'h55 == local_offset_3 ? phv_data_85 : _GEN_3423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3425 = 8'h56 == local_offset_3 ? phv_data_86 : _GEN_3424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3426 = 8'h57 == local_offset_3 ? phv_data_87 : _GEN_3425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3427 = 8'h58 == local_offset_3 ? phv_data_88 : _GEN_3426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3428 = 8'h59 == local_offset_3 ? phv_data_89 : _GEN_3427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3429 = 8'h5a == local_offset_3 ? phv_data_90 : _GEN_3428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3430 = 8'h5b == local_offset_3 ? phv_data_91 : _GEN_3429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3431 = 8'h5c == local_offset_3 ? phv_data_92 : _GEN_3430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3432 = 8'h5d == local_offset_3 ? phv_data_93 : _GEN_3431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3433 = 8'h5e == local_offset_3 ? phv_data_94 : _GEN_3432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3434 = 8'h5f == local_offset_3 ? phv_data_95 : _GEN_3433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3435 = 8'h60 == local_offset_3 ? phv_data_96 : _GEN_3434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3436 = 8'h61 == local_offset_3 ? phv_data_97 : _GEN_3435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3437 = 8'h62 == local_offset_3 ? phv_data_98 : _GEN_3436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3438 = 8'h63 == local_offset_3 ? phv_data_99 : _GEN_3437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3439 = 8'h64 == local_offset_3 ? phv_data_100 : _GEN_3438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3440 = 8'h65 == local_offset_3 ? phv_data_101 : _GEN_3439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3441 = 8'h66 == local_offset_3 ? phv_data_102 : _GEN_3440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3442 = 8'h67 == local_offset_3 ? phv_data_103 : _GEN_3441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3443 = 8'h68 == local_offset_3 ? phv_data_104 : _GEN_3442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3444 = 8'h69 == local_offset_3 ? phv_data_105 : _GEN_3443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3445 = 8'h6a == local_offset_3 ? phv_data_106 : _GEN_3444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3446 = 8'h6b == local_offset_3 ? phv_data_107 : _GEN_3445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3447 = 8'h6c == local_offset_3 ? phv_data_108 : _GEN_3446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3448 = 8'h6d == local_offset_3 ? phv_data_109 : _GEN_3447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3449 = 8'h6e == local_offset_3 ? phv_data_110 : _GEN_3448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3450 = 8'h6f == local_offset_3 ? phv_data_111 : _GEN_3449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3451 = 8'h70 == local_offset_3 ? phv_data_112 : _GEN_3450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3452 = 8'h71 == local_offset_3 ? phv_data_113 : _GEN_3451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3453 = 8'h72 == local_offset_3 ? phv_data_114 : _GEN_3452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3454 = 8'h73 == local_offset_3 ? phv_data_115 : _GEN_3453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3455 = 8'h74 == local_offset_3 ? phv_data_116 : _GEN_3454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3456 = 8'h75 == local_offset_3 ? phv_data_117 : _GEN_3455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3457 = 8'h76 == local_offset_3 ? phv_data_118 : _GEN_3456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3458 = 8'h77 == local_offset_3 ? phv_data_119 : _GEN_3457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3459 = 8'h78 == local_offset_3 ? phv_data_120 : _GEN_3458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3460 = 8'h79 == local_offset_3 ? phv_data_121 : _GEN_3459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3461 = 8'h7a == local_offset_3 ? phv_data_122 : _GEN_3460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3462 = 8'h7b == local_offset_3 ? phv_data_123 : _GEN_3461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3463 = 8'h7c == local_offset_3 ? phv_data_124 : _GEN_3462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3464 = 8'h7d == local_offset_3 ? phv_data_125 : _GEN_3463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3465 = 8'h7e == local_offset_3 ? phv_data_126 : _GEN_3464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3466 = 8'h7f == local_offset_3 ? phv_data_127 : _GEN_3465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3467 = 8'h80 == local_offset_3 ? phv_data_128 : _GEN_3466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3468 = 8'h81 == local_offset_3 ? phv_data_129 : _GEN_3467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3469 = 8'h82 == local_offset_3 ? phv_data_130 : _GEN_3468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3470 = 8'h83 == local_offset_3 ? phv_data_131 : _GEN_3469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3471 = 8'h84 == local_offset_3 ? phv_data_132 : _GEN_3470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3472 = 8'h85 == local_offset_3 ? phv_data_133 : _GEN_3471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3473 = 8'h86 == local_offset_3 ? phv_data_134 : _GEN_3472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3474 = 8'h87 == local_offset_3 ? phv_data_135 : _GEN_3473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3475 = 8'h88 == local_offset_3 ? phv_data_136 : _GEN_3474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3476 = 8'h89 == local_offset_3 ? phv_data_137 : _GEN_3475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3477 = 8'h8a == local_offset_3 ? phv_data_138 : _GEN_3476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3478 = 8'h8b == local_offset_3 ? phv_data_139 : _GEN_3477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3479 = 8'h8c == local_offset_3 ? phv_data_140 : _GEN_3478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3480 = 8'h8d == local_offset_3 ? phv_data_141 : _GEN_3479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3481 = 8'h8e == local_offset_3 ? phv_data_142 : _GEN_3480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3482 = 8'h8f == local_offset_3 ? phv_data_143 : _GEN_3481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3483 = 8'h90 == local_offset_3 ? phv_data_144 : _GEN_3482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3484 = 8'h91 == local_offset_3 ? phv_data_145 : _GEN_3483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3485 = 8'h92 == local_offset_3 ? phv_data_146 : _GEN_3484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3486 = 8'h93 == local_offset_3 ? phv_data_147 : _GEN_3485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3487 = 8'h94 == local_offset_3 ? phv_data_148 : _GEN_3486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3488 = 8'h95 == local_offset_3 ? phv_data_149 : _GEN_3487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3489 = 8'h96 == local_offset_3 ? phv_data_150 : _GEN_3488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3490 = 8'h97 == local_offset_3 ? phv_data_151 : _GEN_3489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3491 = 8'h98 == local_offset_3 ? phv_data_152 : _GEN_3490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3492 = 8'h99 == local_offset_3 ? phv_data_153 : _GEN_3491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3493 = 8'h9a == local_offset_3 ? phv_data_154 : _GEN_3492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3494 = 8'h9b == local_offset_3 ? phv_data_155 : _GEN_3493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3495 = 8'h9c == local_offset_3 ? phv_data_156 : _GEN_3494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3496 = 8'h9d == local_offset_3 ? phv_data_157 : _GEN_3495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3497 = 8'h9e == local_offset_3 ? phv_data_158 : _GEN_3496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3498 = 8'h9f == local_offset_3 ? phv_data_159 : _GEN_3497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3499 = 8'ha0 == local_offset_3 ? phv_data_160 : _GEN_3498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3500 = 8'ha1 == local_offset_3 ? phv_data_161 : _GEN_3499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3501 = 8'ha2 == local_offset_3 ? phv_data_162 : _GEN_3500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3502 = 8'ha3 == local_offset_3 ? phv_data_163 : _GEN_3501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3503 = 8'ha4 == local_offset_3 ? phv_data_164 : _GEN_3502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3504 = 8'ha5 == local_offset_3 ? phv_data_165 : _GEN_3503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3505 = 8'ha6 == local_offset_3 ? phv_data_166 : _GEN_3504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3506 = 8'ha7 == local_offset_3 ? phv_data_167 : _GEN_3505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3507 = 8'ha8 == local_offset_3 ? phv_data_168 : _GEN_3506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3508 = 8'ha9 == local_offset_3 ? phv_data_169 : _GEN_3507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3509 = 8'haa == local_offset_3 ? phv_data_170 : _GEN_3508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3510 = 8'hab == local_offset_3 ? phv_data_171 : _GEN_3509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3511 = 8'hac == local_offset_3 ? phv_data_172 : _GEN_3510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3512 = 8'had == local_offset_3 ? phv_data_173 : _GEN_3511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3513 = 8'hae == local_offset_3 ? phv_data_174 : _GEN_3512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3514 = 8'haf == local_offset_3 ? phv_data_175 : _GEN_3513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3515 = 8'hb0 == local_offset_3 ? phv_data_176 : _GEN_3514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3516 = 8'hb1 == local_offset_3 ? phv_data_177 : _GEN_3515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3517 = 8'hb2 == local_offset_3 ? phv_data_178 : _GEN_3516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3518 = 8'hb3 == local_offset_3 ? phv_data_179 : _GEN_3517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3519 = 8'hb4 == local_offset_3 ? phv_data_180 : _GEN_3518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3520 = 8'hb5 == local_offset_3 ? phv_data_181 : _GEN_3519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3521 = 8'hb6 == local_offset_3 ? phv_data_182 : _GEN_3520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3522 = 8'hb7 == local_offset_3 ? phv_data_183 : _GEN_3521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3523 = 8'hb8 == local_offset_3 ? phv_data_184 : _GEN_3522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3524 = 8'hb9 == local_offset_3 ? phv_data_185 : _GEN_3523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3525 = 8'hba == local_offset_3 ? phv_data_186 : _GEN_3524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3526 = 8'hbb == local_offset_3 ? phv_data_187 : _GEN_3525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3527 = 8'hbc == local_offset_3 ? phv_data_188 : _GEN_3526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3528 = 8'hbd == local_offset_3 ? phv_data_189 : _GEN_3527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3529 = 8'hbe == local_offset_3 ? phv_data_190 : _GEN_3528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3530 = 8'hbf == local_offset_3 ? phv_data_191 : _GEN_3529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3531 = 8'hc0 == local_offset_3 ? phv_data_192 : _GEN_3530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3532 = 8'hc1 == local_offset_3 ? phv_data_193 : _GEN_3531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3533 = 8'hc2 == local_offset_3 ? phv_data_194 : _GEN_3532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3534 = 8'hc3 == local_offset_3 ? phv_data_195 : _GEN_3533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3535 = 8'hc4 == local_offset_3 ? phv_data_196 : _GEN_3534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3536 = 8'hc5 == local_offset_3 ? phv_data_197 : _GEN_3535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3537 = 8'hc6 == local_offset_3 ? phv_data_198 : _GEN_3536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3538 = 8'hc7 == local_offset_3 ? phv_data_199 : _GEN_3537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3539 = 8'hc8 == local_offset_3 ? phv_data_200 : _GEN_3538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3540 = 8'hc9 == local_offset_3 ? phv_data_201 : _GEN_3539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3541 = 8'hca == local_offset_3 ? phv_data_202 : _GEN_3540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3542 = 8'hcb == local_offset_3 ? phv_data_203 : _GEN_3541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3543 = 8'hcc == local_offset_3 ? phv_data_204 : _GEN_3542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3544 = 8'hcd == local_offset_3 ? phv_data_205 : _GEN_3543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3545 = 8'hce == local_offset_3 ? phv_data_206 : _GEN_3544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3546 = 8'hcf == local_offset_3 ? phv_data_207 : _GEN_3545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3547 = 8'hd0 == local_offset_3 ? phv_data_208 : _GEN_3546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3548 = 8'hd1 == local_offset_3 ? phv_data_209 : _GEN_3547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3549 = 8'hd2 == local_offset_3 ? phv_data_210 : _GEN_3548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3550 = 8'hd3 == local_offset_3 ? phv_data_211 : _GEN_3549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3551 = 8'hd4 == local_offset_3 ? phv_data_212 : _GEN_3550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3552 = 8'hd5 == local_offset_3 ? phv_data_213 : _GEN_3551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3553 = 8'hd6 == local_offset_3 ? phv_data_214 : _GEN_3552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3554 = 8'hd7 == local_offset_3 ? phv_data_215 : _GEN_3553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3555 = 8'hd8 == local_offset_3 ? phv_data_216 : _GEN_3554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3556 = 8'hd9 == local_offset_3 ? phv_data_217 : _GEN_3555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3557 = 8'hda == local_offset_3 ? phv_data_218 : _GEN_3556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3558 = 8'hdb == local_offset_3 ? phv_data_219 : _GEN_3557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3559 = 8'hdc == local_offset_3 ? phv_data_220 : _GEN_3558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3560 = 8'hdd == local_offset_3 ? phv_data_221 : _GEN_3559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3561 = 8'hde == local_offset_3 ? phv_data_222 : _GEN_3560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3562 = 8'hdf == local_offset_3 ? phv_data_223 : _GEN_3561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3563 = 8'he0 == local_offset_3 ? phv_data_224 : _GEN_3562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3564 = 8'he1 == local_offset_3 ? phv_data_225 : _GEN_3563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3565 = 8'he2 == local_offset_3 ? phv_data_226 : _GEN_3564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3566 = 8'he3 == local_offset_3 ? phv_data_227 : _GEN_3565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3567 = 8'he4 == local_offset_3 ? phv_data_228 : _GEN_3566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3568 = 8'he5 == local_offset_3 ? phv_data_229 : _GEN_3567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3569 = 8'he6 == local_offset_3 ? phv_data_230 : _GEN_3568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3570 = 8'he7 == local_offset_3 ? phv_data_231 : _GEN_3569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3571 = 8'he8 == local_offset_3 ? phv_data_232 : _GEN_3570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3572 = 8'he9 == local_offset_3 ? phv_data_233 : _GEN_3571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3573 = 8'hea == local_offset_3 ? phv_data_234 : _GEN_3572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3574 = 8'heb == local_offset_3 ? phv_data_235 : _GEN_3573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3575 = 8'hec == local_offset_3 ? phv_data_236 : _GEN_3574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3576 = 8'hed == local_offset_3 ? phv_data_237 : _GEN_3575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3577 = 8'hee == local_offset_3 ? phv_data_238 : _GEN_3576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3578 = 8'hef == local_offset_3 ? phv_data_239 : _GEN_3577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3579 = 8'hf0 == local_offset_3 ? phv_data_240 : _GEN_3578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3580 = 8'hf1 == local_offset_3 ? phv_data_241 : _GEN_3579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3581 = 8'hf2 == local_offset_3 ? phv_data_242 : _GEN_3580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3582 = 8'hf3 == local_offset_3 ? phv_data_243 : _GEN_3581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3583 = 8'hf4 == local_offset_3 ? phv_data_244 : _GEN_3582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3584 = 8'hf5 == local_offset_3 ? phv_data_245 : _GEN_3583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3585 = 8'hf6 == local_offset_3 ? phv_data_246 : _GEN_3584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3586 = 8'hf7 == local_offset_3 ? phv_data_247 : _GEN_3585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3587 = 8'hf8 == local_offset_3 ? phv_data_248 : _GEN_3586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3588 = 8'hf9 == local_offset_3 ? phv_data_249 : _GEN_3587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3589 = 8'hfa == local_offset_3 ? phv_data_250 : _GEN_3588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3590 = 8'hfb == local_offset_3 ? phv_data_251 : _GEN_3589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3591 = 8'hfc == local_offset_3 ? phv_data_252 : _GEN_3590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3592 = 8'hfd == local_offset_3 ? phv_data_253 : _GEN_3591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3593 = 8'hfe == local_offset_3 ? phv_data_254 : _GEN_3592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3594 = 8'hff == local_offset_3 ? phv_data_255 : _GEN_3593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3596 = 8'h1 == _match_key_qbytes_3_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3597 = 8'h2 == _match_key_qbytes_3_T ? phv_data_2 : _GEN_3596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3598 = 8'h3 == _match_key_qbytes_3_T ? phv_data_3 : _GEN_3597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3599 = 8'h4 == _match_key_qbytes_3_T ? phv_data_4 : _GEN_3598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3600 = 8'h5 == _match_key_qbytes_3_T ? phv_data_5 : _GEN_3599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3601 = 8'h6 == _match_key_qbytes_3_T ? phv_data_6 : _GEN_3600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3602 = 8'h7 == _match_key_qbytes_3_T ? phv_data_7 : _GEN_3601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3603 = 8'h8 == _match_key_qbytes_3_T ? phv_data_8 : _GEN_3602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3604 = 8'h9 == _match_key_qbytes_3_T ? phv_data_9 : _GEN_3603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3605 = 8'ha == _match_key_qbytes_3_T ? phv_data_10 : _GEN_3604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3606 = 8'hb == _match_key_qbytes_3_T ? phv_data_11 : _GEN_3605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3607 = 8'hc == _match_key_qbytes_3_T ? phv_data_12 : _GEN_3606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3608 = 8'hd == _match_key_qbytes_3_T ? phv_data_13 : _GEN_3607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3609 = 8'he == _match_key_qbytes_3_T ? phv_data_14 : _GEN_3608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3610 = 8'hf == _match_key_qbytes_3_T ? phv_data_15 : _GEN_3609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3611 = 8'h10 == _match_key_qbytes_3_T ? phv_data_16 : _GEN_3610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3612 = 8'h11 == _match_key_qbytes_3_T ? phv_data_17 : _GEN_3611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3613 = 8'h12 == _match_key_qbytes_3_T ? phv_data_18 : _GEN_3612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3614 = 8'h13 == _match_key_qbytes_3_T ? phv_data_19 : _GEN_3613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3615 = 8'h14 == _match_key_qbytes_3_T ? phv_data_20 : _GEN_3614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3616 = 8'h15 == _match_key_qbytes_3_T ? phv_data_21 : _GEN_3615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3617 = 8'h16 == _match_key_qbytes_3_T ? phv_data_22 : _GEN_3616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3618 = 8'h17 == _match_key_qbytes_3_T ? phv_data_23 : _GEN_3617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3619 = 8'h18 == _match_key_qbytes_3_T ? phv_data_24 : _GEN_3618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3620 = 8'h19 == _match_key_qbytes_3_T ? phv_data_25 : _GEN_3619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3621 = 8'h1a == _match_key_qbytes_3_T ? phv_data_26 : _GEN_3620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3622 = 8'h1b == _match_key_qbytes_3_T ? phv_data_27 : _GEN_3621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3623 = 8'h1c == _match_key_qbytes_3_T ? phv_data_28 : _GEN_3622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3624 = 8'h1d == _match_key_qbytes_3_T ? phv_data_29 : _GEN_3623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3625 = 8'h1e == _match_key_qbytes_3_T ? phv_data_30 : _GEN_3624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3626 = 8'h1f == _match_key_qbytes_3_T ? phv_data_31 : _GEN_3625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3627 = 8'h20 == _match_key_qbytes_3_T ? phv_data_32 : _GEN_3626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3628 = 8'h21 == _match_key_qbytes_3_T ? phv_data_33 : _GEN_3627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3629 = 8'h22 == _match_key_qbytes_3_T ? phv_data_34 : _GEN_3628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3630 = 8'h23 == _match_key_qbytes_3_T ? phv_data_35 : _GEN_3629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3631 = 8'h24 == _match_key_qbytes_3_T ? phv_data_36 : _GEN_3630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3632 = 8'h25 == _match_key_qbytes_3_T ? phv_data_37 : _GEN_3631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3633 = 8'h26 == _match_key_qbytes_3_T ? phv_data_38 : _GEN_3632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3634 = 8'h27 == _match_key_qbytes_3_T ? phv_data_39 : _GEN_3633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3635 = 8'h28 == _match_key_qbytes_3_T ? phv_data_40 : _GEN_3634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3636 = 8'h29 == _match_key_qbytes_3_T ? phv_data_41 : _GEN_3635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3637 = 8'h2a == _match_key_qbytes_3_T ? phv_data_42 : _GEN_3636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3638 = 8'h2b == _match_key_qbytes_3_T ? phv_data_43 : _GEN_3637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3639 = 8'h2c == _match_key_qbytes_3_T ? phv_data_44 : _GEN_3638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3640 = 8'h2d == _match_key_qbytes_3_T ? phv_data_45 : _GEN_3639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3641 = 8'h2e == _match_key_qbytes_3_T ? phv_data_46 : _GEN_3640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3642 = 8'h2f == _match_key_qbytes_3_T ? phv_data_47 : _GEN_3641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3643 = 8'h30 == _match_key_qbytes_3_T ? phv_data_48 : _GEN_3642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3644 = 8'h31 == _match_key_qbytes_3_T ? phv_data_49 : _GEN_3643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3645 = 8'h32 == _match_key_qbytes_3_T ? phv_data_50 : _GEN_3644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3646 = 8'h33 == _match_key_qbytes_3_T ? phv_data_51 : _GEN_3645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3647 = 8'h34 == _match_key_qbytes_3_T ? phv_data_52 : _GEN_3646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3648 = 8'h35 == _match_key_qbytes_3_T ? phv_data_53 : _GEN_3647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3649 = 8'h36 == _match_key_qbytes_3_T ? phv_data_54 : _GEN_3648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3650 = 8'h37 == _match_key_qbytes_3_T ? phv_data_55 : _GEN_3649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3651 = 8'h38 == _match_key_qbytes_3_T ? phv_data_56 : _GEN_3650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3652 = 8'h39 == _match_key_qbytes_3_T ? phv_data_57 : _GEN_3651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3653 = 8'h3a == _match_key_qbytes_3_T ? phv_data_58 : _GEN_3652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3654 = 8'h3b == _match_key_qbytes_3_T ? phv_data_59 : _GEN_3653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3655 = 8'h3c == _match_key_qbytes_3_T ? phv_data_60 : _GEN_3654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3656 = 8'h3d == _match_key_qbytes_3_T ? phv_data_61 : _GEN_3655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3657 = 8'h3e == _match_key_qbytes_3_T ? phv_data_62 : _GEN_3656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3658 = 8'h3f == _match_key_qbytes_3_T ? phv_data_63 : _GEN_3657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3659 = 8'h40 == _match_key_qbytes_3_T ? phv_data_64 : _GEN_3658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3660 = 8'h41 == _match_key_qbytes_3_T ? phv_data_65 : _GEN_3659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3661 = 8'h42 == _match_key_qbytes_3_T ? phv_data_66 : _GEN_3660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3662 = 8'h43 == _match_key_qbytes_3_T ? phv_data_67 : _GEN_3661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3663 = 8'h44 == _match_key_qbytes_3_T ? phv_data_68 : _GEN_3662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3664 = 8'h45 == _match_key_qbytes_3_T ? phv_data_69 : _GEN_3663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3665 = 8'h46 == _match_key_qbytes_3_T ? phv_data_70 : _GEN_3664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3666 = 8'h47 == _match_key_qbytes_3_T ? phv_data_71 : _GEN_3665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3667 = 8'h48 == _match_key_qbytes_3_T ? phv_data_72 : _GEN_3666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3668 = 8'h49 == _match_key_qbytes_3_T ? phv_data_73 : _GEN_3667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3669 = 8'h4a == _match_key_qbytes_3_T ? phv_data_74 : _GEN_3668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3670 = 8'h4b == _match_key_qbytes_3_T ? phv_data_75 : _GEN_3669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3671 = 8'h4c == _match_key_qbytes_3_T ? phv_data_76 : _GEN_3670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3672 = 8'h4d == _match_key_qbytes_3_T ? phv_data_77 : _GEN_3671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3673 = 8'h4e == _match_key_qbytes_3_T ? phv_data_78 : _GEN_3672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3674 = 8'h4f == _match_key_qbytes_3_T ? phv_data_79 : _GEN_3673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3675 = 8'h50 == _match_key_qbytes_3_T ? phv_data_80 : _GEN_3674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3676 = 8'h51 == _match_key_qbytes_3_T ? phv_data_81 : _GEN_3675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3677 = 8'h52 == _match_key_qbytes_3_T ? phv_data_82 : _GEN_3676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3678 = 8'h53 == _match_key_qbytes_3_T ? phv_data_83 : _GEN_3677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3679 = 8'h54 == _match_key_qbytes_3_T ? phv_data_84 : _GEN_3678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3680 = 8'h55 == _match_key_qbytes_3_T ? phv_data_85 : _GEN_3679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3681 = 8'h56 == _match_key_qbytes_3_T ? phv_data_86 : _GEN_3680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3682 = 8'h57 == _match_key_qbytes_3_T ? phv_data_87 : _GEN_3681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3683 = 8'h58 == _match_key_qbytes_3_T ? phv_data_88 : _GEN_3682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3684 = 8'h59 == _match_key_qbytes_3_T ? phv_data_89 : _GEN_3683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3685 = 8'h5a == _match_key_qbytes_3_T ? phv_data_90 : _GEN_3684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3686 = 8'h5b == _match_key_qbytes_3_T ? phv_data_91 : _GEN_3685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3687 = 8'h5c == _match_key_qbytes_3_T ? phv_data_92 : _GEN_3686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3688 = 8'h5d == _match_key_qbytes_3_T ? phv_data_93 : _GEN_3687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3689 = 8'h5e == _match_key_qbytes_3_T ? phv_data_94 : _GEN_3688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3690 = 8'h5f == _match_key_qbytes_3_T ? phv_data_95 : _GEN_3689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3691 = 8'h60 == _match_key_qbytes_3_T ? phv_data_96 : _GEN_3690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3692 = 8'h61 == _match_key_qbytes_3_T ? phv_data_97 : _GEN_3691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3693 = 8'h62 == _match_key_qbytes_3_T ? phv_data_98 : _GEN_3692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3694 = 8'h63 == _match_key_qbytes_3_T ? phv_data_99 : _GEN_3693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3695 = 8'h64 == _match_key_qbytes_3_T ? phv_data_100 : _GEN_3694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3696 = 8'h65 == _match_key_qbytes_3_T ? phv_data_101 : _GEN_3695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3697 = 8'h66 == _match_key_qbytes_3_T ? phv_data_102 : _GEN_3696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3698 = 8'h67 == _match_key_qbytes_3_T ? phv_data_103 : _GEN_3697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3699 = 8'h68 == _match_key_qbytes_3_T ? phv_data_104 : _GEN_3698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3700 = 8'h69 == _match_key_qbytes_3_T ? phv_data_105 : _GEN_3699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3701 = 8'h6a == _match_key_qbytes_3_T ? phv_data_106 : _GEN_3700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3702 = 8'h6b == _match_key_qbytes_3_T ? phv_data_107 : _GEN_3701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3703 = 8'h6c == _match_key_qbytes_3_T ? phv_data_108 : _GEN_3702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3704 = 8'h6d == _match_key_qbytes_3_T ? phv_data_109 : _GEN_3703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3705 = 8'h6e == _match_key_qbytes_3_T ? phv_data_110 : _GEN_3704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3706 = 8'h6f == _match_key_qbytes_3_T ? phv_data_111 : _GEN_3705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3707 = 8'h70 == _match_key_qbytes_3_T ? phv_data_112 : _GEN_3706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3708 = 8'h71 == _match_key_qbytes_3_T ? phv_data_113 : _GEN_3707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3709 = 8'h72 == _match_key_qbytes_3_T ? phv_data_114 : _GEN_3708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3710 = 8'h73 == _match_key_qbytes_3_T ? phv_data_115 : _GEN_3709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3711 = 8'h74 == _match_key_qbytes_3_T ? phv_data_116 : _GEN_3710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3712 = 8'h75 == _match_key_qbytes_3_T ? phv_data_117 : _GEN_3711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3713 = 8'h76 == _match_key_qbytes_3_T ? phv_data_118 : _GEN_3712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3714 = 8'h77 == _match_key_qbytes_3_T ? phv_data_119 : _GEN_3713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3715 = 8'h78 == _match_key_qbytes_3_T ? phv_data_120 : _GEN_3714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3716 = 8'h79 == _match_key_qbytes_3_T ? phv_data_121 : _GEN_3715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3717 = 8'h7a == _match_key_qbytes_3_T ? phv_data_122 : _GEN_3716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3718 = 8'h7b == _match_key_qbytes_3_T ? phv_data_123 : _GEN_3717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3719 = 8'h7c == _match_key_qbytes_3_T ? phv_data_124 : _GEN_3718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3720 = 8'h7d == _match_key_qbytes_3_T ? phv_data_125 : _GEN_3719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3721 = 8'h7e == _match_key_qbytes_3_T ? phv_data_126 : _GEN_3720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3722 = 8'h7f == _match_key_qbytes_3_T ? phv_data_127 : _GEN_3721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3723 = 8'h80 == _match_key_qbytes_3_T ? phv_data_128 : _GEN_3722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3724 = 8'h81 == _match_key_qbytes_3_T ? phv_data_129 : _GEN_3723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3725 = 8'h82 == _match_key_qbytes_3_T ? phv_data_130 : _GEN_3724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3726 = 8'h83 == _match_key_qbytes_3_T ? phv_data_131 : _GEN_3725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3727 = 8'h84 == _match_key_qbytes_3_T ? phv_data_132 : _GEN_3726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3728 = 8'h85 == _match_key_qbytes_3_T ? phv_data_133 : _GEN_3727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3729 = 8'h86 == _match_key_qbytes_3_T ? phv_data_134 : _GEN_3728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3730 = 8'h87 == _match_key_qbytes_3_T ? phv_data_135 : _GEN_3729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3731 = 8'h88 == _match_key_qbytes_3_T ? phv_data_136 : _GEN_3730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3732 = 8'h89 == _match_key_qbytes_3_T ? phv_data_137 : _GEN_3731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3733 = 8'h8a == _match_key_qbytes_3_T ? phv_data_138 : _GEN_3732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3734 = 8'h8b == _match_key_qbytes_3_T ? phv_data_139 : _GEN_3733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3735 = 8'h8c == _match_key_qbytes_3_T ? phv_data_140 : _GEN_3734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3736 = 8'h8d == _match_key_qbytes_3_T ? phv_data_141 : _GEN_3735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3737 = 8'h8e == _match_key_qbytes_3_T ? phv_data_142 : _GEN_3736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3738 = 8'h8f == _match_key_qbytes_3_T ? phv_data_143 : _GEN_3737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3739 = 8'h90 == _match_key_qbytes_3_T ? phv_data_144 : _GEN_3738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3740 = 8'h91 == _match_key_qbytes_3_T ? phv_data_145 : _GEN_3739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3741 = 8'h92 == _match_key_qbytes_3_T ? phv_data_146 : _GEN_3740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3742 = 8'h93 == _match_key_qbytes_3_T ? phv_data_147 : _GEN_3741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3743 = 8'h94 == _match_key_qbytes_3_T ? phv_data_148 : _GEN_3742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3744 = 8'h95 == _match_key_qbytes_3_T ? phv_data_149 : _GEN_3743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3745 = 8'h96 == _match_key_qbytes_3_T ? phv_data_150 : _GEN_3744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3746 = 8'h97 == _match_key_qbytes_3_T ? phv_data_151 : _GEN_3745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3747 = 8'h98 == _match_key_qbytes_3_T ? phv_data_152 : _GEN_3746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3748 = 8'h99 == _match_key_qbytes_3_T ? phv_data_153 : _GEN_3747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3749 = 8'h9a == _match_key_qbytes_3_T ? phv_data_154 : _GEN_3748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3750 = 8'h9b == _match_key_qbytes_3_T ? phv_data_155 : _GEN_3749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3751 = 8'h9c == _match_key_qbytes_3_T ? phv_data_156 : _GEN_3750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3752 = 8'h9d == _match_key_qbytes_3_T ? phv_data_157 : _GEN_3751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3753 = 8'h9e == _match_key_qbytes_3_T ? phv_data_158 : _GEN_3752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3754 = 8'h9f == _match_key_qbytes_3_T ? phv_data_159 : _GEN_3753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3755 = 8'ha0 == _match_key_qbytes_3_T ? phv_data_160 : _GEN_3754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3756 = 8'ha1 == _match_key_qbytes_3_T ? phv_data_161 : _GEN_3755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3757 = 8'ha2 == _match_key_qbytes_3_T ? phv_data_162 : _GEN_3756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3758 = 8'ha3 == _match_key_qbytes_3_T ? phv_data_163 : _GEN_3757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3759 = 8'ha4 == _match_key_qbytes_3_T ? phv_data_164 : _GEN_3758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3760 = 8'ha5 == _match_key_qbytes_3_T ? phv_data_165 : _GEN_3759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3761 = 8'ha6 == _match_key_qbytes_3_T ? phv_data_166 : _GEN_3760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3762 = 8'ha7 == _match_key_qbytes_3_T ? phv_data_167 : _GEN_3761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3763 = 8'ha8 == _match_key_qbytes_3_T ? phv_data_168 : _GEN_3762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3764 = 8'ha9 == _match_key_qbytes_3_T ? phv_data_169 : _GEN_3763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3765 = 8'haa == _match_key_qbytes_3_T ? phv_data_170 : _GEN_3764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3766 = 8'hab == _match_key_qbytes_3_T ? phv_data_171 : _GEN_3765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3767 = 8'hac == _match_key_qbytes_3_T ? phv_data_172 : _GEN_3766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3768 = 8'had == _match_key_qbytes_3_T ? phv_data_173 : _GEN_3767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3769 = 8'hae == _match_key_qbytes_3_T ? phv_data_174 : _GEN_3768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3770 = 8'haf == _match_key_qbytes_3_T ? phv_data_175 : _GEN_3769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3771 = 8'hb0 == _match_key_qbytes_3_T ? phv_data_176 : _GEN_3770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3772 = 8'hb1 == _match_key_qbytes_3_T ? phv_data_177 : _GEN_3771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3773 = 8'hb2 == _match_key_qbytes_3_T ? phv_data_178 : _GEN_3772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3774 = 8'hb3 == _match_key_qbytes_3_T ? phv_data_179 : _GEN_3773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3775 = 8'hb4 == _match_key_qbytes_3_T ? phv_data_180 : _GEN_3774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3776 = 8'hb5 == _match_key_qbytes_3_T ? phv_data_181 : _GEN_3775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3777 = 8'hb6 == _match_key_qbytes_3_T ? phv_data_182 : _GEN_3776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3778 = 8'hb7 == _match_key_qbytes_3_T ? phv_data_183 : _GEN_3777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3779 = 8'hb8 == _match_key_qbytes_3_T ? phv_data_184 : _GEN_3778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3780 = 8'hb9 == _match_key_qbytes_3_T ? phv_data_185 : _GEN_3779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3781 = 8'hba == _match_key_qbytes_3_T ? phv_data_186 : _GEN_3780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3782 = 8'hbb == _match_key_qbytes_3_T ? phv_data_187 : _GEN_3781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3783 = 8'hbc == _match_key_qbytes_3_T ? phv_data_188 : _GEN_3782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3784 = 8'hbd == _match_key_qbytes_3_T ? phv_data_189 : _GEN_3783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3785 = 8'hbe == _match_key_qbytes_3_T ? phv_data_190 : _GEN_3784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3786 = 8'hbf == _match_key_qbytes_3_T ? phv_data_191 : _GEN_3785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3787 = 8'hc0 == _match_key_qbytes_3_T ? phv_data_192 : _GEN_3786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3788 = 8'hc1 == _match_key_qbytes_3_T ? phv_data_193 : _GEN_3787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3789 = 8'hc2 == _match_key_qbytes_3_T ? phv_data_194 : _GEN_3788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3790 = 8'hc3 == _match_key_qbytes_3_T ? phv_data_195 : _GEN_3789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3791 = 8'hc4 == _match_key_qbytes_3_T ? phv_data_196 : _GEN_3790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3792 = 8'hc5 == _match_key_qbytes_3_T ? phv_data_197 : _GEN_3791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3793 = 8'hc6 == _match_key_qbytes_3_T ? phv_data_198 : _GEN_3792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3794 = 8'hc7 == _match_key_qbytes_3_T ? phv_data_199 : _GEN_3793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3795 = 8'hc8 == _match_key_qbytes_3_T ? phv_data_200 : _GEN_3794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3796 = 8'hc9 == _match_key_qbytes_3_T ? phv_data_201 : _GEN_3795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3797 = 8'hca == _match_key_qbytes_3_T ? phv_data_202 : _GEN_3796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3798 = 8'hcb == _match_key_qbytes_3_T ? phv_data_203 : _GEN_3797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3799 = 8'hcc == _match_key_qbytes_3_T ? phv_data_204 : _GEN_3798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3800 = 8'hcd == _match_key_qbytes_3_T ? phv_data_205 : _GEN_3799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3801 = 8'hce == _match_key_qbytes_3_T ? phv_data_206 : _GEN_3800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3802 = 8'hcf == _match_key_qbytes_3_T ? phv_data_207 : _GEN_3801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3803 = 8'hd0 == _match_key_qbytes_3_T ? phv_data_208 : _GEN_3802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3804 = 8'hd1 == _match_key_qbytes_3_T ? phv_data_209 : _GEN_3803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3805 = 8'hd2 == _match_key_qbytes_3_T ? phv_data_210 : _GEN_3804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3806 = 8'hd3 == _match_key_qbytes_3_T ? phv_data_211 : _GEN_3805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3807 = 8'hd4 == _match_key_qbytes_3_T ? phv_data_212 : _GEN_3806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3808 = 8'hd5 == _match_key_qbytes_3_T ? phv_data_213 : _GEN_3807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3809 = 8'hd6 == _match_key_qbytes_3_T ? phv_data_214 : _GEN_3808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3810 = 8'hd7 == _match_key_qbytes_3_T ? phv_data_215 : _GEN_3809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3811 = 8'hd8 == _match_key_qbytes_3_T ? phv_data_216 : _GEN_3810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3812 = 8'hd9 == _match_key_qbytes_3_T ? phv_data_217 : _GEN_3811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3813 = 8'hda == _match_key_qbytes_3_T ? phv_data_218 : _GEN_3812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3814 = 8'hdb == _match_key_qbytes_3_T ? phv_data_219 : _GEN_3813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3815 = 8'hdc == _match_key_qbytes_3_T ? phv_data_220 : _GEN_3814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3816 = 8'hdd == _match_key_qbytes_3_T ? phv_data_221 : _GEN_3815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3817 = 8'hde == _match_key_qbytes_3_T ? phv_data_222 : _GEN_3816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3818 = 8'hdf == _match_key_qbytes_3_T ? phv_data_223 : _GEN_3817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3819 = 8'he0 == _match_key_qbytes_3_T ? phv_data_224 : _GEN_3818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3820 = 8'he1 == _match_key_qbytes_3_T ? phv_data_225 : _GEN_3819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3821 = 8'he2 == _match_key_qbytes_3_T ? phv_data_226 : _GEN_3820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3822 = 8'he3 == _match_key_qbytes_3_T ? phv_data_227 : _GEN_3821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3823 = 8'he4 == _match_key_qbytes_3_T ? phv_data_228 : _GEN_3822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3824 = 8'he5 == _match_key_qbytes_3_T ? phv_data_229 : _GEN_3823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3825 = 8'he6 == _match_key_qbytes_3_T ? phv_data_230 : _GEN_3824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3826 = 8'he7 == _match_key_qbytes_3_T ? phv_data_231 : _GEN_3825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3827 = 8'he8 == _match_key_qbytes_3_T ? phv_data_232 : _GEN_3826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3828 = 8'he9 == _match_key_qbytes_3_T ? phv_data_233 : _GEN_3827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3829 = 8'hea == _match_key_qbytes_3_T ? phv_data_234 : _GEN_3828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3830 = 8'heb == _match_key_qbytes_3_T ? phv_data_235 : _GEN_3829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3831 = 8'hec == _match_key_qbytes_3_T ? phv_data_236 : _GEN_3830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3832 = 8'hed == _match_key_qbytes_3_T ? phv_data_237 : _GEN_3831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3833 = 8'hee == _match_key_qbytes_3_T ? phv_data_238 : _GEN_3832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3834 = 8'hef == _match_key_qbytes_3_T ? phv_data_239 : _GEN_3833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3835 = 8'hf0 == _match_key_qbytes_3_T ? phv_data_240 : _GEN_3834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3836 = 8'hf1 == _match_key_qbytes_3_T ? phv_data_241 : _GEN_3835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3837 = 8'hf2 == _match_key_qbytes_3_T ? phv_data_242 : _GEN_3836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3838 = 8'hf3 == _match_key_qbytes_3_T ? phv_data_243 : _GEN_3837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3839 = 8'hf4 == _match_key_qbytes_3_T ? phv_data_244 : _GEN_3838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3840 = 8'hf5 == _match_key_qbytes_3_T ? phv_data_245 : _GEN_3839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3841 = 8'hf6 == _match_key_qbytes_3_T ? phv_data_246 : _GEN_3840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3842 = 8'hf7 == _match_key_qbytes_3_T ? phv_data_247 : _GEN_3841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3843 = 8'hf8 == _match_key_qbytes_3_T ? phv_data_248 : _GEN_3842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3844 = 8'hf9 == _match_key_qbytes_3_T ? phv_data_249 : _GEN_3843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3845 = 8'hfa == _match_key_qbytes_3_T ? phv_data_250 : _GEN_3844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3846 = 8'hfb == _match_key_qbytes_3_T ? phv_data_251 : _GEN_3845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3847 = 8'hfc == _match_key_qbytes_3_T ? phv_data_252 : _GEN_3846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3848 = 8'hfd == _match_key_qbytes_3_T ? phv_data_253 : _GEN_3847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3849 = 8'hfe == _match_key_qbytes_3_T ? phv_data_254 : _GEN_3848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3850 = 8'hff == _match_key_qbytes_3_T ? phv_data_255 : _GEN_3849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3852 = 8'h1 == _match_key_qbytes_3_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3853 = 8'h2 == _match_key_qbytes_3_T_1 ? phv_data_2 : _GEN_3852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3854 = 8'h3 == _match_key_qbytes_3_T_1 ? phv_data_3 : _GEN_3853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3855 = 8'h4 == _match_key_qbytes_3_T_1 ? phv_data_4 : _GEN_3854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3856 = 8'h5 == _match_key_qbytes_3_T_1 ? phv_data_5 : _GEN_3855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3857 = 8'h6 == _match_key_qbytes_3_T_1 ? phv_data_6 : _GEN_3856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3858 = 8'h7 == _match_key_qbytes_3_T_1 ? phv_data_7 : _GEN_3857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3859 = 8'h8 == _match_key_qbytes_3_T_1 ? phv_data_8 : _GEN_3858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3860 = 8'h9 == _match_key_qbytes_3_T_1 ? phv_data_9 : _GEN_3859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3861 = 8'ha == _match_key_qbytes_3_T_1 ? phv_data_10 : _GEN_3860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3862 = 8'hb == _match_key_qbytes_3_T_1 ? phv_data_11 : _GEN_3861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3863 = 8'hc == _match_key_qbytes_3_T_1 ? phv_data_12 : _GEN_3862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3864 = 8'hd == _match_key_qbytes_3_T_1 ? phv_data_13 : _GEN_3863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3865 = 8'he == _match_key_qbytes_3_T_1 ? phv_data_14 : _GEN_3864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3866 = 8'hf == _match_key_qbytes_3_T_1 ? phv_data_15 : _GEN_3865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3867 = 8'h10 == _match_key_qbytes_3_T_1 ? phv_data_16 : _GEN_3866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3868 = 8'h11 == _match_key_qbytes_3_T_1 ? phv_data_17 : _GEN_3867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3869 = 8'h12 == _match_key_qbytes_3_T_1 ? phv_data_18 : _GEN_3868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3870 = 8'h13 == _match_key_qbytes_3_T_1 ? phv_data_19 : _GEN_3869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3871 = 8'h14 == _match_key_qbytes_3_T_1 ? phv_data_20 : _GEN_3870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3872 = 8'h15 == _match_key_qbytes_3_T_1 ? phv_data_21 : _GEN_3871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3873 = 8'h16 == _match_key_qbytes_3_T_1 ? phv_data_22 : _GEN_3872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3874 = 8'h17 == _match_key_qbytes_3_T_1 ? phv_data_23 : _GEN_3873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3875 = 8'h18 == _match_key_qbytes_3_T_1 ? phv_data_24 : _GEN_3874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3876 = 8'h19 == _match_key_qbytes_3_T_1 ? phv_data_25 : _GEN_3875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3877 = 8'h1a == _match_key_qbytes_3_T_1 ? phv_data_26 : _GEN_3876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3878 = 8'h1b == _match_key_qbytes_3_T_1 ? phv_data_27 : _GEN_3877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3879 = 8'h1c == _match_key_qbytes_3_T_1 ? phv_data_28 : _GEN_3878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3880 = 8'h1d == _match_key_qbytes_3_T_1 ? phv_data_29 : _GEN_3879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3881 = 8'h1e == _match_key_qbytes_3_T_1 ? phv_data_30 : _GEN_3880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3882 = 8'h1f == _match_key_qbytes_3_T_1 ? phv_data_31 : _GEN_3881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3883 = 8'h20 == _match_key_qbytes_3_T_1 ? phv_data_32 : _GEN_3882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3884 = 8'h21 == _match_key_qbytes_3_T_1 ? phv_data_33 : _GEN_3883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3885 = 8'h22 == _match_key_qbytes_3_T_1 ? phv_data_34 : _GEN_3884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3886 = 8'h23 == _match_key_qbytes_3_T_1 ? phv_data_35 : _GEN_3885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3887 = 8'h24 == _match_key_qbytes_3_T_1 ? phv_data_36 : _GEN_3886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3888 = 8'h25 == _match_key_qbytes_3_T_1 ? phv_data_37 : _GEN_3887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3889 = 8'h26 == _match_key_qbytes_3_T_1 ? phv_data_38 : _GEN_3888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3890 = 8'h27 == _match_key_qbytes_3_T_1 ? phv_data_39 : _GEN_3889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3891 = 8'h28 == _match_key_qbytes_3_T_1 ? phv_data_40 : _GEN_3890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3892 = 8'h29 == _match_key_qbytes_3_T_1 ? phv_data_41 : _GEN_3891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3893 = 8'h2a == _match_key_qbytes_3_T_1 ? phv_data_42 : _GEN_3892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3894 = 8'h2b == _match_key_qbytes_3_T_1 ? phv_data_43 : _GEN_3893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3895 = 8'h2c == _match_key_qbytes_3_T_1 ? phv_data_44 : _GEN_3894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3896 = 8'h2d == _match_key_qbytes_3_T_1 ? phv_data_45 : _GEN_3895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3897 = 8'h2e == _match_key_qbytes_3_T_1 ? phv_data_46 : _GEN_3896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3898 = 8'h2f == _match_key_qbytes_3_T_1 ? phv_data_47 : _GEN_3897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3899 = 8'h30 == _match_key_qbytes_3_T_1 ? phv_data_48 : _GEN_3898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3900 = 8'h31 == _match_key_qbytes_3_T_1 ? phv_data_49 : _GEN_3899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3901 = 8'h32 == _match_key_qbytes_3_T_1 ? phv_data_50 : _GEN_3900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3902 = 8'h33 == _match_key_qbytes_3_T_1 ? phv_data_51 : _GEN_3901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3903 = 8'h34 == _match_key_qbytes_3_T_1 ? phv_data_52 : _GEN_3902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3904 = 8'h35 == _match_key_qbytes_3_T_1 ? phv_data_53 : _GEN_3903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3905 = 8'h36 == _match_key_qbytes_3_T_1 ? phv_data_54 : _GEN_3904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3906 = 8'h37 == _match_key_qbytes_3_T_1 ? phv_data_55 : _GEN_3905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3907 = 8'h38 == _match_key_qbytes_3_T_1 ? phv_data_56 : _GEN_3906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3908 = 8'h39 == _match_key_qbytes_3_T_1 ? phv_data_57 : _GEN_3907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3909 = 8'h3a == _match_key_qbytes_3_T_1 ? phv_data_58 : _GEN_3908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3910 = 8'h3b == _match_key_qbytes_3_T_1 ? phv_data_59 : _GEN_3909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3911 = 8'h3c == _match_key_qbytes_3_T_1 ? phv_data_60 : _GEN_3910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3912 = 8'h3d == _match_key_qbytes_3_T_1 ? phv_data_61 : _GEN_3911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3913 = 8'h3e == _match_key_qbytes_3_T_1 ? phv_data_62 : _GEN_3912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3914 = 8'h3f == _match_key_qbytes_3_T_1 ? phv_data_63 : _GEN_3913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3915 = 8'h40 == _match_key_qbytes_3_T_1 ? phv_data_64 : _GEN_3914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3916 = 8'h41 == _match_key_qbytes_3_T_1 ? phv_data_65 : _GEN_3915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3917 = 8'h42 == _match_key_qbytes_3_T_1 ? phv_data_66 : _GEN_3916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3918 = 8'h43 == _match_key_qbytes_3_T_1 ? phv_data_67 : _GEN_3917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3919 = 8'h44 == _match_key_qbytes_3_T_1 ? phv_data_68 : _GEN_3918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3920 = 8'h45 == _match_key_qbytes_3_T_1 ? phv_data_69 : _GEN_3919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3921 = 8'h46 == _match_key_qbytes_3_T_1 ? phv_data_70 : _GEN_3920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3922 = 8'h47 == _match_key_qbytes_3_T_1 ? phv_data_71 : _GEN_3921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3923 = 8'h48 == _match_key_qbytes_3_T_1 ? phv_data_72 : _GEN_3922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3924 = 8'h49 == _match_key_qbytes_3_T_1 ? phv_data_73 : _GEN_3923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3925 = 8'h4a == _match_key_qbytes_3_T_1 ? phv_data_74 : _GEN_3924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3926 = 8'h4b == _match_key_qbytes_3_T_1 ? phv_data_75 : _GEN_3925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3927 = 8'h4c == _match_key_qbytes_3_T_1 ? phv_data_76 : _GEN_3926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3928 = 8'h4d == _match_key_qbytes_3_T_1 ? phv_data_77 : _GEN_3927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3929 = 8'h4e == _match_key_qbytes_3_T_1 ? phv_data_78 : _GEN_3928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3930 = 8'h4f == _match_key_qbytes_3_T_1 ? phv_data_79 : _GEN_3929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3931 = 8'h50 == _match_key_qbytes_3_T_1 ? phv_data_80 : _GEN_3930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3932 = 8'h51 == _match_key_qbytes_3_T_1 ? phv_data_81 : _GEN_3931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3933 = 8'h52 == _match_key_qbytes_3_T_1 ? phv_data_82 : _GEN_3932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3934 = 8'h53 == _match_key_qbytes_3_T_1 ? phv_data_83 : _GEN_3933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3935 = 8'h54 == _match_key_qbytes_3_T_1 ? phv_data_84 : _GEN_3934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3936 = 8'h55 == _match_key_qbytes_3_T_1 ? phv_data_85 : _GEN_3935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3937 = 8'h56 == _match_key_qbytes_3_T_1 ? phv_data_86 : _GEN_3936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3938 = 8'h57 == _match_key_qbytes_3_T_1 ? phv_data_87 : _GEN_3937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3939 = 8'h58 == _match_key_qbytes_3_T_1 ? phv_data_88 : _GEN_3938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3940 = 8'h59 == _match_key_qbytes_3_T_1 ? phv_data_89 : _GEN_3939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3941 = 8'h5a == _match_key_qbytes_3_T_1 ? phv_data_90 : _GEN_3940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3942 = 8'h5b == _match_key_qbytes_3_T_1 ? phv_data_91 : _GEN_3941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3943 = 8'h5c == _match_key_qbytes_3_T_1 ? phv_data_92 : _GEN_3942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3944 = 8'h5d == _match_key_qbytes_3_T_1 ? phv_data_93 : _GEN_3943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3945 = 8'h5e == _match_key_qbytes_3_T_1 ? phv_data_94 : _GEN_3944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3946 = 8'h5f == _match_key_qbytes_3_T_1 ? phv_data_95 : _GEN_3945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3947 = 8'h60 == _match_key_qbytes_3_T_1 ? phv_data_96 : _GEN_3946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3948 = 8'h61 == _match_key_qbytes_3_T_1 ? phv_data_97 : _GEN_3947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3949 = 8'h62 == _match_key_qbytes_3_T_1 ? phv_data_98 : _GEN_3948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3950 = 8'h63 == _match_key_qbytes_3_T_1 ? phv_data_99 : _GEN_3949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3951 = 8'h64 == _match_key_qbytes_3_T_1 ? phv_data_100 : _GEN_3950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3952 = 8'h65 == _match_key_qbytes_3_T_1 ? phv_data_101 : _GEN_3951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3953 = 8'h66 == _match_key_qbytes_3_T_1 ? phv_data_102 : _GEN_3952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3954 = 8'h67 == _match_key_qbytes_3_T_1 ? phv_data_103 : _GEN_3953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3955 = 8'h68 == _match_key_qbytes_3_T_1 ? phv_data_104 : _GEN_3954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3956 = 8'h69 == _match_key_qbytes_3_T_1 ? phv_data_105 : _GEN_3955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3957 = 8'h6a == _match_key_qbytes_3_T_1 ? phv_data_106 : _GEN_3956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3958 = 8'h6b == _match_key_qbytes_3_T_1 ? phv_data_107 : _GEN_3957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3959 = 8'h6c == _match_key_qbytes_3_T_1 ? phv_data_108 : _GEN_3958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3960 = 8'h6d == _match_key_qbytes_3_T_1 ? phv_data_109 : _GEN_3959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3961 = 8'h6e == _match_key_qbytes_3_T_1 ? phv_data_110 : _GEN_3960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3962 = 8'h6f == _match_key_qbytes_3_T_1 ? phv_data_111 : _GEN_3961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3963 = 8'h70 == _match_key_qbytes_3_T_1 ? phv_data_112 : _GEN_3962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3964 = 8'h71 == _match_key_qbytes_3_T_1 ? phv_data_113 : _GEN_3963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3965 = 8'h72 == _match_key_qbytes_3_T_1 ? phv_data_114 : _GEN_3964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3966 = 8'h73 == _match_key_qbytes_3_T_1 ? phv_data_115 : _GEN_3965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3967 = 8'h74 == _match_key_qbytes_3_T_1 ? phv_data_116 : _GEN_3966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3968 = 8'h75 == _match_key_qbytes_3_T_1 ? phv_data_117 : _GEN_3967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3969 = 8'h76 == _match_key_qbytes_3_T_1 ? phv_data_118 : _GEN_3968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3970 = 8'h77 == _match_key_qbytes_3_T_1 ? phv_data_119 : _GEN_3969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3971 = 8'h78 == _match_key_qbytes_3_T_1 ? phv_data_120 : _GEN_3970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3972 = 8'h79 == _match_key_qbytes_3_T_1 ? phv_data_121 : _GEN_3971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3973 = 8'h7a == _match_key_qbytes_3_T_1 ? phv_data_122 : _GEN_3972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3974 = 8'h7b == _match_key_qbytes_3_T_1 ? phv_data_123 : _GEN_3973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3975 = 8'h7c == _match_key_qbytes_3_T_1 ? phv_data_124 : _GEN_3974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3976 = 8'h7d == _match_key_qbytes_3_T_1 ? phv_data_125 : _GEN_3975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3977 = 8'h7e == _match_key_qbytes_3_T_1 ? phv_data_126 : _GEN_3976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3978 = 8'h7f == _match_key_qbytes_3_T_1 ? phv_data_127 : _GEN_3977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3979 = 8'h80 == _match_key_qbytes_3_T_1 ? phv_data_128 : _GEN_3978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3980 = 8'h81 == _match_key_qbytes_3_T_1 ? phv_data_129 : _GEN_3979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3981 = 8'h82 == _match_key_qbytes_3_T_1 ? phv_data_130 : _GEN_3980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3982 = 8'h83 == _match_key_qbytes_3_T_1 ? phv_data_131 : _GEN_3981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3983 = 8'h84 == _match_key_qbytes_3_T_1 ? phv_data_132 : _GEN_3982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3984 = 8'h85 == _match_key_qbytes_3_T_1 ? phv_data_133 : _GEN_3983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3985 = 8'h86 == _match_key_qbytes_3_T_1 ? phv_data_134 : _GEN_3984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3986 = 8'h87 == _match_key_qbytes_3_T_1 ? phv_data_135 : _GEN_3985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3987 = 8'h88 == _match_key_qbytes_3_T_1 ? phv_data_136 : _GEN_3986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3988 = 8'h89 == _match_key_qbytes_3_T_1 ? phv_data_137 : _GEN_3987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3989 = 8'h8a == _match_key_qbytes_3_T_1 ? phv_data_138 : _GEN_3988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3990 = 8'h8b == _match_key_qbytes_3_T_1 ? phv_data_139 : _GEN_3989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3991 = 8'h8c == _match_key_qbytes_3_T_1 ? phv_data_140 : _GEN_3990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3992 = 8'h8d == _match_key_qbytes_3_T_1 ? phv_data_141 : _GEN_3991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3993 = 8'h8e == _match_key_qbytes_3_T_1 ? phv_data_142 : _GEN_3992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3994 = 8'h8f == _match_key_qbytes_3_T_1 ? phv_data_143 : _GEN_3993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3995 = 8'h90 == _match_key_qbytes_3_T_1 ? phv_data_144 : _GEN_3994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3996 = 8'h91 == _match_key_qbytes_3_T_1 ? phv_data_145 : _GEN_3995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3997 = 8'h92 == _match_key_qbytes_3_T_1 ? phv_data_146 : _GEN_3996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3998 = 8'h93 == _match_key_qbytes_3_T_1 ? phv_data_147 : _GEN_3997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3999 = 8'h94 == _match_key_qbytes_3_T_1 ? phv_data_148 : _GEN_3998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4000 = 8'h95 == _match_key_qbytes_3_T_1 ? phv_data_149 : _GEN_3999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4001 = 8'h96 == _match_key_qbytes_3_T_1 ? phv_data_150 : _GEN_4000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4002 = 8'h97 == _match_key_qbytes_3_T_1 ? phv_data_151 : _GEN_4001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4003 = 8'h98 == _match_key_qbytes_3_T_1 ? phv_data_152 : _GEN_4002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4004 = 8'h99 == _match_key_qbytes_3_T_1 ? phv_data_153 : _GEN_4003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4005 = 8'h9a == _match_key_qbytes_3_T_1 ? phv_data_154 : _GEN_4004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4006 = 8'h9b == _match_key_qbytes_3_T_1 ? phv_data_155 : _GEN_4005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4007 = 8'h9c == _match_key_qbytes_3_T_1 ? phv_data_156 : _GEN_4006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4008 = 8'h9d == _match_key_qbytes_3_T_1 ? phv_data_157 : _GEN_4007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4009 = 8'h9e == _match_key_qbytes_3_T_1 ? phv_data_158 : _GEN_4008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4010 = 8'h9f == _match_key_qbytes_3_T_1 ? phv_data_159 : _GEN_4009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4011 = 8'ha0 == _match_key_qbytes_3_T_1 ? phv_data_160 : _GEN_4010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4012 = 8'ha1 == _match_key_qbytes_3_T_1 ? phv_data_161 : _GEN_4011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4013 = 8'ha2 == _match_key_qbytes_3_T_1 ? phv_data_162 : _GEN_4012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4014 = 8'ha3 == _match_key_qbytes_3_T_1 ? phv_data_163 : _GEN_4013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4015 = 8'ha4 == _match_key_qbytes_3_T_1 ? phv_data_164 : _GEN_4014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4016 = 8'ha5 == _match_key_qbytes_3_T_1 ? phv_data_165 : _GEN_4015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4017 = 8'ha6 == _match_key_qbytes_3_T_1 ? phv_data_166 : _GEN_4016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4018 = 8'ha7 == _match_key_qbytes_3_T_1 ? phv_data_167 : _GEN_4017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4019 = 8'ha8 == _match_key_qbytes_3_T_1 ? phv_data_168 : _GEN_4018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4020 = 8'ha9 == _match_key_qbytes_3_T_1 ? phv_data_169 : _GEN_4019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4021 = 8'haa == _match_key_qbytes_3_T_1 ? phv_data_170 : _GEN_4020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4022 = 8'hab == _match_key_qbytes_3_T_1 ? phv_data_171 : _GEN_4021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4023 = 8'hac == _match_key_qbytes_3_T_1 ? phv_data_172 : _GEN_4022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4024 = 8'had == _match_key_qbytes_3_T_1 ? phv_data_173 : _GEN_4023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4025 = 8'hae == _match_key_qbytes_3_T_1 ? phv_data_174 : _GEN_4024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4026 = 8'haf == _match_key_qbytes_3_T_1 ? phv_data_175 : _GEN_4025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4027 = 8'hb0 == _match_key_qbytes_3_T_1 ? phv_data_176 : _GEN_4026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4028 = 8'hb1 == _match_key_qbytes_3_T_1 ? phv_data_177 : _GEN_4027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4029 = 8'hb2 == _match_key_qbytes_3_T_1 ? phv_data_178 : _GEN_4028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4030 = 8'hb3 == _match_key_qbytes_3_T_1 ? phv_data_179 : _GEN_4029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4031 = 8'hb4 == _match_key_qbytes_3_T_1 ? phv_data_180 : _GEN_4030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4032 = 8'hb5 == _match_key_qbytes_3_T_1 ? phv_data_181 : _GEN_4031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4033 = 8'hb6 == _match_key_qbytes_3_T_1 ? phv_data_182 : _GEN_4032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4034 = 8'hb7 == _match_key_qbytes_3_T_1 ? phv_data_183 : _GEN_4033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4035 = 8'hb8 == _match_key_qbytes_3_T_1 ? phv_data_184 : _GEN_4034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4036 = 8'hb9 == _match_key_qbytes_3_T_1 ? phv_data_185 : _GEN_4035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4037 = 8'hba == _match_key_qbytes_3_T_1 ? phv_data_186 : _GEN_4036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4038 = 8'hbb == _match_key_qbytes_3_T_1 ? phv_data_187 : _GEN_4037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4039 = 8'hbc == _match_key_qbytes_3_T_1 ? phv_data_188 : _GEN_4038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4040 = 8'hbd == _match_key_qbytes_3_T_1 ? phv_data_189 : _GEN_4039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4041 = 8'hbe == _match_key_qbytes_3_T_1 ? phv_data_190 : _GEN_4040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4042 = 8'hbf == _match_key_qbytes_3_T_1 ? phv_data_191 : _GEN_4041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4043 = 8'hc0 == _match_key_qbytes_3_T_1 ? phv_data_192 : _GEN_4042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4044 = 8'hc1 == _match_key_qbytes_3_T_1 ? phv_data_193 : _GEN_4043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4045 = 8'hc2 == _match_key_qbytes_3_T_1 ? phv_data_194 : _GEN_4044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4046 = 8'hc3 == _match_key_qbytes_3_T_1 ? phv_data_195 : _GEN_4045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4047 = 8'hc4 == _match_key_qbytes_3_T_1 ? phv_data_196 : _GEN_4046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4048 = 8'hc5 == _match_key_qbytes_3_T_1 ? phv_data_197 : _GEN_4047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4049 = 8'hc6 == _match_key_qbytes_3_T_1 ? phv_data_198 : _GEN_4048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4050 = 8'hc7 == _match_key_qbytes_3_T_1 ? phv_data_199 : _GEN_4049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4051 = 8'hc8 == _match_key_qbytes_3_T_1 ? phv_data_200 : _GEN_4050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4052 = 8'hc9 == _match_key_qbytes_3_T_1 ? phv_data_201 : _GEN_4051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4053 = 8'hca == _match_key_qbytes_3_T_1 ? phv_data_202 : _GEN_4052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4054 = 8'hcb == _match_key_qbytes_3_T_1 ? phv_data_203 : _GEN_4053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4055 = 8'hcc == _match_key_qbytes_3_T_1 ? phv_data_204 : _GEN_4054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4056 = 8'hcd == _match_key_qbytes_3_T_1 ? phv_data_205 : _GEN_4055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4057 = 8'hce == _match_key_qbytes_3_T_1 ? phv_data_206 : _GEN_4056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4058 = 8'hcf == _match_key_qbytes_3_T_1 ? phv_data_207 : _GEN_4057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4059 = 8'hd0 == _match_key_qbytes_3_T_1 ? phv_data_208 : _GEN_4058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4060 = 8'hd1 == _match_key_qbytes_3_T_1 ? phv_data_209 : _GEN_4059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4061 = 8'hd2 == _match_key_qbytes_3_T_1 ? phv_data_210 : _GEN_4060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4062 = 8'hd3 == _match_key_qbytes_3_T_1 ? phv_data_211 : _GEN_4061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4063 = 8'hd4 == _match_key_qbytes_3_T_1 ? phv_data_212 : _GEN_4062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4064 = 8'hd5 == _match_key_qbytes_3_T_1 ? phv_data_213 : _GEN_4063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4065 = 8'hd6 == _match_key_qbytes_3_T_1 ? phv_data_214 : _GEN_4064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4066 = 8'hd7 == _match_key_qbytes_3_T_1 ? phv_data_215 : _GEN_4065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4067 = 8'hd8 == _match_key_qbytes_3_T_1 ? phv_data_216 : _GEN_4066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4068 = 8'hd9 == _match_key_qbytes_3_T_1 ? phv_data_217 : _GEN_4067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4069 = 8'hda == _match_key_qbytes_3_T_1 ? phv_data_218 : _GEN_4068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4070 = 8'hdb == _match_key_qbytes_3_T_1 ? phv_data_219 : _GEN_4069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4071 = 8'hdc == _match_key_qbytes_3_T_1 ? phv_data_220 : _GEN_4070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4072 = 8'hdd == _match_key_qbytes_3_T_1 ? phv_data_221 : _GEN_4071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4073 = 8'hde == _match_key_qbytes_3_T_1 ? phv_data_222 : _GEN_4072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4074 = 8'hdf == _match_key_qbytes_3_T_1 ? phv_data_223 : _GEN_4073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4075 = 8'he0 == _match_key_qbytes_3_T_1 ? phv_data_224 : _GEN_4074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4076 = 8'he1 == _match_key_qbytes_3_T_1 ? phv_data_225 : _GEN_4075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4077 = 8'he2 == _match_key_qbytes_3_T_1 ? phv_data_226 : _GEN_4076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4078 = 8'he3 == _match_key_qbytes_3_T_1 ? phv_data_227 : _GEN_4077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4079 = 8'he4 == _match_key_qbytes_3_T_1 ? phv_data_228 : _GEN_4078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4080 = 8'he5 == _match_key_qbytes_3_T_1 ? phv_data_229 : _GEN_4079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4081 = 8'he6 == _match_key_qbytes_3_T_1 ? phv_data_230 : _GEN_4080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4082 = 8'he7 == _match_key_qbytes_3_T_1 ? phv_data_231 : _GEN_4081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4083 = 8'he8 == _match_key_qbytes_3_T_1 ? phv_data_232 : _GEN_4082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4084 = 8'he9 == _match_key_qbytes_3_T_1 ? phv_data_233 : _GEN_4083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4085 = 8'hea == _match_key_qbytes_3_T_1 ? phv_data_234 : _GEN_4084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4086 = 8'heb == _match_key_qbytes_3_T_1 ? phv_data_235 : _GEN_4085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4087 = 8'hec == _match_key_qbytes_3_T_1 ? phv_data_236 : _GEN_4086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4088 = 8'hed == _match_key_qbytes_3_T_1 ? phv_data_237 : _GEN_4087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4089 = 8'hee == _match_key_qbytes_3_T_1 ? phv_data_238 : _GEN_4088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4090 = 8'hef == _match_key_qbytes_3_T_1 ? phv_data_239 : _GEN_4089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4091 = 8'hf0 == _match_key_qbytes_3_T_1 ? phv_data_240 : _GEN_4090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4092 = 8'hf1 == _match_key_qbytes_3_T_1 ? phv_data_241 : _GEN_4091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4093 = 8'hf2 == _match_key_qbytes_3_T_1 ? phv_data_242 : _GEN_4092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4094 = 8'hf3 == _match_key_qbytes_3_T_1 ? phv_data_243 : _GEN_4093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4095 = 8'hf4 == _match_key_qbytes_3_T_1 ? phv_data_244 : _GEN_4094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4096 = 8'hf5 == _match_key_qbytes_3_T_1 ? phv_data_245 : _GEN_4095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4097 = 8'hf6 == _match_key_qbytes_3_T_1 ? phv_data_246 : _GEN_4096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4098 = 8'hf7 == _match_key_qbytes_3_T_1 ? phv_data_247 : _GEN_4097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4099 = 8'hf8 == _match_key_qbytes_3_T_1 ? phv_data_248 : _GEN_4098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4100 = 8'hf9 == _match_key_qbytes_3_T_1 ? phv_data_249 : _GEN_4099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4101 = 8'hfa == _match_key_qbytes_3_T_1 ? phv_data_250 : _GEN_4100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4102 = 8'hfb == _match_key_qbytes_3_T_1 ? phv_data_251 : _GEN_4101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4103 = 8'hfc == _match_key_qbytes_3_T_1 ? phv_data_252 : _GEN_4102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4104 = 8'hfd == _match_key_qbytes_3_T_1 ? phv_data_253 : _GEN_4103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4105 = 8'hfe == _match_key_qbytes_3_T_1 ? phv_data_254 : _GEN_4104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4106 = 8'hff == _match_key_qbytes_3_T_1 ? phv_data_255 : _GEN_4105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_3_T_3 = {_GEN_3850,_GEN_4106,_GEN_3338,_GEN_3594}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_3 = local_offset_3 < end_offset ? _match_key_qbytes_3_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_4 = 8'h10 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_4_hi = local_offset_4[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_4_T = {match_key_qbytes_4_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_4_T_1 = {match_key_qbytes_4_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_4_T_2 = {match_key_qbytes_4_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_4109 = 8'h1 == _match_key_qbytes_4_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4110 = 8'h2 == _match_key_qbytes_4_T_2 ? phv_data_2 : _GEN_4109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4111 = 8'h3 == _match_key_qbytes_4_T_2 ? phv_data_3 : _GEN_4110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4112 = 8'h4 == _match_key_qbytes_4_T_2 ? phv_data_4 : _GEN_4111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4113 = 8'h5 == _match_key_qbytes_4_T_2 ? phv_data_5 : _GEN_4112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4114 = 8'h6 == _match_key_qbytes_4_T_2 ? phv_data_6 : _GEN_4113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4115 = 8'h7 == _match_key_qbytes_4_T_2 ? phv_data_7 : _GEN_4114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4116 = 8'h8 == _match_key_qbytes_4_T_2 ? phv_data_8 : _GEN_4115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4117 = 8'h9 == _match_key_qbytes_4_T_2 ? phv_data_9 : _GEN_4116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4118 = 8'ha == _match_key_qbytes_4_T_2 ? phv_data_10 : _GEN_4117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4119 = 8'hb == _match_key_qbytes_4_T_2 ? phv_data_11 : _GEN_4118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4120 = 8'hc == _match_key_qbytes_4_T_2 ? phv_data_12 : _GEN_4119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4121 = 8'hd == _match_key_qbytes_4_T_2 ? phv_data_13 : _GEN_4120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4122 = 8'he == _match_key_qbytes_4_T_2 ? phv_data_14 : _GEN_4121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4123 = 8'hf == _match_key_qbytes_4_T_2 ? phv_data_15 : _GEN_4122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4124 = 8'h10 == _match_key_qbytes_4_T_2 ? phv_data_16 : _GEN_4123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4125 = 8'h11 == _match_key_qbytes_4_T_2 ? phv_data_17 : _GEN_4124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4126 = 8'h12 == _match_key_qbytes_4_T_2 ? phv_data_18 : _GEN_4125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4127 = 8'h13 == _match_key_qbytes_4_T_2 ? phv_data_19 : _GEN_4126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4128 = 8'h14 == _match_key_qbytes_4_T_2 ? phv_data_20 : _GEN_4127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4129 = 8'h15 == _match_key_qbytes_4_T_2 ? phv_data_21 : _GEN_4128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4130 = 8'h16 == _match_key_qbytes_4_T_2 ? phv_data_22 : _GEN_4129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4131 = 8'h17 == _match_key_qbytes_4_T_2 ? phv_data_23 : _GEN_4130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4132 = 8'h18 == _match_key_qbytes_4_T_2 ? phv_data_24 : _GEN_4131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4133 = 8'h19 == _match_key_qbytes_4_T_2 ? phv_data_25 : _GEN_4132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4134 = 8'h1a == _match_key_qbytes_4_T_2 ? phv_data_26 : _GEN_4133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4135 = 8'h1b == _match_key_qbytes_4_T_2 ? phv_data_27 : _GEN_4134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4136 = 8'h1c == _match_key_qbytes_4_T_2 ? phv_data_28 : _GEN_4135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4137 = 8'h1d == _match_key_qbytes_4_T_2 ? phv_data_29 : _GEN_4136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4138 = 8'h1e == _match_key_qbytes_4_T_2 ? phv_data_30 : _GEN_4137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4139 = 8'h1f == _match_key_qbytes_4_T_2 ? phv_data_31 : _GEN_4138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4140 = 8'h20 == _match_key_qbytes_4_T_2 ? phv_data_32 : _GEN_4139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4141 = 8'h21 == _match_key_qbytes_4_T_2 ? phv_data_33 : _GEN_4140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4142 = 8'h22 == _match_key_qbytes_4_T_2 ? phv_data_34 : _GEN_4141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4143 = 8'h23 == _match_key_qbytes_4_T_2 ? phv_data_35 : _GEN_4142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4144 = 8'h24 == _match_key_qbytes_4_T_2 ? phv_data_36 : _GEN_4143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4145 = 8'h25 == _match_key_qbytes_4_T_2 ? phv_data_37 : _GEN_4144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4146 = 8'h26 == _match_key_qbytes_4_T_2 ? phv_data_38 : _GEN_4145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4147 = 8'h27 == _match_key_qbytes_4_T_2 ? phv_data_39 : _GEN_4146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4148 = 8'h28 == _match_key_qbytes_4_T_2 ? phv_data_40 : _GEN_4147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4149 = 8'h29 == _match_key_qbytes_4_T_2 ? phv_data_41 : _GEN_4148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4150 = 8'h2a == _match_key_qbytes_4_T_2 ? phv_data_42 : _GEN_4149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4151 = 8'h2b == _match_key_qbytes_4_T_2 ? phv_data_43 : _GEN_4150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4152 = 8'h2c == _match_key_qbytes_4_T_2 ? phv_data_44 : _GEN_4151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4153 = 8'h2d == _match_key_qbytes_4_T_2 ? phv_data_45 : _GEN_4152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4154 = 8'h2e == _match_key_qbytes_4_T_2 ? phv_data_46 : _GEN_4153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4155 = 8'h2f == _match_key_qbytes_4_T_2 ? phv_data_47 : _GEN_4154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4156 = 8'h30 == _match_key_qbytes_4_T_2 ? phv_data_48 : _GEN_4155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4157 = 8'h31 == _match_key_qbytes_4_T_2 ? phv_data_49 : _GEN_4156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4158 = 8'h32 == _match_key_qbytes_4_T_2 ? phv_data_50 : _GEN_4157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4159 = 8'h33 == _match_key_qbytes_4_T_2 ? phv_data_51 : _GEN_4158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4160 = 8'h34 == _match_key_qbytes_4_T_2 ? phv_data_52 : _GEN_4159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4161 = 8'h35 == _match_key_qbytes_4_T_2 ? phv_data_53 : _GEN_4160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4162 = 8'h36 == _match_key_qbytes_4_T_2 ? phv_data_54 : _GEN_4161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4163 = 8'h37 == _match_key_qbytes_4_T_2 ? phv_data_55 : _GEN_4162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4164 = 8'h38 == _match_key_qbytes_4_T_2 ? phv_data_56 : _GEN_4163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4165 = 8'h39 == _match_key_qbytes_4_T_2 ? phv_data_57 : _GEN_4164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4166 = 8'h3a == _match_key_qbytes_4_T_2 ? phv_data_58 : _GEN_4165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4167 = 8'h3b == _match_key_qbytes_4_T_2 ? phv_data_59 : _GEN_4166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4168 = 8'h3c == _match_key_qbytes_4_T_2 ? phv_data_60 : _GEN_4167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4169 = 8'h3d == _match_key_qbytes_4_T_2 ? phv_data_61 : _GEN_4168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4170 = 8'h3e == _match_key_qbytes_4_T_2 ? phv_data_62 : _GEN_4169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4171 = 8'h3f == _match_key_qbytes_4_T_2 ? phv_data_63 : _GEN_4170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4172 = 8'h40 == _match_key_qbytes_4_T_2 ? phv_data_64 : _GEN_4171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4173 = 8'h41 == _match_key_qbytes_4_T_2 ? phv_data_65 : _GEN_4172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4174 = 8'h42 == _match_key_qbytes_4_T_2 ? phv_data_66 : _GEN_4173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4175 = 8'h43 == _match_key_qbytes_4_T_2 ? phv_data_67 : _GEN_4174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4176 = 8'h44 == _match_key_qbytes_4_T_2 ? phv_data_68 : _GEN_4175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4177 = 8'h45 == _match_key_qbytes_4_T_2 ? phv_data_69 : _GEN_4176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4178 = 8'h46 == _match_key_qbytes_4_T_2 ? phv_data_70 : _GEN_4177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4179 = 8'h47 == _match_key_qbytes_4_T_2 ? phv_data_71 : _GEN_4178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4180 = 8'h48 == _match_key_qbytes_4_T_2 ? phv_data_72 : _GEN_4179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4181 = 8'h49 == _match_key_qbytes_4_T_2 ? phv_data_73 : _GEN_4180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4182 = 8'h4a == _match_key_qbytes_4_T_2 ? phv_data_74 : _GEN_4181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4183 = 8'h4b == _match_key_qbytes_4_T_2 ? phv_data_75 : _GEN_4182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4184 = 8'h4c == _match_key_qbytes_4_T_2 ? phv_data_76 : _GEN_4183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4185 = 8'h4d == _match_key_qbytes_4_T_2 ? phv_data_77 : _GEN_4184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4186 = 8'h4e == _match_key_qbytes_4_T_2 ? phv_data_78 : _GEN_4185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4187 = 8'h4f == _match_key_qbytes_4_T_2 ? phv_data_79 : _GEN_4186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4188 = 8'h50 == _match_key_qbytes_4_T_2 ? phv_data_80 : _GEN_4187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4189 = 8'h51 == _match_key_qbytes_4_T_2 ? phv_data_81 : _GEN_4188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4190 = 8'h52 == _match_key_qbytes_4_T_2 ? phv_data_82 : _GEN_4189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4191 = 8'h53 == _match_key_qbytes_4_T_2 ? phv_data_83 : _GEN_4190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4192 = 8'h54 == _match_key_qbytes_4_T_2 ? phv_data_84 : _GEN_4191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4193 = 8'h55 == _match_key_qbytes_4_T_2 ? phv_data_85 : _GEN_4192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4194 = 8'h56 == _match_key_qbytes_4_T_2 ? phv_data_86 : _GEN_4193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4195 = 8'h57 == _match_key_qbytes_4_T_2 ? phv_data_87 : _GEN_4194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4196 = 8'h58 == _match_key_qbytes_4_T_2 ? phv_data_88 : _GEN_4195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4197 = 8'h59 == _match_key_qbytes_4_T_2 ? phv_data_89 : _GEN_4196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4198 = 8'h5a == _match_key_qbytes_4_T_2 ? phv_data_90 : _GEN_4197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4199 = 8'h5b == _match_key_qbytes_4_T_2 ? phv_data_91 : _GEN_4198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4200 = 8'h5c == _match_key_qbytes_4_T_2 ? phv_data_92 : _GEN_4199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4201 = 8'h5d == _match_key_qbytes_4_T_2 ? phv_data_93 : _GEN_4200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4202 = 8'h5e == _match_key_qbytes_4_T_2 ? phv_data_94 : _GEN_4201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4203 = 8'h5f == _match_key_qbytes_4_T_2 ? phv_data_95 : _GEN_4202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4204 = 8'h60 == _match_key_qbytes_4_T_2 ? phv_data_96 : _GEN_4203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4205 = 8'h61 == _match_key_qbytes_4_T_2 ? phv_data_97 : _GEN_4204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4206 = 8'h62 == _match_key_qbytes_4_T_2 ? phv_data_98 : _GEN_4205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4207 = 8'h63 == _match_key_qbytes_4_T_2 ? phv_data_99 : _GEN_4206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4208 = 8'h64 == _match_key_qbytes_4_T_2 ? phv_data_100 : _GEN_4207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4209 = 8'h65 == _match_key_qbytes_4_T_2 ? phv_data_101 : _GEN_4208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4210 = 8'h66 == _match_key_qbytes_4_T_2 ? phv_data_102 : _GEN_4209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4211 = 8'h67 == _match_key_qbytes_4_T_2 ? phv_data_103 : _GEN_4210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4212 = 8'h68 == _match_key_qbytes_4_T_2 ? phv_data_104 : _GEN_4211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4213 = 8'h69 == _match_key_qbytes_4_T_2 ? phv_data_105 : _GEN_4212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4214 = 8'h6a == _match_key_qbytes_4_T_2 ? phv_data_106 : _GEN_4213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4215 = 8'h6b == _match_key_qbytes_4_T_2 ? phv_data_107 : _GEN_4214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4216 = 8'h6c == _match_key_qbytes_4_T_2 ? phv_data_108 : _GEN_4215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4217 = 8'h6d == _match_key_qbytes_4_T_2 ? phv_data_109 : _GEN_4216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4218 = 8'h6e == _match_key_qbytes_4_T_2 ? phv_data_110 : _GEN_4217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4219 = 8'h6f == _match_key_qbytes_4_T_2 ? phv_data_111 : _GEN_4218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4220 = 8'h70 == _match_key_qbytes_4_T_2 ? phv_data_112 : _GEN_4219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4221 = 8'h71 == _match_key_qbytes_4_T_2 ? phv_data_113 : _GEN_4220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4222 = 8'h72 == _match_key_qbytes_4_T_2 ? phv_data_114 : _GEN_4221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4223 = 8'h73 == _match_key_qbytes_4_T_2 ? phv_data_115 : _GEN_4222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4224 = 8'h74 == _match_key_qbytes_4_T_2 ? phv_data_116 : _GEN_4223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4225 = 8'h75 == _match_key_qbytes_4_T_2 ? phv_data_117 : _GEN_4224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4226 = 8'h76 == _match_key_qbytes_4_T_2 ? phv_data_118 : _GEN_4225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4227 = 8'h77 == _match_key_qbytes_4_T_2 ? phv_data_119 : _GEN_4226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4228 = 8'h78 == _match_key_qbytes_4_T_2 ? phv_data_120 : _GEN_4227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4229 = 8'h79 == _match_key_qbytes_4_T_2 ? phv_data_121 : _GEN_4228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4230 = 8'h7a == _match_key_qbytes_4_T_2 ? phv_data_122 : _GEN_4229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4231 = 8'h7b == _match_key_qbytes_4_T_2 ? phv_data_123 : _GEN_4230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4232 = 8'h7c == _match_key_qbytes_4_T_2 ? phv_data_124 : _GEN_4231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4233 = 8'h7d == _match_key_qbytes_4_T_2 ? phv_data_125 : _GEN_4232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4234 = 8'h7e == _match_key_qbytes_4_T_2 ? phv_data_126 : _GEN_4233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4235 = 8'h7f == _match_key_qbytes_4_T_2 ? phv_data_127 : _GEN_4234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4236 = 8'h80 == _match_key_qbytes_4_T_2 ? phv_data_128 : _GEN_4235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4237 = 8'h81 == _match_key_qbytes_4_T_2 ? phv_data_129 : _GEN_4236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4238 = 8'h82 == _match_key_qbytes_4_T_2 ? phv_data_130 : _GEN_4237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4239 = 8'h83 == _match_key_qbytes_4_T_2 ? phv_data_131 : _GEN_4238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4240 = 8'h84 == _match_key_qbytes_4_T_2 ? phv_data_132 : _GEN_4239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4241 = 8'h85 == _match_key_qbytes_4_T_2 ? phv_data_133 : _GEN_4240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4242 = 8'h86 == _match_key_qbytes_4_T_2 ? phv_data_134 : _GEN_4241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4243 = 8'h87 == _match_key_qbytes_4_T_2 ? phv_data_135 : _GEN_4242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4244 = 8'h88 == _match_key_qbytes_4_T_2 ? phv_data_136 : _GEN_4243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4245 = 8'h89 == _match_key_qbytes_4_T_2 ? phv_data_137 : _GEN_4244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4246 = 8'h8a == _match_key_qbytes_4_T_2 ? phv_data_138 : _GEN_4245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4247 = 8'h8b == _match_key_qbytes_4_T_2 ? phv_data_139 : _GEN_4246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4248 = 8'h8c == _match_key_qbytes_4_T_2 ? phv_data_140 : _GEN_4247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4249 = 8'h8d == _match_key_qbytes_4_T_2 ? phv_data_141 : _GEN_4248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4250 = 8'h8e == _match_key_qbytes_4_T_2 ? phv_data_142 : _GEN_4249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4251 = 8'h8f == _match_key_qbytes_4_T_2 ? phv_data_143 : _GEN_4250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4252 = 8'h90 == _match_key_qbytes_4_T_2 ? phv_data_144 : _GEN_4251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4253 = 8'h91 == _match_key_qbytes_4_T_2 ? phv_data_145 : _GEN_4252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4254 = 8'h92 == _match_key_qbytes_4_T_2 ? phv_data_146 : _GEN_4253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4255 = 8'h93 == _match_key_qbytes_4_T_2 ? phv_data_147 : _GEN_4254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4256 = 8'h94 == _match_key_qbytes_4_T_2 ? phv_data_148 : _GEN_4255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4257 = 8'h95 == _match_key_qbytes_4_T_2 ? phv_data_149 : _GEN_4256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4258 = 8'h96 == _match_key_qbytes_4_T_2 ? phv_data_150 : _GEN_4257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4259 = 8'h97 == _match_key_qbytes_4_T_2 ? phv_data_151 : _GEN_4258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4260 = 8'h98 == _match_key_qbytes_4_T_2 ? phv_data_152 : _GEN_4259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4261 = 8'h99 == _match_key_qbytes_4_T_2 ? phv_data_153 : _GEN_4260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4262 = 8'h9a == _match_key_qbytes_4_T_2 ? phv_data_154 : _GEN_4261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4263 = 8'h9b == _match_key_qbytes_4_T_2 ? phv_data_155 : _GEN_4262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4264 = 8'h9c == _match_key_qbytes_4_T_2 ? phv_data_156 : _GEN_4263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4265 = 8'h9d == _match_key_qbytes_4_T_2 ? phv_data_157 : _GEN_4264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4266 = 8'h9e == _match_key_qbytes_4_T_2 ? phv_data_158 : _GEN_4265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4267 = 8'h9f == _match_key_qbytes_4_T_2 ? phv_data_159 : _GEN_4266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4268 = 8'ha0 == _match_key_qbytes_4_T_2 ? phv_data_160 : _GEN_4267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4269 = 8'ha1 == _match_key_qbytes_4_T_2 ? phv_data_161 : _GEN_4268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4270 = 8'ha2 == _match_key_qbytes_4_T_2 ? phv_data_162 : _GEN_4269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4271 = 8'ha3 == _match_key_qbytes_4_T_2 ? phv_data_163 : _GEN_4270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4272 = 8'ha4 == _match_key_qbytes_4_T_2 ? phv_data_164 : _GEN_4271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4273 = 8'ha5 == _match_key_qbytes_4_T_2 ? phv_data_165 : _GEN_4272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4274 = 8'ha6 == _match_key_qbytes_4_T_2 ? phv_data_166 : _GEN_4273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4275 = 8'ha7 == _match_key_qbytes_4_T_2 ? phv_data_167 : _GEN_4274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4276 = 8'ha8 == _match_key_qbytes_4_T_2 ? phv_data_168 : _GEN_4275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4277 = 8'ha9 == _match_key_qbytes_4_T_2 ? phv_data_169 : _GEN_4276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4278 = 8'haa == _match_key_qbytes_4_T_2 ? phv_data_170 : _GEN_4277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4279 = 8'hab == _match_key_qbytes_4_T_2 ? phv_data_171 : _GEN_4278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4280 = 8'hac == _match_key_qbytes_4_T_2 ? phv_data_172 : _GEN_4279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4281 = 8'had == _match_key_qbytes_4_T_2 ? phv_data_173 : _GEN_4280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4282 = 8'hae == _match_key_qbytes_4_T_2 ? phv_data_174 : _GEN_4281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4283 = 8'haf == _match_key_qbytes_4_T_2 ? phv_data_175 : _GEN_4282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4284 = 8'hb0 == _match_key_qbytes_4_T_2 ? phv_data_176 : _GEN_4283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4285 = 8'hb1 == _match_key_qbytes_4_T_2 ? phv_data_177 : _GEN_4284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4286 = 8'hb2 == _match_key_qbytes_4_T_2 ? phv_data_178 : _GEN_4285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4287 = 8'hb3 == _match_key_qbytes_4_T_2 ? phv_data_179 : _GEN_4286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4288 = 8'hb4 == _match_key_qbytes_4_T_2 ? phv_data_180 : _GEN_4287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4289 = 8'hb5 == _match_key_qbytes_4_T_2 ? phv_data_181 : _GEN_4288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4290 = 8'hb6 == _match_key_qbytes_4_T_2 ? phv_data_182 : _GEN_4289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4291 = 8'hb7 == _match_key_qbytes_4_T_2 ? phv_data_183 : _GEN_4290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4292 = 8'hb8 == _match_key_qbytes_4_T_2 ? phv_data_184 : _GEN_4291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4293 = 8'hb9 == _match_key_qbytes_4_T_2 ? phv_data_185 : _GEN_4292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4294 = 8'hba == _match_key_qbytes_4_T_2 ? phv_data_186 : _GEN_4293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4295 = 8'hbb == _match_key_qbytes_4_T_2 ? phv_data_187 : _GEN_4294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4296 = 8'hbc == _match_key_qbytes_4_T_2 ? phv_data_188 : _GEN_4295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4297 = 8'hbd == _match_key_qbytes_4_T_2 ? phv_data_189 : _GEN_4296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4298 = 8'hbe == _match_key_qbytes_4_T_2 ? phv_data_190 : _GEN_4297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4299 = 8'hbf == _match_key_qbytes_4_T_2 ? phv_data_191 : _GEN_4298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4300 = 8'hc0 == _match_key_qbytes_4_T_2 ? phv_data_192 : _GEN_4299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4301 = 8'hc1 == _match_key_qbytes_4_T_2 ? phv_data_193 : _GEN_4300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4302 = 8'hc2 == _match_key_qbytes_4_T_2 ? phv_data_194 : _GEN_4301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4303 = 8'hc3 == _match_key_qbytes_4_T_2 ? phv_data_195 : _GEN_4302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4304 = 8'hc4 == _match_key_qbytes_4_T_2 ? phv_data_196 : _GEN_4303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4305 = 8'hc5 == _match_key_qbytes_4_T_2 ? phv_data_197 : _GEN_4304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4306 = 8'hc6 == _match_key_qbytes_4_T_2 ? phv_data_198 : _GEN_4305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4307 = 8'hc7 == _match_key_qbytes_4_T_2 ? phv_data_199 : _GEN_4306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4308 = 8'hc8 == _match_key_qbytes_4_T_2 ? phv_data_200 : _GEN_4307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4309 = 8'hc9 == _match_key_qbytes_4_T_2 ? phv_data_201 : _GEN_4308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4310 = 8'hca == _match_key_qbytes_4_T_2 ? phv_data_202 : _GEN_4309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4311 = 8'hcb == _match_key_qbytes_4_T_2 ? phv_data_203 : _GEN_4310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4312 = 8'hcc == _match_key_qbytes_4_T_2 ? phv_data_204 : _GEN_4311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4313 = 8'hcd == _match_key_qbytes_4_T_2 ? phv_data_205 : _GEN_4312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4314 = 8'hce == _match_key_qbytes_4_T_2 ? phv_data_206 : _GEN_4313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4315 = 8'hcf == _match_key_qbytes_4_T_2 ? phv_data_207 : _GEN_4314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4316 = 8'hd0 == _match_key_qbytes_4_T_2 ? phv_data_208 : _GEN_4315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4317 = 8'hd1 == _match_key_qbytes_4_T_2 ? phv_data_209 : _GEN_4316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4318 = 8'hd2 == _match_key_qbytes_4_T_2 ? phv_data_210 : _GEN_4317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4319 = 8'hd3 == _match_key_qbytes_4_T_2 ? phv_data_211 : _GEN_4318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4320 = 8'hd4 == _match_key_qbytes_4_T_2 ? phv_data_212 : _GEN_4319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4321 = 8'hd5 == _match_key_qbytes_4_T_2 ? phv_data_213 : _GEN_4320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4322 = 8'hd6 == _match_key_qbytes_4_T_2 ? phv_data_214 : _GEN_4321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4323 = 8'hd7 == _match_key_qbytes_4_T_2 ? phv_data_215 : _GEN_4322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4324 = 8'hd8 == _match_key_qbytes_4_T_2 ? phv_data_216 : _GEN_4323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4325 = 8'hd9 == _match_key_qbytes_4_T_2 ? phv_data_217 : _GEN_4324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4326 = 8'hda == _match_key_qbytes_4_T_2 ? phv_data_218 : _GEN_4325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4327 = 8'hdb == _match_key_qbytes_4_T_2 ? phv_data_219 : _GEN_4326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4328 = 8'hdc == _match_key_qbytes_4_T_2 ? phv_data_220 : _GEN_4327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4329 = 8'hdd == _match_key_qbytes_4_T_2 ? phv_data_221 : _GEN_4328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4330 = 8'hde == _match_key_qbytes_4_T_2 ? phv_data_222 : _GEN_4329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4331 = 8'hdf == _match_key_qbytes_4_T_2 ? phv_data_223 : _GEN_4330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4332 = 8'he0 == _match_key_qbytes_4_T_2 ? phv_data_224 : _GEN_4331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4333 = 8'he1 == _match_key_qbytes_4_T_2 ? phv_data_225 : _GEN_4332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4334 = 8'he2 == _match_key_qbytes_4_T_2 ? phv_data_226 : _GEN_4333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4335 = 8'he3 == _match_key_qbytes_4_T_2 ? phv_data_227 : _GEN_4334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4336 = 8'he4 == _match_key_qbytes_4_T_2 ? phv_data_228 : _GEN_4335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4337 = 8'he5 == _match_key_qbytes_4_T_2 ? phv_data_229 : _GEN_4336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4338 = 8'he6 == _match_key_qbytes_4_T_2 ? phv_data_230 : _GEN_4337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4339 = 8'he7 == _match_key_qbytes_4_T_2 ? phv_data_231 : _GEN_4338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4340 = 8'he8 == _match_key_qbytes_4_T_2 ? phv_data_232 : _GEN_4339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4341 = 8'he9 == _match_key_qbytes_4_T_2 ? phv_data_233 : _GEN_4340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4342 = 8'hea == _match_key_qbytes_4_T_2 ? phv_data_234 : _GEN_4341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4343 = 8'heb == _match_key_qbytes_4_T_2 ? phv_data_235 : _GEN_4342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4344 = 8'hec == _match_key_qbytes_4_T_2 ? phv_data_236 : _GEN_4343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4345 = 8'hed == _match_key_qbytes_4_T_2 ? phv_data_237 : _GEN_4344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4346 = 8'hee == _match_key_qbytes_4_T_2 ? phv_data_238 : _GEN_4345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4347 = 8'hef == _match_key_qbytes_4_T_2 ? phv_data_239 : _GEN_4346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4348 = 8'hf0 == _match_key_qbytes_4_T_2 ? phv_data_240 : _GEN_4347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4349 = 8'hf1 == _match_key_qbytes_4_T_2 ? phv_data_241 : _GEN_4348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4350 = 8'hf2 == _match_key_qbytes_4_T_2 ? phv_data_242 : _GEN_4349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4351 = 8'hf3 == _match_key_qbytes_4_T_2 ? phv_data_243 : _GEN_4350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4352 = 8'hf4 == _match_key_qbytes_4_T_2 ? phv_data_244 : _GEN_4351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4353 = 8'hf5 == _match_key_qbytes_4_T_2 ? phv_data_245 : _GEN_4352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4354 = 8'hf6 == _match_key_qbytes_4_T_2 ? phv_data_246 : _GEN_4353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4355 = 8'hf7 == _match_key_qbytes_4_T_2 ? phv_data_247 : _GEN_4354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4356 = 8'hf8 == _match_key_qbytes_4_T_2 ? phv_data_248 : _GEN_4355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4357 = 8'hf9 == _match_key_qbytes_4_T_2 ? phv_data_249 : _GEN_4356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4358 = 8'hfa == _match_key_qbytes_4_T_2 ? phv_data_250 : _GEN_4357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4359 = 8'hfb == _match_key_qbytes_4_T_2 ? phv_data_251 : _GEN_4358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4360 = 8'hfc == _match_key_qbytes_4_T_2 ? phv_data_252 : _GEN_4359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4361 = 8'hfd == _match_key_qbytes_4_T_2 ? phv_data_253 : _GEN_4360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4362 = 8'hfe == _match_key_qbytes_4_T_2 ? phv_data_254 : _GEN_4361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4363 = 8'hff == _match_key_qbytes_4_T_2 ? phv_data_255 : _GEN_4362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4365 = 8'h1 == local_offset_4 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4366 = 8'h2 == local_offset_4 ? phv_data_2 : _GEN_4365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4367 = 8'h3 == local_offset_4 ? phv_data_3 : _GEN_4366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4368 = 8'h4 == local_offset_4 ? phv_data_4 : _GEN_4367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4369 = 8'h5 == local_offset_4 ? phv_data_5 : _GEN_4368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4370 = 8'h6 == local_offset_4 ? phv_data_6 : _GEN_4369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4371 = 8'h7 == local_offset_4 ? phv_data_7 : _GEN_4370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4372 = 8'h8 == local_offset_4 ? phv_data_8 : _GEN_4371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4373 = 8'h9 == local_offset_4 ? phv_data_9 : _GEN_4372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4374 = 8'ha == local_offset_4 ? phv_data_10 : _GEN_4373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4375 = 8'hb == local_offset_4 ? phv_data_11 : _GEN_4374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4376 = 8'hc == local_offset_4 ? phv_data_12 : _GEN_4375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4377 = 8'hd == local_offset_4 ? phv_data_13 : _GEN_4376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4378 = 8'he == local_offset_4 ? phv_data_14 : _GEN_4377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4379 = 8'hf == local_offset_4 ? phv_data_15 : _GEN_4378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4380 = 8'h10 == local_offset_4 ? phv_data_16 : _GEN_4379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4381 = 8'h11 == local_offset_4 ? phv_data_17 : _GEN_4380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4382 = 8'h12 == local_offset_4 ? phv_data_18 : _GEN_4381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4383 = 8'h13 == local_offset_4 ? phv_data_19 : _GEN_4382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4384 = 8'h14 == local_offset_4 ? phv_data_20 : _GEN_4383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4385 = 8'h15 == local_offset_4 ? phv_data_21 : _GEN_4384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4386 = 8'h16 == local_offset_4 ? phv_data_22 : _GEN_4385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4387 = 8'h17 == local_offset_4 ? phv_data_23 : _GEN_4386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4388 = 8'h18 == local_offset_4 ? phv_data_24 : _GEN_4387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4389 = 8'h19 == local_offset_4 ? phv_data_25 : _GEN_4388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4390 = 8'h1a == local_offset_4 ? phv_data_26 : _GEN_4389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4391 = 8'h1b == local_offset_4 ? phv_data_27 : _GEN_4390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4392 = 8'h1c == local_offset_4 ? phv_data_28 : _GEN_4391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4393 = 8'h1d == local_offset_4 ? phv_data_29 : _GEN_4392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4394 = 8'h1e == local_offset_4 ? phv_data_30 : _GEN_4393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4395 = 8'h1f == local_offset_4 ? phv_data_31 : _GEN_4394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4396 = 8'h20 == local_offset_4 ? phv_data_32 : _GEN_4395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4397 = 8'h21 == local_offset_4 ? phv_data_33 : _GEN_4396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4398 = 8'h22 == local_offset_4 ? phv_data_34 : _GEN_4397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4399 = 8'h23 == local_offset_4 ? phv_data_35 : _GEN_4398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4400 = 8'h24 == local_offset_4 ? phv_data_36 : _GEN_4399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4401 = 8'h25 == local_offset_4 ? phv_data_37 : _GEN_4400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4402 = 8'h26 == local_offset_4 ? phv_data_38 : _GEN_4401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4403 = 8'h27 == local_offset_4 ? phv_data_39 : _GEN_4402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4404 = 8'h28 == local_offset_4 ? phv_data_40 : _GEN_4403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4405 = 8'h29 == local_offset_4 ? phv_data_41 : _GEN_4404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4406 = 8'h2a == local_offset_4 ? phv_data_42 : _GEN_4405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4407 = 8'h2b == local_offset_4 ? phv_data_43 : _GEN_4406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4408 = 8'h2c == local_offset_4 ? phv_data_44 : _GEN_4407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4409 = 8'h2d == local_offset_4 ? phv_data_45 : _GEN_4408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4410 = 8'h2e == local_offset_4 ? phv_data_46 : _GEN_4409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4411 = 8'h2f == local_offset_4 ? phv_data_47 : _GEN_4410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4412 = 8'h30 == local_offset_4 ? phv_data_48 : _GEN_4411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4413 = 8'h31 == local_offset_4 ? phv_data_49 : _GEN_4412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4414 = 8'h32 == local_offset_4 ? phv_data_50 : _GEN_4413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4415 = 8'h33 == local_offset_4 ? phv_data_51 : _GEN_4414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4416 = 8'h34 == local_offset_4 ? phv_data_52 : _GEN_4415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4417 = 8'h35 == local_offset_4 ? phv_data_53 : _GEN_4416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4418 = 8'h36 == local_offset_4 ? phv_data_54 : _GEN_4417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4419 = 8'h37 == local_offset_4 ? phv_data_55 : _GEN_4418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4420 = 8'h38 == local_offset_4 ? phv_data_56 : _GEN_4419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4421 = 8'h39 == local_offset_4 ? phv_data_57 : _GEN_4420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4422 = 8'h3a == local_offset_4 ? phv_data_58 : _GEN_4421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4423 = 8'h3b == local_offset_4 ? phv_data_59 : _GEN_4422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4424 = 8'h3c == local_offset_4 ? phv_data_60 : _GEN_4423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4425 = 8'h3d == local_offset_4 ? phv_data_61 : _GEN_4424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4426 = 8'h3e == local_offset_4 ? phv_data_62 : _GEN_4425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4427 = 8'h3f == local_offset_4 ? phv_data_63 : _GEN_4426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4428 = 8'h40 == local_offset_4 ? phv_data_64 : _GEN_4427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4429 = 8'h41 == local_offset_4 ? phv_data_65 : _GEN_4428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4430 = 8'h42 == local_offset_4 ? phv_data_66 : _GEN_4429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4431 = 8'h43 == local_offset_4 ? phv_data_67 : _GEN_4430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4432 = 8'h44 == local_offset_4 ? phv_data_68 : _GEN_4431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4433 = 8'h45 == local_offset_4 ? phv_data_69 : _GEN_4432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4434 = 8'h46 == local_offset_4 ? phv_data_70 : _GEN_4433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4435 = 8'h47 == local_offset_4 ? phv_data_71 : _GEN_4434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4436 = 8'h48 == local_offset_4 ? phv_data_72 : _GEN_4435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4437 = 8'h49 == local_offset_4 ? phv_data_73 : _GEN_4436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4438 = 8'h4a == local_offset_4 ? phv_data_74 : _GEN_4437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4439 = 8'h4b == local_offset_4 ? phv_data_75 : _GEN_4438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4440 = 8'h4c == local_offset_4 ? phv_data_76 : _GEN_4439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4441 = 8'h4d == local_offset_4 ? phv_data_77 : _GEN_4440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4442 = 8'h4e == local_offset_4 ? phv_data_78 : _GEN_4441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4443 = 8'h4f == local_offset_4 ? phv_data_79 : _GEN_4442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4444 = 8'h50 == local_offset_4 ? phv_data_80 : _GEN_4443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4445 = 8'h51 == local_offset_4 ? phv_data_81 : _GEN_4444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4446 = 8'h52 == local_offset_4 ? phv_data_82 : _GEN_4445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4447 = 8'h53 == local_offset_4 ? phv_data_83 : _GEN_4446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4448 = 8'h54 == local_offset_4 ? phv_data_84 : _GEN_4447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4449 = 8'h55 == local_offset_4 ? phv_data_85 : _GEN_4448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4450 = 8'h56 == local_offset_4 ? phv_data_86 : _GEN_4449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4451 = 8'h57 == local_offset_4 ? phv_data_87 : _GEN_4450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4452 = 8'h58 == local_offset_4 ? phv_data_88 : _GEN_4451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4453 = 8'h59 == local_offset_4 ? phv_data_89 : _GEN_4452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4454 = 8'h5a == local_offset_4 ? phv_data_90 : _GEN_4453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4455 = 8'h5b == local_offset_4 ? phv_data_91 : _GEN_4454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4456 = 8'h5c == local_offset_4 ? phv_data_92 : _GEN_4455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4457 = 8'h5d == local_offset_4 ? phv_data_93 : _GEN_4456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4458 = 8'h5e == local_offset_4 ? phv_data_94 : _GEN_4457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4459 = 8'h5f == local_offset_4 ? phv_data_95 : _GEN_4458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4460 = 8'h60 == local_offset_4 ? phv_data_96 : _GEN_4459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4461 = 8'h61 == local_offset_4 ? phv_data_97 : _GEN_4460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4462 = 8'h62 == local_offset_4 ? phv_data_98 : _GEN_4461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4463 = 8'h63 == local_offset_4 ? phv_data_99 : _GEN_4462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4464 = 8'h64 == local_offset_4 ? phv_data_100 : _GEN_4463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4465 = 8'h65 == local_offset_4 ? phv_data_101 : _GEN_4464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4466 = 8'h66 == local_offset_4 ? phv_data_102 : _GEN_4465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4467 = 8'h67 == local_offset_4 ? phv_data_103 : _GEN_4466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4468 = 8'h68 == local_offset_4 ? phv_data_104 : _GEN_4467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4469 = 8'h69 == local_offset_4 ? phv_data_105 : _GEN_4468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4470 = 8'h6a == local_offset_4 ? phv_data_106 : _GEN_4469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4471 = 8'h6b == local_offset_4 ? phv_data_107 : _GEN_4470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4472 = 8'h6c == local_offset_4 ? phv_data_108 : _GEN_4471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4473 = 8'h6d == local_offset_4 ? phv_data_109 : _GEN_4472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4474 = 8'h6e == local_offset_4 ? phv_data_110 : _GEN_4473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4475 = 8'h6f == local_offset_4 ? phv_data_111 : _GEN_4474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4476 = 8'h70 == local_offset_4 ? phv_data_112 : _GEN_4475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4477 = 8'h71 == local_offset_4 ? phv_data_113 : _GEN_4476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4478 = 8'h72 == local_offset_4 ? phv_data_114 : _GEN_4477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4479 = 8'h73 == local_offset_4 ? phv_data_115 : _GEN_4478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4480 = 8'h74 == local_offset_4 ? phv_data_116 : _GEN_4479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4481 = 8'h75 == local_offset_4 ? phv_data_117 : _GEN_4480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4482 = 8'h76 == local_offset_4 ? phv_data_118 : _GEN_4481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4483 = 8'h77 == local_offset_4 ? phv_data_119 : _GEN_4482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4484 = 8'h78 == local_offset_4 ? phv_data_120 : _GEN_4483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4485 = 8'h79 == local_offset_4 ? phv_data_121 : _GEN_4484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4486 = 8'h7a == local_offset_4 ? phv_data_122 : _GEN_4485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4487 = 8'h7b == local_offset_4 ? phv_data_123 : _GEN_4486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4488 = 8'h7c == local_offset_4 ? phv_data_124 : _GEN_4487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4489 = 8'h7d == local_offset_4 ? phv_data_125 : _GEN_4488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4490 = 8'h7e == local_offset_4 ? phv_data_126 : _GEN_4489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4491 = 8'h7f == local_offset_4 ? phv_data_127 : _GEN_4490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4492 = 8'h80 == local_offset_4 ? phv_data_128 : _GEN_4491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4493 = 8'h81 == local_offset_4 ? phv_data_129 : _GEN_4492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4494 = 8'h82 == local_offset_4 ? phv_data_130 : _GEN_4493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4495 = 8'h83 == local_offset_4 ? phv_data_131 : _GEN_4494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4496 = 8'h84 == local_offset_4 ? phv_data_132 : _GEN_4495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4497 = 8'h85 == local_offset_4 ? phv_data_133 : _GEN_4496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4498 = 8'h86 == local_offset_4 ? phv_data_134 : _GEN_4497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4499 = 8'h87 == local_offset_4 ? phv_data_135 : _GEN_4498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4500 = 8'h88 == local_offset_4 ? phv_data_136 : _GEN_4499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4501 = 8'h89 == local_offset_4 ? phv_data_137 : _GEN_4500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4502 = 8'h8a == local_offset_4 ? phv_data_138 : _GEN_4501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4503 = 8'h8b == local_offset_4 ? phv_data_139 : _GEN_4502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4504 = 8'h8c == local_offset_4 ? phv_data_140 : _GEN_4503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4505 = 8'h8d == local_offset_4 ? phv_data_141 : _GEN_4504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4506 = 8'h8e == local_offset_4 ? phv_data_142 : _GEN_4505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4507 = 8'h8f == local_offset_4 ? phv_data_143 : _GEN_4506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4508 = 8'h90 == local_offset_4 ? phv_data_144 : _GEN_4507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4509 = 8'h91 == local_offset_4 ? phv_data_145 : _GEN_4508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4510 = 8'h92 == local_offset_4 ? phv_data_146 : _GEN_4509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4511 = 8'h93 == local_offset_4 ? phv_data_147 : _GEN_4510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4512 = 8'h94 == local_offset_4 ? phv_data_148 : _GEN_4511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4513 = 8'h95 == local_offset_4 ? phv_data_149 : _GEN_4512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4514 = 8'h96 == local_offset_4 ? phv_data_150 : _GEN_4513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4515 = 8'h97 == local_offset_4 ? phv_data_151 : _GEN_4514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4516 = 8'h98 == local_offset_4 ? phv_data_152 : _GEN_4515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4517 = 8'h99 == local_offset_4 ? phv_data_153 : _GEN_4516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4518 = 8'h9a == local_offset_4 ? phv_data_154 : _GEN_4517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4519 = 8'h9b == local_offset_4 ? phv_data_155 : _GEN_4518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4520 = 8'h9c == local_offset_4 ? phv_data_156 : _GEN_4519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4521 = 8'h9d == local_offset_4 ? phv_data_157 : _GEN_4520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4522 = 8'h9e == local_offset_4 ? phv_data_158 : _GEN_4521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4523 = 8'h9f == local_offset_4 ? phv_data_159 : _GEN_4522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4524 = 8'ha0 == local_offset_4 ? phv_data_160 : _GEN_4523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4525 = 8'ha1 == local_offset_4 ? phv_data_161 : _GEN_4524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4526 = 8'ha2 == local_offset_4 ? phv_data_162 : _GEN_4525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4527 = 8'ha3 == local_offset_4 ? phv_data_163 : _GEN_4526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4528 = 8'ha4 == local_offset_4 ? phv_data_164 : _GEN_4527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4529 = 8'ha5 == local_offset_4 ? phv_data_165 : _GEN_4528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4530 = 8'ha6 == local_offset_4 ? phv_data_166 : _GEN_4529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4531 = 8'ha7 == local_offset_4 ? phv_data_167 : _GEN_4530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4532 = 8'ha8 == local_offset_4 ? phv_data_168 : _GEN_4531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4533 = 8'ha9 == local_offset_4 ? phv_data_169 : _GEN_4532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4534 = 8'haa == local_offset_4 ? phv_data_170 : _GEN_4533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4535 = 8'hab == local_offset_4 ? phv_data_171 : _GEN_4534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4536 = 8'hac == local_offset_4 ? phv_data_172 : _GEN_4535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4537 = 8'had == local_offset_4 ? phv_data_173 : _GEN_4536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4538 = 8'hae == local_offset_4 ? phv_data_174 : _GEN_4537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4539 = 8'haf == local_offset_4 ? phv_data_175 : _GEN_4538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4540 = 8'hb0 == local_offset_4 ? phv_data_176 : _GEN_4539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4541 = 8'hb1 == local_offset_4 ? phv_data_177 : _GEN_4540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4542 = 8'hb2 == local_offset_4 ? phv_data_178 : _GEN_4541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4543 = 8'hb3 == local_offset_4 ? phv_data_179 : _GEN_4542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4544 = 8'hb4 == local_offset_4 ? phv_data_180 : _GEN_4543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4545 = 8'hb5 == local_offset_4 ? phv_data_181 : _GEN_4544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4546 = 8'hb6 == local_offset_4 ? phv_data_182 : _GEN_4545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4547 = 8'hb7 == local_offset_4 ? phv_data_183 : _GEN_4546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4548 = 8'hb8 == local_offset_4 ? phv_data_184 : _GEN_4547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4549 = 8'hb9 == local_offset_4 ? phv_data_185 : _GEN_4548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4550 = 8'hba == local_offset_4 ? phv_data_186 : _GEN_4549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4551 = 8'hbb == local_offset_4 ? phv_data_187 : _GEN_4550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4552 = 8'hbc == local_offset_4 ? phv_data_188 : _GEN_4551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4553 = 8'hbd == local_offset_4 ? phv_data_189 : _GEN_4552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4554 = 8'hbe == local_offset_4 ? phv_data_190 : _GEN_4553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4555 = 8'hbf == local_offset_4 ? phv_data_191 : _GEN_4554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4556 = 8'hc0 == local_offset_4 ? phv_data_192 : _GEN_4555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4557 = 8'hc1 == local_offset_4 ? phv_data_193 : _GEN_4556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4558 = 8'hc2 == local_offset_4 ? phv_data_194 : _GEN_4557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4559 = 8'hc3 == local_offset_4 ? phv_data_195 : _GEN_4558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4560 = 8'hc4 == local_offset_4 ? phv_data_196 : _GEN_4559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4561 = 8'hc5 == local_offset_4 ? phv_data_197 : _GEN_4560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4562 = 8'hc6 == local_offset_4 ? phv_data_198 : _GEN_4561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4563 = 8'hc7 == local_offset_4 ? phv_data_199 : _GEN_4562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4564 = 8'hc8 == local_offset_4 ? phv_data_200 : _GEN_4563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4565 = 8'hc9 == local_offset_4 ? phv_data_201 : _GEN_4564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4566 = 8'hca == local_offset_4 ? phv_data_202 : _GEN_4565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4567 = 8'hcb == local_offset_4 ? phv_data_203 : _GEN_4566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4568 = 8'hcc == local_offset_4 ? phv_data_204 : _GEN_4567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4569 = 8'hcd == local_offset_4 ? phv_data_205 : _GEN_4568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4570 = 8'hce == local_offset_4 ? phv_data_206 : _GEN_4569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4571 = 8'hcf == local_offset_4 ? phv_data_207 : _GEN_4570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4572 = 8'hd0 == local_offset_4 ? phv_data_208 : _GEN_4571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4573 = 8'hd1 == local_offset_4 ? phv_data_209 : _GEN_4572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4574 = 8'hd2 == local_offset_4 ? phv_data_210 : _GEN_4573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4575 = 8'hd3 == local_offset_4 ? phv_data_211 : _GEN_4574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4576 = 8'hd4 == local_offset_4 ? phv_data_212 : _GEN_4575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4577 = 8'hd5 == local_offset_4 ? phv_data_213 : _GEN_4576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4578 = 8'hd6 == local_offset_4 ? phv_data_214 : _GEN_4577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4579 = 8'hd7 == local_offset_4 ? phv_data_215 : _GEN_4578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4580 = 8'hd8 == local_offset_4 ? phv_data_216 : _GEN_4579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4581 = 8'hd9 == local_offset_4 ? phv_data_217 : _GEN_4580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4582 = 8'hda == local_offset_4 ? phv_data_218 : _GEN_4581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4583 = 8'hdb == local_offset_4 ? phv_data_219 : _GEN_4582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4584 = 8'hdc == local_offset_4 ? phv_data_220 : _GEN_4583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4585 = 8'hdd == local_offset_4 ? phv_data_221 : _GEN_4584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4586 = 8'hde == local_offset_4 ? phv_data_222 : _GEN_4585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4587 = 8'hdf == local_offset_4 ? phv_data_223 : _GEN_4586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4588 = 8'he0 == local_offset_4 ? phv_data_224 : _GEN_4587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4589 = 8'he1 == local_offset_4 ? phv_data_225 : _GEN_4588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4590 = 8'he2 == local_offset_4 ? phv_data_226 : _GEN_4589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4591 = 8'he3 == local_offset_4 ? phv_data_227 : _GEN_4590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4592 = 8'he4 == local_offset_4 ? phv_data_228 : _GEN_4591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4593 = 8'he5 == local_offset_4 ? phv_data_229 : _GEN_4592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4594 = 8'he6 == local_offset_4 ? phv_data_230 : _GEN_4593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4595 = 8'he7 == local_offset_4 ? phv_data_231 : _GEN_4594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4596 = 8'he8 == local_offset_4 ? phv_data_232 : _GEN_4595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4597 = 8'he9 == local_offset_4 ? phv_data_233 : _GEN_4596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4598 = 8'hea == local_offset_4 ? phv_data_234 : _GEN_4597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4599 = 8'heb == local_offset_4 ? phv_data_235 : _GEN_4598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4600 = 8'hec == local_offset_4 ? phv_data_236 : _GEN_4599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4601 = 8'hed == local_offset_4 ? phv_data_237 : _GEN_4600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4602 = 8'hee == local_offset_4 ? phv_data_238 : _GEN_4601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4603 = 8'hef == local_offset_4 ? phv_data_239 : _GEN_4602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4604 = 8'hf0 == local_offset_4 ? phv_data_240 : _GEN_4603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4605 = 8'hf1 == local_offset_4 ? phv_data_241 : _GEN_4604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4606 = 8'hf2 == local_offset_4 ? phv_data_242 : _GEN_4605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4607 = 8'hf3 == local_offset_4 ? phv_data_243 : _GEN_4606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4608 = 8'hf4 == local_offset_4 ? phv_data_244 : _GEN_4607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4609 = 8'hf5 == local_offset_4 ? phv_data_245 : _GEN_4608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4610 = 8'hf6 == local_offset_4 ? phv_data_246 : _GEN_4609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4611 = 8'hf7 == local_offset_4 ? phv_data_247 : _GEN_4610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4612 = 8'hf8 == local_offset_4 ? phv_data_248 : _GEN_4611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4613 = 8'hf9 == local_offset_4 ? phv_data_249 : _GEN_4612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4614 = 8'hfa == local_offset_4 ? phv_data_250 : _GEN_4613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4615 = 8'hfb == local_offset_4 ? phv_data_251 : _GEN_4614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4616 = 8'hfc == local_offset_4 ? phv_data_252 : _GEN_4615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4617 = 8'hfd == local_offset_4 ? phv_data_253 : _GEN_4616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4618 = 8'hfe == local_offset_4 ? phv_data_254 : _GEN_4617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4619 = 8'hff == local_offset_4 ? phv_data_255 : _GEN_4618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4621 = 8'h1 == _match_key_qbytes_4_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4622 = 8'h2 == _match_key_qbytes_4_T ? phv_data_2 : _GEN_4621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4623 = 8'h3 == _match_key_qbytes_4_T ? phv_data_3 : _GEN_4622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4624 = 8'h4 == _match_key_qbytes_4_T ? phv_data_4 : _GEN_4623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4625 = 8'h5 == _match_key_qbytes_4_T ? phv_data_5 : _GEN_4624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4626 = 8'h6 == _match_key_qbytes_4_T ? phv_data_6 : _GEN_4625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4627 = 8'h7 == _match_key_qbytes_4_T ? phv_data_7 : _GEN_4626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4628 = 8'h8 == _match_key_qbytes_4_T ? phv_data_8 : _GEN_4627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4629 = 8'h9 == _match_key_qbytes_4_T ? phv_data_9 : _GEN_4628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4630 = 8'ha == _match_key_qbytes_4_T ? phv_data_10 : _GEN_4629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4631 = 8'hb == _match_key_qbytes_4_T ? phv_data_11 : _GEN_4630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4632 = 8'hc == _match_key_qbytes_4_T ? phv_data_12 : _GEN_4631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4633 = 8'hd == _match_key_qbytes_4_T ? phv_data_13 : _GEN_4632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4634 = 8'he == _match_key_qbytes_4_T ? phv_data_14 : _GEN_4633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4635 = 8'hf == _match_key_qbytes_4_T ? phv_data_15 : _GEN_4634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4636 = 8'h10 == _match_key_qbytes_4_T ? phv_data_16 : _GEN_4635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4637 = 8'h11 == _match_key_qbytes_4_T ? phv_data_17 : _GEN_4636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4638 = 8'h12 == _match_key_qbytes_4_T ? phv_data_18 : _GEN_4637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4639 = 8'h13 == _match_key_qbytes_4_T ? phv_data_19 : _GEN_4638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4640 = 8'h14 == _match_key_qbytes_4_T ? phv_data_20 : _GEN_4639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4641 = 8'h15 == _match_key_qbytes_4_T ? phv_data_21 : _GEN_4640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4642 = 8'h16 == _match_key_qbytes_4_T ? phv_data_22 : _GEN_4641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4643 = 8'h17 == _match_key_qbytes_4_T ? phv_data_23 : _GEN_4642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4644 = 8'h18 == _match_key_qbytes_4_T ? phv_data_24 : _GEN_4643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4645 = 8'h19 == _match_key_qbytes_4_T ? phv_data_25 : _GEN_4644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4646 = 8'h1a == _match_key_qbytes_4_T ? phv_data_26 : _GEN_4645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4647 = 8'h1b == _match_key_qbytes_4_T ? phv_data_27 : _GEN_4646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4648 = 8'h1c == _match_key_qbytes_4_T ? phv_data_28 : _GEN_4647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4649 = 8'h1d == _match_key_qbytes_4_T ? phv_data_29 : _GEN_4648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4650 = 8'h1e == _match_key_qbytes_4_T ? phv_data_30 : _GEN_4649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4651 = 8'h1f == _match_key_qbytes_4_T ? phv_data_31 : _GEN_4650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4652 = 8'h20 == _match_key_qbytes_4_T ? phv_data_32 : _GEN_4651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4653 = 8'h21 == _match_key_qbytes_4_T ? phv_data_33 : _GEN_4652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4654 = 8'h22 == _match_key_qbytes_4_T ? phv_data_34 : _GEN_4653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4655 = 8'h23 == _match_key_qbytes_4_T ? phv_data_35 : _GEN_4654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4656 = 8'h24 == _match_key_qbytes_4_T ? phv_data_36 : _GEN_4655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4657 = 8'h25 == _match_key_qbytes_4_T ? phv_data_37 : _GEN_4656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4658 = 8'h26 == _match_key_qbytes_4_T ? phv_data_38 : _GEN_4657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4659 = 8'h27 == _match_key_qbytes_4_T ? phv_data_39 : _GEN_4658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4660 = 8'h28 == _match_key_qbytes_4_T ? phv_data_40 : _GEN_4659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4661 = 8'h29 == _match_key_qbytes_4_T ? phv_data_41 : _GEN_4660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4662 = 8'h2a == _match_key_qbytes_4_T ? phv_data_42 : _GEN_4661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4663 = 8'h2b == _match_key_qbytes_4_T ? phv_data_43 : _GEN_4662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4664 = 8'h2c == _match_key_qbytes_4_T ? phv_data_44 : _GEN_4663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4665 = 8'h2d == _match_key_qbytes_4_T ? phv_data_45 : _GEN_4664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4666 = 8'h2e == _match_key_qbytes_4_T ? phv_data_46 : _GEN_4665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4667 = 8'h2f == _match_key_qbytes_4_T ? phv_data_47 : _GEN_4666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4668 = 8'h30 == _match_key_qbytes_4_T ? phv_data_48 : _GEN_4667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4669 = 8'h31 == _match_key_qbytes_4_T ? phv_data_49 : _GEN_4668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4670 = 8'h32 == _match_key_qbytes_4_T ? phv_data_50 : _GEN_4669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4671 = 8'h33 == _match_key_qbytes_4_T ? phv_data_51 : _GEN_4670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4672 = 8'h34 == _match_key_qbytes_4_T ? phv_data_52 : _GEN_4671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4673 = 8'h35 == _match_key_qbytes_4_T ? phv_data_53 : _GEN_4672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4674 = 8'h36 == _match_key_qbytes_4_T ? phv_data_54 : _GEN_4673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4675 = 8'h37 == _match_key_qbytes_4_T ? phv_data_55 : _GEN_4674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4676 = 8'h38 == _match_key_qbytes_4_T ? phv_data_56 : _GEN_4675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4677 = 8'h39 == _match_key_qbytes_4_T ? phv_data_57 : _GEN_4676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4678 = 8'h3a == _match_key_qbytes_4_T ? phv_data_58 : _GEN_4677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4679 = 8'h3b == _match_key_qbytes_4_T ? phv_data_59 : _GEN_4678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4680 = 8'h3c == _match_key_qbytes_4_T ? phv_data_60 : _GEN_4679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4681 = 8'h3d == _match_key_qbytes_4_T ? phv_data_61 : _GEN_4680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4682 = 8'h3e == _match_key_qbytes_4_T ? phv_data_62 : _GEN_4681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4683 = 8'h3f == _match_key_qbytes_4_T ? phv_data_63 : _GEN_4682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4684 = 8'h40 == _match_key_qbytes_4_T ? phv_data_64 : _GEN_4683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4685 = 8'h41 == _match_key_qbytes_4_T ? phv_data_65 : _GEN_4684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4686 = 8'h42 == _match_key_qbytes_4_T ? phv_data_66 : _GEN_4685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4687 = 8'h43 == _match_key_qbytes_4_T ? phv_data_67 : _GEN_4686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4688 = 8'h44 == _match_key_qbytes_4_T ? phv_data_68 : _GEN_4687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4689 = 8'h45 == _match_key_qbytes_4_T ? phv_data_69 : _GEN_4688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4690 = 8'h46 == _match_key_qbytes_4_T ? phv_data_70 : _GEN_4689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4691 = 8'h47 == _match_key_qbytes_4_T ? phv_data_71 : _GEN_4690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4692 = 8'h48 == _match_key_qbytes_4_T ? phv_data_72 : _GEN_4691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4693 = 8'h49 == _match_key_qbytes_4_T ? phv_data_73 : _GEN_4692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4694 = 8'h4a == _match_key_qbytes_4_T ? phv_data_74 : _GEN_4693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4695 = 8'h4b == _match_key_qbytes_4_T ? phv_data_75 : _GEN_4694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4696 = 8'h4c == _match_key_qbytes_4_T ? phv_data_76 : _GEN_4695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4697 = 8'h4d == _match_key_qbytes_4_T ? phv_data_77 : _GEN_4696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4698 = 8'h4e == _match_key_qbytes_4_T ? phv_data_78 : _GEN_4697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4699 = 8'h4f == _match_key_qbytes_4_T ? phv_data_79 : _GEN_4698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4700 = 8'h50 == _match_key_qbytes_4_T ? phv_data_80 : _GEN_4699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4701 = 8'h51 == _match_key_qbytes_4_T ? phv_data_81 : _GEN_4700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4702 = 8'h52 == _match_key_qbytes_4_T ? phv_data_82 : _GEN_4701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4703 = 8'h53 == _match_key_qbytes_4_T ? phv_data_83 : _GEN_4702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4704 = 8'h54 == _match_key_qbytes_4_T ? phv_data_84 : _GEN_4703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4705 = 8'h55 == _match_key_qbytes_4_T ? phv_data_85 : _GEN_4704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4706 = 8'h56 == _match_key_qbytes_4_T ? phv_data_86 : _GEN_4705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4707 = 8'h57 == _match_key_qbytes_4_T ? phv_data_87 : _GEN_4706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4708 = 8'h58 == _match_key_qbytes_4_T ? phv_data_88 : _GEN_4707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4709 = 8'h59 == _match_key_qbytes_4_T ? phv_data_89 : _GEN_4708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4710 = 8'h5a == _match_key_qbytes_4_T ? phv_data_90 : _GEN_4709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4711 = 8'h5b == _match_key_qbytes_4_T ? phv_data_91 : _GEN_4710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4712 = 8'h5c == _match_key_qbytes_4_T ? phv_data_92 : _GEN_4711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4713 = 8'h5d == _match_key_qbytes_4_T ? phv_data_93 : _GEN_4712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4714 = 8'h5e == _match_key_qbytes_4_T ? phv_data_94 : _GEN_4713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4715 = 8'h5f == _match_key_qbytes_4_T ? phv_data_95 : _GEN_4714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4716 = 8'h60 == _match_key_qbytes_4_T ? phv_data_96 : _GEN_4715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4717 = 8'h61 == _match_key_qbytes_4_T ? phv_data_97 : _GEN_4716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4718 = 8'h62 == _match_key_qbytes_4_T ? phv_data_98 : _GEN_4717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4719 = 8'h63 == _match_key_qbytes_4_T ? phv_data_99 : _GEN_4718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4720 = 8'h64 == _match_key_qbytes_4_T ? phv_data_100 : _GEN_4719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4721 = 8'h65 == _match_key_qbytes_4_T ? phv_data_101 : _GEN_4720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4722 = 8'h66 == _match_key_qbytes_4_T ? phv_data_102 : _GEN_4721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4723 = 8'h67 == _match_key_qbytes_4_T ? phv_data_103 : _GEN_4722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4724 = 8'h68 == _match_key_qbytes_4_T ? phv_data_104 : _GEN_4723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4725 = 8'h69 == _match_key_qbytes_4_T ? phv_data_105 : _GEN_4724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4726 = 8'h6a == _match_key_qbytes_4_T ? phv_data_106 : _GEN_4725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4727 = 8'h6b == _match_key_qbytes_4_T ? phv_data_107 : _GEN_4726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4728 = 8'h6c == _match_key_qbytes_4_T ? phv_data_108 : _GEN_4727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4729 = 8'h6d == _match_key_qbytes_4_T ? phv_data_109 : _GEN_4728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4730 = 8'h6e == _match_key_qbytes_4_T ? phv_data_110 : _GEN_4729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4731 = 8'h6f == _match_key_qbytes_4_T ? phv_data_111 : _GEN_4730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4732 = 8'h70 == _match_key_qbytes_4_T ? phv_data_112 : _GEN_4731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4733 = 8'h71 == _match_key_qbytes_4_T ? phv_data_113 : _GEN_4732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4734 = 8'h72 == _match_key_qbytes_4_T ? phv_data_114 : _GEN_4733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4735 = 8'h73 == _match_key_qbytes_4_T ? phv_data_115 : _GEN_4734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4736 = 8'h74 == _match_key_qbytes_4_T ? phv_data_116 : _GEN_4735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4737 = 8'h75 == _match_key_qbytes_4_T ? phv_data_117 : _GEN_4736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4738 = 8'h76 == _match_key_qbytes_4_T ? phv_data_118 : _GEN_4737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4739 = 8'h77 == _match_key_qbytes_4_T ? phv_data_119 : _GEN_4738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4740 = 8'h78 == _match_key_qbytes_4_T ? phv_data_120 : _GEN_4739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4741 = 8'h79 == _match_key_qbytes_4_T ? phv_data_121 : _GEN_4740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4742 = 8'h7a == _match_key_qbytes_4_T ? phv_data_122 : _GEN_4741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4743 = 8'h7b == _match_key_qbytes_4_T ? phv_data_123 : _GEN_4742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4744 = 8'h7c == _match_key_qbytes_4_T ? phv_data_124 : _GEN_4743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4745 = 8'h7d == _match_key_qbytes_4_T ? phv_data_125 : _GEN_4744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4746 = 8'h7e == _match_key_qbytes_4_T ? phv_data_126 : _GEN_4745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4747 = 8'h7f == _match_key_qbytes_4_T ? phv_data_127 : _GEN_4746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4748 = 8'h80 == _match_key_qbytes_4_T ? phv_data_128 : _GEN_4747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4749 = 8'h81 == _match_key_qbytes_4_T ? phv_data_129 : _GEN_4748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4750 = 8'h82 == _match_key_qbytes_4_T ? phv_data_130 : _GEN_4749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4751 = 8'h83 == _match_key_qbytes_4_T ? phv_data_131 : _GEN_4750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4752 = 8'h84 == _match_key_qbytes_4_T ? phv_data_132 : _GEN_4751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4753 = 8'h85 == _match_key_qbytes_4_T ? phv_data_133 : _GEN_4752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4754 = 8'h86 == _match_key_qbytes_4_T ? phv_data_134 : _GEN_4753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4755 = 8'h87 == _match_key_qbytes_4_T ? phv_data_135 : _GEN_4754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4756 = 8'h88 == _match_key_qbytes_4_T ? phv_data_136 : _GEN_4755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4757 = 8'h89 == _match_key_qbytes_4_T ? phv_data_137 : _GEN_4756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4758 = 8'h8a == _match_key_qbytes_4_T ? phv_data_138 : _GEN_4757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4759 = 8'h8b == _match_key_qbytes_4_T ? phv_data_139 : _GEN_4758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4760 = 8'h8c == _match_key_qbytes_4_T ? phv_data_140 : _GEN_4759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4761 = 8'h8d == _match_key_qbytes_4_T ? phv_data_141 : _GEN_4760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4762 = 8'h8e == _match_key_qbytes_4_T ? phv_data_142 : _GEN_4761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4763 = 8'h8f == _match_key_qbytes_4_T ? phv_data_143 : _GEN_4762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4764 = 8'h90 == _match_key_qbytes_4_T ? phv_data_144 : _GEN_4763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4765 = 8'h91 == _match_key_qbytes_4_T ? phv_data_145 : _GEN_4764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4766 = 8'h92 == _match_key_qbytes_4_T ? phv_data_146 : _GEN_4765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4767 = 8'h93 == _match_key_qbytes_4_T ? phv_data_147 : _GEN_4766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4768 = 8'h94 == _match_key_qbytes_4_T ? phv_data_148 : _GEN_4767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4769 = 8'h95 == _match_key_qbytes_4_T ? phv_data_149 : _GEN_4768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4770 = 8'h96 == _match_key_qbytes_4_T ? phv_data_150 : _GEN_4769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4771 = 8'h97 == _match_key_qbytes_4_T ? phv_data_151 : _GEN_4770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4772 = 8'h98 == _match_key_qbytes_4_T ? phv_data_152 : _GEN_4771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4773 = 8'h99 == _match_key_qbytes_4_T ? phv_data_153 : _GEN_4772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4774 = 8'h9a == _match_key_qbytes_4_T ? phv_data_154 : _GEN_4773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4775 = 8'h9b == _match_key_qbytes_4_T ? phv_data_155 : _GEN_4774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4776 = 8'h9c == _match_key_qbytes_4_T ? phv_data_156 : _GEN_4775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4777 = 8'h9d == _match_key_qbytes_4_T ? phv_data_157 : _GEN_4776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4778 = 8'h9e == _match_key_qbytes_4_T ? phv_data_158 : _GEN_4777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4779 = 8'h9f == _match_key_qbytes_4_T ? phv_data_159 : _GEN_4778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4780 = 8'ha0 == _match_key_qbytes_4_T ? phv_data_160 : _GEN_4779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4781 = 8'ha1 == _match_key_qbytes_4_T ? phv_data_161 : _GEN_4780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4782 = 8'ha2 == _match_key_qbytes_4_T ? phv_data_162 : _GEN_4781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4783 = 8'ha3 == _match_key_qbytes_4_T ? phv_data_163 : _GEN_4782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4784 = 8'ha4 == _match_key_qbytes_4_T ? phv_data_164 : _GEN_4783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4785 = 8'ha5 == _match_key_qbytes_4_T ? phv_data_165 : _GEN_4784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4786 = 8'ha6 == _match_key_qbytes_4_T ? phv_data_166 : _GEN_4785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4787 = 8'ha7 == _match_key_qbytes_4_T ? phv_data_167 : _GEN_4786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4788 = 8'ha8 == _match_key_qbytes_4_T ? phv_data_168 : _GEN_4787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4789 = 8'ha9 == _match_key_qbytes_4_T ? phv_data_169 : _GEN_4788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4790 = 8'haa == _match_key_qbytes_4_T ? phv_data_170 : _GEN_4789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4791 = 8'hab == _match_key_qbytes_4_T ? phv_data_171 : _GEN_4790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4792 = 8'hac == _match_key_qbytes_4_T ? phv_data_172 : _GEN_4791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4793 = 8'had == _match_key_qbytes_4_T ? phv_data_173 : _GEN_4792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4794 = 8'hae == _match_key_qbytes_4_T ? phv_data_174 : _GEN_4793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4795 = 8'haf == _match_key_qbytes_4_T ? phv_data_175 : _GEN_4794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4796 = 8'hb0 == _match_key_qbytes_4_T ? phv_data_176 : _GEN_4795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4797 = 8'hb1 == _match_key_qbytes_4_T ? phv_data_177 : _GEN_4796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4798 = 8'hb2 == _match_key_qbytes_4_T ? phv_data_178 : _GEN_4797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4799 = 8'hb3 == _match_key_qbytes_4_T ? phv_data_179 : _GEN_4798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4800 = 8'hb4 == _match_key_qbytes_4_T ? phv_data_180 : _GEN_4799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4801 = 8'hb5 == _match_key_qbytes_4_T ? phv_data_181 : _GEN_4800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4802 = 8'hb6 == _match_key_qbytes_4_T ? phv_data_182 : _GEN_4801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4803 = 8'hb7 == _match_key_qbytes_4_T ? phv_data_183 : _GEN_4802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4804 = 8'hb8 == _match_key_qbytes_4_T ? phv_data_184 : _GEN_4803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4805 = 8'hb9 == _match_key_qbytes_4_T ? phv_data_185 : _GEN_4804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4806 = 8'hba == _match_key_qbytes_4_T ? phv_data_186 : _GEN_4805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4807 = 8'hbb == _match_key_qbytes_4_T ? phv_data_187 : _GEN_4806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4808 = 8'hbc == _match_key_qbytes_4_T ? phv_data_188 : _GEN_4807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4809 = 8'hbd == _match_key_qbytes_4_T ? phv_data_189 : _GEN_4808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4810 = 8'hbe == _match_key_qbytes_4_T ? phv_data_190 : _GEN_4809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4811 = 8'hbf == _match_key_qbytes_4_T ? phv_data_191 : _GEN_4810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4812 = 8'hc0 == _match_key_qbytes_4_T ? phv_data_192 : _GEN_4811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4813 = 8'hc1 == _match_key_qbytes_4_T ? phv_data_193 : _GEN_4812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4814 = 8'hc2 == _match_key_qbytes_4_T ? phv_data_194 : _GEN_4813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4815 = 8'hc3 == _match_key_qbytes_4_T ? phv_data_195 : _GEN_4814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4816 = 8'hc4 == _match_key_qbytes_4_T ? phv_data_196 : _GEN_4815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4817 = 8'hc5 == _match_key_qbytes_4_T ? phv_data_197 : _GEN_4816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4818 = 8'hc6 == _match_key_qbytes_4_T ? phv_data_198 : _GEN_4817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4819 = 8'hc7 == _match_key_qbytes_4_T ? phv_data_199 : _GEN_4818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4820 = 8'hc8 == _match_key_qbytes_4_T ? phv_data_200 : _GEN_4819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4821 = 8'hc9 == _match_key_qbytes_4_T ? phv_data_201 : _GEN_4820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4822 = 8'hca == _match_key_qbytes_4_T ? phv_data_202 : _GEN_4821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4823 = 8'hcb == _match_key_qbytes_4_T ? phv_data_203 : _GEN_4822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4824 = 8'hcc == _match_key_qbytes_4_T ? phv_data_204 : _GEN_4823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4825 = 8'hcd == _match_key_qbytes_4_T ? phv_data_205 : _GEN_4824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4826 = 8'hce == _match_key_qbytes_4_T ? phv_data_206 : _GEN_4825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4827 = 8'hcf == _match_key_qbytes_4_T ? phv_data_207 : _GEN_4826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4828 = 8'hd0 == _match_key_qbytes_4_T ? phv_data_208 : _GEN_4827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4829 = 8'hd1 == _match_key_qbytes_4_T ? phv_data_209 : _GEN_4828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4830 = 8'hd2 == _match_key_qbytes_4_T ? phv_data_210 : _GEN_4829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4831 = 8'hd3 == _match_key_qbytes_4_T ? phv_data_211 : _GEN_4830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4832 = 8'hd4 == _match_key_qbytes_4_T ? phv_data_212 : _GEN_4831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4833 = 8'hd5 == _match_key_qbytes_4_T ? phv_data_213 : _GEN_4832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4834 = 8'hd6 == _match_key_qbytes_4_T ? phv_data_214 : _GEN_4833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4835 = 8'hd7 == _match_key_qbytes_4_T ? phv_data_215 : _GEN_4834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4836 = 8'hd8 == _match_key_qbytes_4_T ? phv_data_216 : _GEN_4835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4837 = 8'hd9 == _match_key_qbytes_4_T ? phv_data_217 : _GEN_4836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4838 = 8'hda == _match_key_qbytes_4_T ? phv_data_218 : _GEN_4837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4839 = 8'hdb == _match_key_qbytes_4_T ? phv_data_219 : _GEN_4838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4840 = 8'hdc == _match_key_qbytes_4_T ? phv_data_220 : _GEN_4839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4841 = 8'hdd == _match_key_qbytes_4_T ? phv_data_221 : _GEN_4840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4842 = 8'hde == _match_key_qbytes_4_T ? phv_data_222 : _GEN_4841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4843 = 8'hdf == _match_key_qbytes_4_T ? phv_data_223 : _GEN_4842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4844 = 8'he0 == _match_key_qbytes_4_T ? phv_data_224 : _GEN_4843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4845 = 8'he1 == _match_key_qbytes_4_T ? phv_data_225 : _GEN_4844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4846 = 8'he2 == _match_key_qbytes_4_T ? phv_data_226 : _GEN_4845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4847 = 8'he3 == _match_key_qbytes_4_T ? phv_data_227 : _GEN_4846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4848 = 8'he4 == _match_key_qbytes_4_T ? phv_data_228 : _GEN_4847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4849 = 8'he5 == _match_key_qbytes_4_T ? phv_data_229 : _GEN_4848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4850 = 8'he6 == _match_key_qbytes_4_T ? phv_data_230 : _GEN_4849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4851 = 8'he7 == _match_key_qbytes_4_T ? phv_data_231 : _GEN_4850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4852 = 8'he8 == _match_key_qbytes_4_T ? phv_data_232 : _GEN_4851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4853 = 8'he9 == _match_key_qbytes_4_T ? phv_data_233 : _GEN_4852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4854 = 8'hea == _match_key_qbytes_4_T ? phv_data_234 : _GEN_4853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4855 = 8'heb == _match_key_qbytes_4_T ? phv_data_235 : _GEN_4854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4856 = 8'hec == _match_key_qbytes_4_T ? phv_data_236 : _GEN_4855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4857 = 8'hed == _match_key_qbytes_4_T ? phv_data_237 : _GEN_4856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4858 = 8'hee == _match_key_qbytes_4_T ? phv_data_238 : _GEN_4857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4859 = 8'hef == _match_key_qbytes_4_T ? phv_data_239 : _GEN_4858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4860 = 8'hf0 == _match_key_qbytes_4_T ? phv_data_240 : _GEN_4859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4861 = 8'hf1 == _match_key_qbytes_4_T ? phv_data_241 : _GEN_4860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4862 = 8'hf2 == _match_key_qbytes_4_T ? phv_data_242 : _GEN_4861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4863 = 8'hf3 == _match_key_qbytes_4_T ? phv_data_243 : _GEN_4862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4864 = 8'hf4 == _match_key_qbytes_4_T ? phv_data_244 : _GEN_4863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4865 = 8'hf5 == _match_key_qbytes_4_T ? phv_data_245 : _GEN_4864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4866 = 8'hf6 == _match_key_qbytes_4_T ? phv_data_246 : _GEN_4865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4867 = 8'hf7 == _match_key_qbytes_4_T ? phv_data_247 : _GEN_4866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4868 = 8'hf8 == _match_key_qbytes_4_T ? phv_data_248 : _GEN_4867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4869 = 8'hf9 == _match_key_qbytes_4_T ? phv_data_249 : _GEN_4868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4870 = 8'hfa == _match_key_qbytes_4_T ? phv_data_250 : _GEN_4869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4871 = 8'hfb == _match_key_qbytes_4_T ? phv_data_251 : _GEN_4870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4872 = 8'hfc == _match_key_qbytes_4_T ? phv_data_252 : _GEN_4871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4873 = 8'hfd == _match_key_qbytes_4_T ? phv_data_253 : _GEN_4872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4874 = 8'hfe == _match_key_qbytes_4_T ? phv_data_254 : _GEN_4873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4875 = 8'hff == _match_key_qbytes_4_T ? phv_data_255 : _GEN_4874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4877 = 8'h1 == _match_key_qbytes_4_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4878 = 8'h2 == _match_key_qbytes_4_T_1 ? phv_data_2 : _GEN_4877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4879 = 8'h3 == _match_key_qbytes_4_T_1 ? phv_data_3 : _GEN_4878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4880 = 8'h4 == _match_key_qbytes_4_T_1 ? phv_data_4 : _GEN_4879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4881 = 8'h5 == _match_key_qbytes_4_T_1 ? phv_data_5 : _GEN_4880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4882 = 8'h6 == _match_key_qbytes_4_T_1 ? phv_data_6 : _GEN_4881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4883 = 8'h7 == _match_key_qbytes_4_T_1 ? phv_data_7 : _GEN_4882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4884 = 8'h8 == _match_key_qbytes_4_T_1 ? phv_data_8 : _GEN_4883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4885 = 8'h9 == _match_key_qbytes_4_T_1 ? phv_data_9 : _GEN_4884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4886 = 8'ha == _match_key_qbytes_4_T_1 ? phv_data_10 : _GEN_4885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4887 = 8'hb == _match_key_qbytes_4_T_1 ? phv_data_11 : _GEN_4886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4888 = 8'hc == _match_key_qbytes_4_T_1 ? phv_data_12 : _GEN_4887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4889 = 8'hd == _match_key_qbytes_4_T_1 ? phv_data_13 : _GEN_4888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4890 = 8'he == _match_key_qbytes_4_T_1 ? phv_data_14 : _GEN_4889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4891 = 8'hf == _match_key_qbytes_4_T_1 ? phv_data_15 : _GEN_4890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4892 = 8'h10 == _match_key_qbytes_4_T_1 ? phv_data_16 : _GEN_4891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4893 = 8'h11 == _match_key_qbytes_4_T_1 ? phv_data_17 : _GEN_4892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4894 = 8'h12 == _match_key_qbytes_4_T_1 ? phv_data_18 : _GEN_4893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4895 = 8'h13 == _match_key_qbytes_4_T_1 ? phv_data_19 : _GEN_4894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4896 = 8'h14 == _match_key_qbytes_4_T_1 ? phv_data_20 : _GEN_4895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4897 = 8'h15 == _match_key_qbytes_4_T_1 ? phv_data_21 : _GEN_4896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4898 = 8'h16 == _match_key_qbytes_4_T_1 ? phv_data_22 : _GEN_4897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4899 = 8'h17 == _match_key_qbytes_4_T_1 ? phv_data_23 : _GEN_4898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4900 = 8'h18 == _match_key_qbytes_4_T_1 ? phv_data_24 : _GEN_4899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4901 = 8'h19 == _match_key_qbytes_4_T_1 ? phv_data_25 : _GEN_4900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4902 = 8'h1a == _match_key_qbytes_4_T_1 ? phv_data_26 : _GEN_4901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4903 = 8'h1b == _match_key_qbytes_4_T_1 ? phv_data_27 : _GEN_4902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4904 = 8'h1c == _match_key_qbytes_4_T_1 ? phv_data_28 : _GEN_4903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4905 = 8'h1d == _match_key_qbytes_4_T_1 ? phv_data_29 : _GEN_4904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4906 = 8'h1e == _match_key_qbytes_4_T_1 ? phv_data_30 : _GEN_4905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4907 = 8'h1f == _match_key_qbytes_4_T_1 ? phv_data_31 : _GEN_4906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4908 = 8'h20 == _match_key_qbytes_4_T_1 ? phv_data_32 : _GEN_4907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4909 = 8'h21 == _match_key_qbytes_4_T_1 ? phv_data_33 : _GEN_4908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4910 = 8'h22 == _match_key_qbytes_4_T_1 ? phv_data_34 : _GEN_4909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4911 = 8'h23 == _match_key_qbytes_4_T_1 ? phv_data_35 : _GEN_4910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4912 = 8'h24 == _match_key_qbytes_4_T_1 ? phv_data_36 : _GEN_4911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4913 = 8'h25 == _match_key_qbytes_4_T_1 ? phv_data_37 : _GEN_4912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4914 = 8'h26 == _match_key_qbytes_4_T_1 ? phv_data_38 : _GEN_4913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4915 = 8'h27 == _match_key_qbytes_4_T_1 ? phv_data_39 : _GEN_4914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4916 = 8'h28 == _match_key_qbytes_4_T_1 ? phv_data_40 : _GEN_4915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4917 = 8'h29 == _match_key_qbytes_4_T_1 ? phv_data_41 : _GEN_4916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4918 = 8'h2a == _match_key_qbytes_4_T_1 ? phv_data_42 : _GEN_4917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4919 = 8'h2b == _match_key_qbytes_4_T_1 ? phv_data_43 : _GEN_4918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4920 = 8'h2c == _match_key_qbytes_4_T_1 ? phv_data_44 : _GEN_4919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4921 = 8'h2d == _match_key_qbytes_4_T_1 ? phv_data_45 : _GEN_4920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4922 = 8'h2e == _match_key_qbytes_4_T_1 ? phv_data_46 : _GEN_4921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4923 = 8'h2f == _match_key_qbytes_4_T_1 ? phv_data_47 : _GEN_4922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4924 = 8'h30 == _match_key_qbytes_4_T_1 ? phv_data_48 : _GEN_4923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4925 = 8'h31 == _match_key_qbytes_4_T_1 ? phv_data_49 : _GEN_4924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4926 = 8'h32 == _match_key_qbytes_4_T_1 ? phv_data_50 : _GEN_4925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4927 = 8'h33 == _match_key_qbytes_4_T_1 ? phv_data_51 : _GEN_4926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4928 = 8'h34 == _match_key_qbytes_4_T_1 ? phv_data_52 : _GEN_4927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4929 = 8'h35 == _match_key_qbytes_4_T_1 ? phv_data_53 : _GEN_4928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4930 = 8'h36 == _match_key_qbytes_4_T_1 ? phv_data_54 : _GEN_4929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4931 = 8'h37 == _match_key_qbytes_4_T_1 ? phv_data_55 : _GEN_4930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4932 = 8'h38 == _match_key_qbytes_4_T_1 ? phv_data_56 : _GEN_4931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4933 = 8'h39 == _match_key_qbytes_4_T_1 ? phv_data_57 : _GEN_4932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4934 = 8'h3a == _match_key_qbytes_4_T_1 ? phv_data_58 : _GEN_4933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4935 = 8'h3b == _match_key_qbytes_4_T_1 ? phv_data_59 : _GEN_4934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4936 = 8'h3c == _match_key_qbytes_4_T_1 ? phv_data_60 : _GEN_4935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4937 = 8'h3d == _match_key_qbytes_4_T_1 ? phv_data_61 : _GEN_4936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4938 = 8'h3e == _match_key_qbytes_4_T_1 ? phv_data_62 : _GEN_4937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4939 = 8'h3f == _match_key_qbytes_4_T_1 ? phv_data_63 : _GEN_4938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4940 = 8'h40 == _match_key_qbytes_4_T_1 ? phv_data_64 : _GEN_4939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4941 = 8'h41 == _match_key_qbytes_4_T_1 ? phv_data_65 : _GEN_4940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4942 = 8'h42 == _match_key_qbytes_4_T_1 ? phv_data_66 : _GEN_4941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4943 = 8'h43 == _match_key_qbytes_4_T_1 ? phv_data_67 : _GEN_4942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4944 = 8'h44 == _match_key_qbytes_4_T_1 ? phv_data_68 : _GEN_4943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4945 = 8'h45 == _match_key_qbytes_4_T_1 ? phv_data_69 : _GEN_4944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4946 = 8'h46 == _match_key_qbytes_4_T_1 ? phv_data_70 : _GEN_4945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4947 = 8'h47 == _match_key_qbytes_4_T_1 ? phv_data_71 : _GEN_4946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4948 = 8'h48 == _match_key_qbytes_4_T_1 ? phv_data_72 : _GEN_4947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4949 = 8'h49 == _match_key_qbytes_4_T_1 ? phv_data_73 : _GEN_4948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4950 = 8'h4a == _match_key_qbytes_4_T_1 ? phv_data_74 : _GEN_4949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4951 = 8'h4b == _match_key_qbytes_4_T_1 ? phv_data_75 : _GEN_4950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4952 = 8'h4c == _match_key_qbytes_4_T_1 ? phv_data_76 : _GEN_4951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4953 = 8'h4d == _match_key_qbytes_4_T_1 ? phv_data_77 : _GEN_4952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4954 = 8'h4e == _match_key_qbytes_4_T_1 ? phv_data_78 : _GEN_4953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4955 = 8'h4f == _match_key_qbytes_4_T_1 ? phv_data_79 : _GEN_4954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4956 = 8'h50 == _match_key_qbytes_4_T_1 ? phv_data_80 : _GEN_4955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4957 = 8'h51 == _match_key_qbytes_4_T_1 ? phv_data_81 : _GEN_4956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4958 = 8'h52 == _match_key_qbytes_4_T_1 ? phv_data_82 : _GEN_4957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4959 = 8'h53 == _match_key_qbytes_4_T_1 ? phv_data_83 : _GEN_4958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4960 = 8'h54 == _match_key_qbytes_4_T_1 ? phv_data_84 : _GEN_4959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4961 = 8'h55 == _match_key_qbytes_4_T_1 ? phv_data_85 : _GEN_4960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4962 = 8'h56 == _match_key_qbytes_4_T_1 ? phv_data_86 : _GEN_4961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4963 = 8'h57 == _match_key_qbytes_4_T_1 ? phv_data_87 : _GEN_4962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4964 = 8'h58 == _match_key_qbytes_4_T_1 ? phv_data_88 : _GEN_4963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4965 = 8'h59 == _match_key_qbytes_4_T_1 ? phv_data_89 : _GEN_4964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4966 = 8'h5a == _match_key_qbytes_4_T_1 ? phv_data_90 : _GEN_4965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4967 = 8'h5b == _match_key_qbytes_4_T_1 ? phv_data_91 : _GEN_4966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4968 = 8'h5c == _match_key_qbytes_4_T_1 ? phv_data_92 : _GEN_4967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4969 = 8'h5d == _match_key_qbytes_4_T_1 ? phv_data_93 : _GEN_4968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4970 = 8'h5e == _match_key_qbytes_4_T_1 ? phv_data_94 : _GEN_4969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4971 = 8'h5f == _match_key_qbytes_4_T_1 ? phv_data_95 : _GEN_4970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4972 = 8'h60 == _match_key_qbytes_4_T_1 ? phv_data_96 : _GEN_4971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4973 = 8'h61 == _match_key_qbytes_4_T_1 ? phv_data_97 : _GEN_4972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4974 = 8'h62 == _match_key_qbytes_4_T_1 ? phv_data_98 : _GEN_4973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4975 = 8'h63 == _match_key_qbytes_4_T_1 ? phv_data_99 : _GEN_4974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4976 = 8'h64 == _match_key_qbytes_4_T_1 ? phv_data_100 : _GEN_4975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4977 = 8'h65 == _match_key_qbytes_4_T_1 ? phv_data_101 : _GEN_4976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4978 = 8'h66 == _match_key_qbytes_4_T_1 ? phv_data_102 : _GEN_4977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4979 = 8'h67 == _match_key_qbytes_4_T_1 ? phv_data_103 : _GEN_4978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4980 = 8'h68 == _match_key_qbytes_4_T_1 ? phv_data_104 : _GEN_4979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4981 = 8'h69 == _match_key_qbytes_4_T_1 ? phv_data_105 : _GEN_4980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4982 = 8'h6a == _match_key_qbytes_4_T_1 ? phv_data_106 : _GEN_4981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4983 = 8'h6b == _match_key_qbytes_4_T_1 ? phv_data_107 : _GEN_4982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4984 = 8'h6c == _match_key_qbytes_4_T_1 ? phv_data_108 : _GEN_4983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4985 = 8'h6d == _match_key_qbytes_4_T_1 ? phv_data_109 : _GEN_4984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4986 = 8'h6e == _match_key_qbytes_4_T_1 ? phv_data_110 : _GEN_4985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4987 = 8'h6f == _match_key_qbytes_4_T_1 ? phv_data_111 : _GEN_4986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4988 = 8'h70 == _match_key_qbytes_4_T_1 ? phv_data_112 : _GEN_4987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4989 = 8'h71 == _match_key_qbytes_4_T_1 ? phv_data_113 : _GEN_4988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4990 = 8'h72 == _match_key_qbytes_4_T_1 ? phv_data_114 : _GEN_4989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4991 = 8'h73 == _match_key_qbytes_4_T_1 ? phv_data_115 : _GEN_4990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4992 = 8'h74 == _match_key_qbytes_4_T_1 ? phv_data_116 : _GEN_4991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4993 = 8'h75 == _match_key_qbytes_4_T_1 ? phv_data_117 : _GEN_4992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4994 = 8'h76 == _match_key_qbytes_4_T_1 ? phv_data_118 : _GEN_4993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4995 = 8'h77 == _match_key_qbytes_4_T_1 ? phv_data_119 : _GEN_4994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4996 = 8'h78 == _match_key_qbytes_4_T_1 ? phv_data_120 : _GEN_4995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4997 = 8'h79 == _match_key_qbytes_4_T_1 ? phv_data_121 : _GEN_4996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4998 = 8'h7a == _match_key_qbytes_4_T_1 ? phv_data_122 : _GEN_4997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4999 = 8'h7b == _match_key_qbytes_4_T_1 ? phv_data_123 : _GEN_4998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5000 = 8'h7c == _match_key_qbytes_4_T_1 ? phv_data_124 : _GEN_4999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5001 = 8'h7d == _match_key_qbytes_4_T_1 ? phv_data_125 : _GEN_5000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5002 = 8'h7e == _match_key_qbytes_4_T_1 ? phv_data_126 : _GEN_5001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5003 = 8'h7f == _match_key_qbytes_4_T_1 ? phv_data_127 : _GEN_5002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5004 = 8'h80 == _match_key_qbytes_4_T_1 ? phv_data_128 : _GEN_5003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5005 = 8'h81 == _match_key_qbytes_4_T_1 ? phv_data_129 : _GEN_5004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5006 = 8'h82 == _match_key_qbytes_4_T_1 ? phv_data_130 : _GEN_5005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5007 = 8'h83 == _match_key_qbytes_4_T_1 ? phv_data_131 : _GEN_5006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5008 = 8'h84 == _match_key_qbytes_4_T_1 ? phv_data_132 : _GEN_5007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5009 = 8'h85 == _match_key_qbytes_4_T_1 ? phv_data_133 : _GEN_5008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5010 = 8'h86 == _match_key_qbytes_4_T_1 ? phv_data_134 : _GEN_5009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5011 = 8'h87 == _match_key_qbytes_4_T_1 ? phv_data_135 : _GEN_5010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5012 = 8'h88 == _match_key_qbytes_4_T_1 ? phv_data_136 : _GEN_5011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5013 = 8'h89 == _match_key_qbytes_4_T_1 ? phv_data_137 : _GEN_5012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5014 = 8'h8a == _match_key_qbytes_4_T_1 ? phv_data_138 : _GEN_5013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5015 = 8'h8b == _match_key_qbytes_4_T_1 ? phv_data_139 : _GEN_5014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5016 = 8'h8c == _match_key_qbytes_4_T_1 ? phv_data_140 : _GEN_5015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5017 = 8'h8d == _match_key_qbytes_4_T_1 ? phv_data_141 : _GEN_5016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5018 = 8'h8e == _match_key_qbytes_4_T_1 ? phv_data_142 : _GEN_5017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5019 = 8'h8f == _match_key_qbytes_4_T_1 ? phv_data_143 : _GEN_5018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5020 = 8'h90 == _match_key_qbytes_4_T_1 ? phv_data_144 : _GEN_5019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5021 = 8'h91 == _match_key_qbytes_4_T_1 ? phv_data_145 : _GEN_5020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5022 = 8'h92 == _match_key_qbytes_4_T_1 ? phv_data_146 : _GEN_5021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5023 = 8'h93 == _match_key_qbytes_4_T_1 ? phv_data_147 : _GEN_5022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5024 = 8'h94 == _match_key_qbytes_4_T_1 ? phv_data_148 : _GEN_5023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5025 = 8'h95 == _match_key_qbytes_4_T_1 ? phv_data_149 : _GEN_5024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5026 = 8'h96 == _match_key_qbytes_4_T_1 ? phv_data_150 : _GEN_5025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5027 = 8'h97 == _match_key_qbytes_4_T_1 ? phv_data_151 : _GEN_5026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5028 = 8'h98 == _match_key_qbytes_4_T_1 ? phv_data_152 : _GEN_5027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5029 = 8'h99 == _match_key_qbytes_4_T_1 ? phv_data_153 : _GEN_5028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5030 = 8'h9a == _match_key_qbytes_4_T_1 ? phv_data_154 : _GEN_5029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5031 = 8'h9b == _match_key_qbytes_4_T_1 ? phv_data_155 : _GEN_5030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5032 = 8'h9c == _match_key_qbytes_4_T_1 ? phv_data_156 : _GEN_5031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5033 = 8'h9d == _match_key_qbytes_4_T_1 ? phv_data_157 : _GEN_5032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5034 = 8'h9e == _match_key_qbytes_4_T_1 ? phv_data_158 : _GEN_5033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5035 = 8'h9f == _match_key_qbytes_4_T_1 ? phv_data_159 : _GEN_5034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5036 = 8'ha0 == _match_key_qbytes_4_T_1 ? phv_data_160 : _GEN_5035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5037 = 8'ha1 == _match_key_qbytes_4_T_1 ? phv_data_161 : _GEN_5036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5038 = 8'ha2 == _match_key_qbytes_4_T_1 ? phv_data_162 : _GEN_5037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5039 = 8'ha3 == _match_key_qbytes_4_T_1 ? phv_data_163 : _GEN_5038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5040 = 8'ha4 == _match_key_qbytes_4_T_1 ? phv_data_164 : _GEN_5039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5041 = 8'ha5 == _match_key_qbytes_4_T_1 ? phv_data_165 : _GEN_5040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5042 = 8'ha6 == _match_key_qbytes_4_T_1 ? phv_data_166 : _GEN_5041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5043 = 8'ha7 == _match_key_qbytes_4_T_1 ? phv_data_167 : _GEN_5042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5044 = 8'ha8 == _match_key_qbytes_4_T_1 ? phv_data_168 : _GEN_5043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5045 = 8'ha9 == _match_key_qbytes_4_T_1 ? phv_data_169 : _GEN_5044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5046 = 8'haa == _match_key_qbytes_4_T_1 ? phv_data_170 : _GEN_5045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5047 = 8'hab == _match_key_qbytes_4_T_1 ? phv_data_171 : _GEN_5046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5048 = 8'hac == _match_key_qbytes_4_T_1 ? phv_data_172 : _GEN_5047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5049 = 8'had == _match_key_qbytes_4_T_1 ? phv_data_173 : _GEN_5048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5050 = 8'hae == _match_key_qbytes_4_T_1 ? phv_data_174 : _GEN_5049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5051 = 8'haf == _match_key_qbytes_4_T_1 ? phv_data_175 : _GEN_5050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5052 = 8'hb0 == _match_key_qbytes_4_T_1 ? phv_data_176 : _GEN_5051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5053 = 8'hb1 == _match_key_qbytes_4_T_1 ? phv_data_177 : _GEN_5052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5054 = 8'hb2 == _match_key_qbytes_4_T_1 ? phv_data_178 : _GEN_5053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5055 = 8'hb3 == _match_key_qbytes_4_T_1 ? phv_data_179 : _GEN_5054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5056 = 8'hb4 == _match_key_qbytes_4_T_1 ? phv_data_180 : _GEN_5055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5057 = 8'hb5 == _match_key_qbytes_4_T_1 ? phv_data_181 : _GEN_5056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5058 = 8'hb6 == _match_key_qbytes_4_T_1 ? phv_data_182 : _GEN_5057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5059 = 8'hb7 == _match_key_qbytes_4_T_1 ? phv_data_183 : _GEN_5058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5060 = 8'hb8 == _match_key_qbytes_4_T_1 ? phv_data_184 : _GEN_5059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5061 = 8'hb9 == _match_key_qbytes_4_T_1 ? phv_data_185 : _GEN_5060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5062 = 8'hba == _match_key_qbytes_4_T_1 ? phv_data_186 : _GEN_5061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5063 = 8'hbb == _match_key_qbytes_4_T_1 ? phv_data_187 : _GEN_5062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5064 = 8'hbc == _match_key_qbytes_4_T_1 ? phv_data_188 : _GEN_5063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5065 = 8'hbd == _match_key_qbytes_4_T_1 ? phv_data_189 : _GEN_5064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5066 = 8'hbe == _match_key_qbytes_4_T_1 ? phv_data_190 : _GEN_5065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5067 = 8'hbf == _match_key_qbytes_4_T_1 ? phv_data_191 : _GEN_5066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5068 = 8'hc0 == _match_key_qbytes_4_T_1 ? phv_data_192 : _GEN_5067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5069 = 8'hc1 == _match_key_qbytes_4_T_1 ? phv_data_193 : _GEN_5068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5070 = 8'hc2 == _match_key_qbytes_4_T_1 ? phv_data_194 : _GEN_5069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5071 = 8'hc3 == _match_key_qbytes_4_T_1 ? phv_data_195 : _GEN_5070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5072 = 8'hc4 == _match_key_qbytes_4_T_1 ? phv_data_196 : _GEN_5071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5073 = 8'hc5 == _match_key_qbytes_4_T_1 ? phv_data_197 : _GEN_5072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5074 = 8'hc6 == _match_key_qbytes_4_T_1 ? phv_data_198 : _GEN_5073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5075 = 8'hc7 == _match_key_qbytes_4_T_1 ? phv_data_199 : _GEN_5074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5076 = 8'hc8 == _match_key_qbytes_4_T_1 ? phv_data_200 : _GEN_5075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5077 = 8'hc9 == _match_key_qbytes_4_T_1 ? phv_data_201 : _GEN_5076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5078 = 8'hca == _match_key_qbytes_4_T_1 ? phv_data_202 : _GEN_5077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5079 = 8'hcb == _match_key_qbytes_4_T_1 ? phv_data_203 : _GEN_5078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5080 = 8'hcc == _match_key_qbytes_4_T_1 ? phv_data_204 : _GEN_5079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5081 = 8'hcd == _match_key_qbytes_4_T_1 ? phv_data_205 : _GEN_5080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5082 = 8'hce == _match_key_qbytes_4_T_1 ? phv_data_206 : _GEN_5081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5083 = 8'hcf == _match_key_qbytes_4_T_1 ? phv_data_207 : _GEN_5082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5084 = 8'hd0 == _match_key_qbytes_4_T_1 ? phv_data_208 : _GEN_5083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5085 = 8'hd1 == _match_key_qbytes_4_T_1 ? phv_data_209 : _GEN_5084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5086 = 8'hd2 == _match_key_qbytes_4_T_1 ? phv_data_210 : _GEN_5085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5087 = 8'hd3 == _match_key_qbytes_4_T_1 ? phv_data_211 : _GEN_5086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5088 = 8'hd4 == _match_key_qbytes_4_T_1 ? phv_data_212 : _GEN_5087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5089 = 8'hd5 == _match_key_qbytes_4_T_1 ? phv_data_213 : _GEN_5088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5090 = 8'hd6 == _match_key_qbytes_4_T_1 ? phv_data_214 : _GEN_5089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5091 = 8'hd7 == _match_key_qbytes_4_T_1 ? phv_data_215 : _GEN_5090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5092 = 8'hd8 == _match_key_qbytes_4_T_1 ? phv_data_216 : _GEN_5091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5093 = 8'hd9 == _match_key_qbytes_4_T_1 ? phv_data_217 : _GEN_5092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5094 = 8'hda == _match_key_qbytes_4_T_1 ? phv_data_218 : _GEN_5093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5095 = 8'hdb == _match_key_qbytes_4_T_1 ? phv_data_219 : _GEN_5094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5096 = 8'hdc == _match_key_qbytes_4_T_1 ? phv_data_220 : _GEN_5095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5097 = 8'hdd == _match_key_qbytes_4_T_1 ? phv_data_221 : _GEN_5096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5098 = 8'hde == _match_key_qbytes_4_T_1 ? phv_data_222 : _GEN_5097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5099 = 8'hdf == _match_key_qbytes_4_T_1 ? phv_data_223 : _GEN_5098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5100 = 8'he0 == _match_key_qbytes_4_T_1 ? phv_data_224 : _GEN_5099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5101 = 8'he1 == _match_key_qbytes_4_T_1 ? phv_data_225 : _GEN_5100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5102 = 8'he2 == _match_key_qbytes_4_T_1 ? phv_data_226 : _GEN_5101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5103 = 8'he3 == _match_key_qbytes_4_T_1 ? phv_data_227 : _GEN_5102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5104 = 8'he4 == _match_key_qbytes_4_T_1 ? phv_data_228 : _GEN_5103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5105 = 8'he5 == _match_key_qbytes_4_T_1 ? phv_data_229 : _GEN_5104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5106 = 8'he6 == _match_key_qbytes_4_T_1 ? phv_data_230 : _GEN_5105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5107 = 8'he7 == _match_key_qbytes_4_T_1 ? phv_data_231 : _GEN_5106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5108 = 8'he8 == _match_key_qbytes_4_T_1 ? phv_data_232 : _GEN_5107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5109 = 8'he9 == _match_key_qbytes_4_T_1 ? phv_data_233 : _GEN_5108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5110 = 8'hea == _match_key_qbytes_4_T_1 ? phv_data_234 : _GEN_5109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5111 = 8'heb == _match_key_qbytes_4_T_1 ? phv_data_235 : _GEN_5110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5112 = 8'hec == _match_key_qbytes_4_T_1 ? phv_data_236 : _GEN_5111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5113 = 8'hed == _match_key_qbytes_4_T_1 ? phv_data_237 : _GEN_5112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5114 = 8'hee == _match_key_qbytes_4_T_1 ? phv_data_238 : _GEN_5113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5115 = 8'hef == _match_key_qbytes_4_T_1 ? phv_data_239 : _GEN_5114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5116 = 8'hf0 == _match_key_qbytes_4_T_1 ? phv_data_240 : _GEN_5115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5117 = 8'hf1 == _match_key_qbytes_4_T_1 ? phv_data_241 : _GEN_5116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5118 = 8'hf2 == _match_key_qbytes_4_T_1 ? phv_data_242 : _GEN_5117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5119 = 8'hf3 == _match_key_qbytes_4_T_1 ? phv_data_243 : _GEN_5118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5120 = 8'hf4 == _match_key_qbytes_4_T_1 ? phv_data_244 : _GEN_5119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5121 = 8'hf5 == _match_key_qbytes_4_T_1 ? phv_data_245 : _GEN_5120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5122 = 8'hf6 == _match_key_qbytes_4_T_1 ? phv_data_246 : _GEN_5121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5123 = 8'hf7 == _match_key_qbytes_4_T_1 ? phv_data_247 : _GEN_5122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5124 = 8'hf8 == _match_key_qbytes_4_T_1 ? phv_data_248 : _GEN_5123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5125 = 8'hf9 == _match_key_qbytes_4_T_1 ? phv_data_249 : _GEN_5124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5126 = 8'hfa == _match_key_qbytes_4_T_1 ? phv_data_250 : _GEN_5125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5127 = 8'hfb == _match_key_qbytes_4_T_1 ? phv_data_251 : _GEN_5126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5128 = 8'hfc == _match_key_qbytes_4_T_1 ? phv_data_252 : _GEN_5127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5129 = 8'hfd == _match_key_qbytes_4_T_1 ? phv_data_253 : _GEN_5128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5130 = 8'hfe == _match_key_qbytes_4_T_1 ? phv_data_254 : _GEN_5129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5131 = 8'hff == _match_key_qbytes_4_T_1 ? phv_data_255 : _GEN_5130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_4_T_3 = {_GEN_4875,_GEN_5131,_GEN_4363,_GEN_4619}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_4 = local_offset_4 < end_offset ? _match_key_qbytes_4_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_5 = 8'h14 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_5_hi = local_offset_5[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_5_T = {match_key_qbytes_5_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_5_T_1 = {match_key_qbytes_5_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_5_T_2 = {match_key_qbytes_5_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_5134 = 8'h1 == _match_key_qbytes_5_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5135 = 8'h2 == _match_key_qbytes_5_T_2 ? phv_data_2 : _GEN_5134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5136 = 8'h3 == _match_key_qbytes_5_T_2 ? phv_data_3 : _GEN_5135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5137 = 8'h4 == _match_key_qbytes_5_T_2 ? phv_data_4 : _GEN_5136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5138 = 8'h5 == _match_key_qbytes_5_T_2 ? phv_data_5 : _GEN_5137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5139 = 8'h6 == _match_key_qbytes_5_T_2 ? phv_data_6 : _GEN_5138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5140 = 8'h7 == _match_key_qbytes_5_T_2 ? phv_data_7 : _GEN_5139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5141 = 8'h8 == _match_key_qbytes_5_T_2 ? phv_data_8 : _GEN_5140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5142 = 8'h9 == _match_key_qbytes_5_T_2 ? phv_data_9 : _GEN_5141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5143 = 8'ha == _match_key_qbytes_5_T_2 ? phv_data_10 : _GEN_5142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5144 = 8'hb == _match_key_qbytes_5_T_2 ? phv_data_11 : _GEN_5143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5145 = 8'hc == _match_key_qbytes_5_T_2 ? phv_data_12 : _GEN_5144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5146 = 8'hd == _match_key_qbytes_5_T_2 ? phv_data_13 : _GEN_5145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5147 = 8'he == _match_key_qbytes_5_T_2 ? phv_data_14 : _GEN_5146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5148 = 8'hf == _match_key_qbytes_5_T_2 ? phv_data_15 : _GEN_5147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5149 = 8'h10 == _match_key_qbytes_5_T_2 ? phv_data_16 : _GEN_5148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5150 = 8'h11 == _match_key_qbytes_5_T_2 ? phv_data_17 : _GEN_5149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5151 = 8'h12 == _match_key_qbytes_5_T_2 ? phv_data_18 : _GEN_5150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5152 = 8'h13 == _match_key_qbytes_5_T_2 ? phv_data_19 : _GEN_5151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5153 = 8'h14 == _match_key_qbytes_5_T_2 ? phv_data_20 : _GEN_5152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5154 = 8'h15 == _match_key_qbytes_5_T_2 ? phv_data_21 : _GEN_5153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5155 = 8'h16 == _match_key_qbytes_5_T_2 ? phv_data_22 : _GEN_5154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5156 = 8'h17 == _match_key_qbytes_5_T_2 ? phv_data_23 : _GEN_5155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5157 = 8'h18 == _match_key_qbytes_5_T_2 ? phv_data_24 : _GEN_5156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5158 = 8'h19 == _match_key_qbytes_5_T_2 ? phv_data_25 : _GEN_5157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5159 = 8'h1a == _match_key_qbytes_5_T_2 ? phv_data_26 : _GEN_5158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5160 = 8'h1b == _match_key_qbytes_5_T_2 ? phv_data_27 : _GEN_5159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5161 = 8'h1c == _match_key_qbytes_5_T_2 ? phv_data_28 : _GEN_5160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5162 = 8'h1d == _match_key_qbytes_5_T_2 ? phv_data_29 : _GEN_5161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5163 = 8'h1e == _match_key_qbytes_5_T_2 ? phv_data_30 : _GEN_5162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5164 = 8'h1f == _match_key_qbytes_5_T_2 ? phv_data_31 : _GEN_5163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5165 = 8'h20 == _match_key_qbytes_5_T_2 ? phv_data_32 : _GEN_5164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5166 = 8'h21 == _match_key_qbytes_5_T_2 ? phv_data_33 : _GEN_5165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5167 = 8'h22 == _match_key_qbytes_5_T_2 ? phv_data_34 : _GEN_5166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5168 = 8'h23 == _match_key_qbytes_5_T_2 ? phv_data_35 : _GEN_5167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5169 = 8'h24 == _match_key_qbytes_5_T_2 ? phv_data_36 : _GEN_5168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5170 = 8'h25 == _match_key_qbytes_5_T_2 ? phv_data_37 : _GEN_5169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5171 = 8'h26 == _match_key_qbytes_5_T_2 ? phv_data_38 : _GEN_5170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5172 = 8'h27 == _match_key_qbytes_5_T_2 ? phv_data_39 : _GEN_5171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5173 = 8'h28 == _match_key_qbytes_5_T_2 ? phv_data_40 : _GEN_5172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5174 = 8'h29 == _match_key_qbytes_5_T_2 ? phv_data_41 : _GEN_5173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5175 = 8'h2a == _match_key_qbytes_5_T_2 ? phv_data_42 : _GEN_5174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5176 = 8'h2b == _match_key_qbytes_5_T_2 ? phv_data_43 : _GEN_5175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5177 = 8'h2c == _match_key_qbytes_5_T_2 ? phv_data_44 : _GEN_5176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5178 = 8'h2d == _match_key_qbytes_5_T_2 ? phv_data_45 : _GEN_5177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5179 = 8'h2e == _match_key_qbytes_5_T_2 ? phv_data_46 : _GEN_5178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5180 = 8'h2f == _match_key_qbytes_5_T_2 ? phv_data_47 : _GEN_5179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5181 = 8'h30 == _match_key_qbytes_5_T_2 ? phv_data_48 : _GEN_5180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5182 = 8'h31 == _match_key_qbytes_5_T_2 ? phv_data_49 : _GEN_5181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5183 = 8'h32 == _match_key_qbytes_5_T_2 ? phv_data_50 : _GEN_5182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5184 = 8'h33 == _match_key_qbytes_5_T_2 ? phv_data_51 : _GEN_5183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5185 = 8'h34 == _match_key_qbytes_5_T_2 ? phv_data_52 : _GEN_5184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5186 = 8'h35 == _match_key_qbytes_5_T_2 ? phv_data_53 : _GEN_5185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5187 = 8'h36 == _match_key_qbytes_5_T_2 ? phv_data_54 : _GEN_5186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5188 = 8'h37 == _match_key_qbytes_5_T_2 ? phv_data_55 : _GEN_5187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5189 = 8'h38 == _match_key_qbytes_5_T_2 ? phv_data_56 : _GEN_5188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5190 = 8'h39 == _match_key_qbytes_5_T_2 ? phv_data_57 : _GEN_5189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5191 = 8'h3a == _match_key_qbytes_5_T_2 ? phv_data_58 : _GEN_5190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5192 = 8'h3b == _match_key_qbytes_5_T_2 ? phv_data_59 : _GEN_5191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5193 = 8'h3c == _match_key_qbytes_5_T_2 ? phv_data_60 : _GEN_5192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5194 = 8'h3d == _match_key_qbytes_5_T_2 ? phv_data_61 : _GEN_5193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5195 = 8'h3e == _match_key_qbytes_5_T_2 ? phv_data_62 : _GEN_5194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5196 = 8'h3f == _match_key_qbytes_5_T_2 ? phv_data_63 : _GEN_5195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5197 = 8'h40 == _match_key_qbytes_5_T_2 ? phv_data_64 : _GEN_5196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5198 = 8'h41 == _match_key_qbytes_5_T_2 ? phv_data_65 : _GEN_5197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5199 = 8'h42 == _match_key_qbytes_5_T_2 ? phv_data_66 : _GEN_5198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5200 = 8'h43 == _match_key_qbytes_5_T_2 ? phv_data_67 : _GEN_5199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5201 = 8'h44 == _match_key_qbytes_5_T_2 ? phv_data_68 : _GEN_5200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5202 = 8'h45 == _match_key_qbytes_5_T_2 ? phv_data_69 : _GEN_5201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5203 = 8'h46 == _match_key_qbytes_5_T_2 ? phv_data_70 : _GEN_5202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5204 = 8'h47 == _match_key_qbytes_5_T_2 ? phv_data_71 : _GEN_5203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5205 = 8'h48 == _match_key_qbytes_5_T_2 ? phv_data_72 : _GEN_5204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5206 = 8'h49 == _match_key_qbytes_5_T_2 ? phv_data_73 : _GEN_5205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5207 = 8'h4a == _match_key_qbytes_5_T_2 ? phv_data_74 : _GEN_5206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5208 = 8'h4b == _match_key_qbytes_5_T_2 ? phv_data_75 : _GEN_5207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5209 = 8'h4c == _match_key_qbytes_5_T_2 ? phv_data_76 : _GEN_5208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5210 = 8'h4d == _match_key_qbytes_5_T_2 ? phv_data_77 : _GEN_5209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5211 = 8'h4e == _match_key_qbytes_5_T_2 ? phv_data_78 : _GEN_5210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5212 = 8'h4f == _match_key_qbytes_5_T_2 ? phv_data_79 : _GEN_5211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5213 = 8'h50 == _match_key_qbytes_5_T_2 ? phv_data_80 : _GEN_5212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5214 = 8'h51 == _match_key_qbytes_5_T_2 ? phv_data_81 : _GEN_5213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5215 = 8'h52 == _match_key_qbytes_5_T_2 ? phv_data_82 : _GEN_5214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5216 = 8'h53 == _match_key_qbytes_5_T_2 ? phv_data_83 : _GEN_5215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5217 = 8'h54 == _match_key_qbytes_5_T_2 ? phv_data_84 : _GEN_5216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5218 = 8'h55 == _match_key_qbytes_5_T_2 ? phv_data_85 : _GEN_5217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5219 = 8'h56 == _match_key_qbytes_5_T_2 ? phv_data_86 : _GEN_5218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5220 = 8'h57 == _match_key_qbytes_5_T_2 ? phv_data_87 : _GEN_5219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5221 = 8'h58 == _match_key_qbytes_5_T_2 ? phv_data_88 : _GEN_5220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5222 = 8'h59 == _match_key_qbytes_5_T_2 ? phv_data_89 : _GEN_5221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5223 = 8'h5a == _match_key_qbytes_5_T_2 ? phv_data_90 : _GEN_5222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5224 = 8'h5b == _match_key_qbytes_5_T_2 ? phv_data_91 : _GEN_5223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5225 = 8'h5c == _match_key_qbytes_5_T_2 ? phv_data_92 : _GEN_5224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5226 = 8'h5d == _match_key_qbytes_5_T_2 ? phv_data_93 : _GEN_5225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5227 = 8'h5e == _match_key_qbytes_5_T_2 ? phv_data_94 : _GEN_5226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5228 = 8'h5f == _match_key_qbytes_5_T_2 ? phv_data_95 : _GEN_5227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5229 = 8'h60 == _match_key_qbytes_5_T_2 ? phv_data_96 : _GEN_5228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5230 = 8'h61 == _match_key_qbytes_5_T_2 ? phv_data_97 : _GEN_5229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5231 = 8'h62 == _match_key_qbytes_5_T_2 ? phv_data_98 : _GEN_5230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5232 = 8'h63 == _match_key_qbytes_5_T_2 ? phv_data_99 : _GEN_5231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5233 = 8'h64 == _match_key_qbytes_5_T_2 ? phv_data_100 : _GEN_5232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5234 = 8'h65 == _match_key_qbytes_5_T_2 ? phv_data_101 : _GEN_5233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5235 = 8'h66 == _match_key_qbytes_5_T_2 ? phv_data_102 : _GEN_5234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5236 = 8'h67 == _match_key_qbytes_5_T_2 ? phv_data_103 : _GEN_5235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5237 = 8'h68 == _match_key_qbytes_5_T_2 ? phv_data_104 : _GEN_5236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5238 = 8'h69 == _match_key_qbytes_5_T_2 ? phv_data_105 : _GEN_5237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5239 = 8'h6a == _match_key_qbytes_5_T_2 ? phv_data_106 : _GEN_5238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5240 = 8'h6b == _match_key_qbytes_5_T_2 ? phv_data_107 : _GEN_5239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5241 = 8'h6c == _match_key_qbytes_5_T_2 ? phv_data_108 : _GEN_5240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5242 = 8'h6d == _match_key_qbytes_5_T_2 ? phv_data_109 : _GEN_5241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5243 = 8'h6e == _match_key_qbytes_5_T_2 ? phv_data_110 : _GEN_5242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5244 = 8'h6f == _match_key_qbytes_5_T_2 ? phv_data_111 : _GEN_5243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5245 = 8'h70 == _match_key_qbytes_5_T_2 ? phv_data_112 : _GEN_5244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5246 = 8'h71 == _match_key_qbytes_5_T_2 ? phv_data_113 : _GEN_5245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5247 = 8'h72 == _match_key_qbytes_5_T_2 ? phv_data_114 : _GEN_5246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5248 = 8'h73 == _match_key_qbytes_5_T_2 ? phv_data_115 : _GEN_5247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5249 = 8'h74 == _match_key_qbytes_5_T_2 ? phv_data_116 : _GEN_5248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5250 = 8'h75 == _match_key_qbytes_5_T_2 ? phv_data_117 : _GEN_5249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5251 = 8'h76 == _match_key_qbytes_5_T_2 ? phv_data_118 : _GEN_5250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5252 = 8'h77 == _match_key_qbytes_5_T_2 ? phv_data_119 : _GEN_5251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5253 = 8'h78 == _match_key_qbytes_5_T_2 ? phv_data_120 : _GEN_5252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5254 = 8'h79 == _match_key_qbytes_5_T_2 ? phv_data_121 : _GEN_5253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5255 = 8'h7a == _match_key_qbytes_5_T_2 ? phv_data_122 : _GEN_5254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5256 = 8'h7b == _match_key_qbytes_5_T_2 ? phv_data_123 : _GEN_5255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5257 = 8'h7c == _match_key_qbytes_5_T_2 ? phv_data_124 : _GEN_5256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5258 = 8'h7d == _match_key_qbytes_5_T_2 ? phv_data_125 : _GEN_5257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5259 = 8'h7e == _match_key_qbytes_5_T_2 ? phv_data_126 : _GEN_5258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5260 = 8'h7f == _match_key_qbytes_5_T_2 ? phv_data_127 : _GEN_5259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5261 = 8'h80 == _match_key_qbytes_5_T_2 ? phv_data_128 : _GEN_5260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5262 = 8'h81 == _match_key_qbytes_5_T_2 ? phv_data_129 : _GEN_5261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5263 = 8'h82 == _match_key_qbytes_5_T_2 ? phv_data_130 : _GEN_5262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5264 = 8'h83 == _match_key_qbytes_5_T_2 ? phv_data_131 : _GEN_5263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5265 = 8'h84 == _match_key_qbytes_5_T_2 ? phv_data_132 : _GEN_5264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5266 = 8'h85 == _match_key_qbytes_5_T_2 ? phv_data_133 : _GEN_5265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5267 = 8'h86 == _match_key_qbytes_5_T_2 ? phv_data_134 : _GEN_5266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5268 = 8'h87 == _match_key_qbytes_5_T_2 ? phv_data_135 : _GEN_5267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5269 = 8'h88 == _match_key_qbytes_5_T_2 ? phv_data_136 : _GEN_5268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5270 = 8'h89 == _match_key_qbytes_5_T_2 ? phv_data_137 : _GEN_5269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5271 = 8'h8a == _match_key_qbytes_5_T_2 ? phv_data_138 : _GEN_5270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5272 = 8'h8b == _match_key_qbytes_5_T_2 ? phv_data_139 : _GEN_5271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5273 = 8'h8c == _match_key_qbytes_5_T_2 ? phv_data_140 : _GEN_5272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5274 = 8'h8d == _match_key_qbytes_5_T_2 ? phv_data_141 : _GEN_5273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5275 = 8'h8e == _match_key_qbytes_5_T_2 ? phv_data_142 : _GEN_5274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5276 = 8'h8f == _match_key_qbytes_5_T_2 ? phv_data_143 : _GEN_5275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5277 = 8'h90 == _match_key_qbytes_5_T_2 ? phv_data_144 : _GEN_5276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5278 = 8'h91 == _match_key_qbytes_5_T_2 ? phv_data_145 : _GEN_5277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5279 = 8'h92 == _match_key_qbytes_5_T_2 ? phv_data_146 : _GEN_5278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5280 = 8'h93 == _match_key_qbytes_5_T_2 ? phv_data_147 : _GEN_5279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5281 = 8'h94 == _match_key_qbytes_5_T_2 ? phv_data_148 : _GEN_5280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5282 = 8'h95 == _match_key_qbytes_5_T_2 ? phv_data_149 : _GEN_5281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5283 = 8'h96 == _match_key_qbytes_5_T_2 ? phv_data_150 : _GEN_5282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5284 = 8'h97 == _match_key_qbytes_5_T_2 ? phv_data_151 : _GEN_5283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5285 = 8'h98 == _match_key_qbytes_5_T_2 ? phv_data_152 : _GEN_5284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5286 = 8'h99 == _match_key_qbytes_5_T_2 ? phv_data_153 : _GEN_5285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5287 = 8'h9a == _match_key_qbytes_5_T_2 ? phv_data_154 : _GEN_5286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5288 = 8'h9b == _match_key_qbytes_5_T_2 ? phv_data_155 : _GEN_5287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5289 = 8'h9c == _match_key_qbytes_5_T_2 ? phv_data_156 : _GEN_5288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5290 = 8'h9d == _match_key_qbytes_5_T_2 ? phv_data_157 : _GEN_5289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5291 = 8'h9e == _match_key_qbytes_5_T_2 ? phv_data_158 : _GEN_5290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5292 = 8'h9f == _match_key_qbytes_5_T_2 ? phv_data_159 : _GEN_5291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5293 = 8'ha0 == _match_key_qbytes_5_T_2 ? phv_data_160 : _GEN_5292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5294 = 8'ha1 == _match_key_qbytes_5_T_2 ? phv_data_161 : _GEN_5293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5295 = 8'ha2 == _match_key_qbytes_5_T_2 ? phv_data_162 : _GEN_5294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5296 = 8'ha3 == _match_key_qbytes_5_T_2 ? phv_data_163 : _GEN_5295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5297 = 8'ha4 == _match_key_qbytes_5_T_2 ? phv_data_164 : _GEN_5296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5298 = 8'ha5 == _match_key_qbytes_5_T_2 ? phv_data_165 : _GEN_5297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5299 = 8'ha6 == _match_key_qbytes_5_T_2 ? phv_data_166 : _GEN_5298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5300 = 8'ha7 == _match_key_qbytes_5_T_2 ? phv_data_167 : _GEN_5299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5301 = 8'ha8 == _match_key_qbytes_5_T_2 ? phv_data_168 : _GEN_5300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5302 = 8'ha9 == _match_key_qbytes_5_T_2 ? phv_data_169 : _GEN_5301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5303 = 8'haa == _match_key_qbytes_5_T_2 ? phv_data_170 : _GEN_5302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5304 = 8'hab == _match_key_qbytes_5_T_2 ? phv_data_171 : _GEN_5303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5305 = 8'hac == _match_key_qbytes_5_T_2 ? phv_data_172 : _GEN_5304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5306 = 8'had == _match_key_qbytes_5_T_2 ? phv_data_173 : _GEN_5305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5307 = 8'hae == _match_key_qbytes_5_T_2 ? phv_data_174 : _GEN_5306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5308 = 8'haf == _match_key_qbytes_5_T_2 ? phv_data_175 : _GEN_5307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5309 = 8'hb0 == _match_key_qbytes_5_T_2 ? phv_data_176 : _GEN_5308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5310 = 8'hb1 == _match_key_qbytes_5_T_2 ? phv_data_177 : _GEN_5309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5311 = 8'hb2 == _match_key_qbytes_5_T_2 ? phv_data_178 : _GEN_5310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5312 = 8'hb3 == _match_key_qbytes_5_T_2 ? phv_data_179 : _GEN_5311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5313 = 8'hb4 == _match_key_qbytes_5_T_2 ? phv_data_180 : _GEN_5312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5314 = 8'hb5 == _match_key_qbytes_5_T_2 ? phv_data_181 : _GEN_5313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5315 = 8'hb6 == _match_key_qbytes_5_T_2 ? phv_data_182 : _GEN_5314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5316 = 8'hb7 == _match_key_qbytes_5_T_2 ? phv_data_183 : _GEN_5315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5317 = 8'hb8 == _match_key_qbytes_5_T_2 ? phv_data_184 : _GEN_5316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5318 = 8'hb9 == _match_key_qbytes_5_T_2 ? phv_data_185 : _GEN_5317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5319 = 8'hba == _match_key_qbytes_5_T_2 ? phv_data_186 : _GEN_5318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5320 = 8'hbb == _match_key_qbytes_5_T_2 ? phv_data_187 : _GEN_5319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5321 = 8'hbc == _match_key_qbytes_5_T_2 ? phv_data_188 : _GEN_5320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5322 = 8'hbd == _match_key_qbytes_5_T_2 ? phv_data_189 : _GEN_5321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5323 = 8'hbe == _match_key_qbytes_5_T_2 ? phv_data_190 : _GEN_5322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5324 = 8'hbf == _match_key_qbytes_5_T_2 ? phv_data_191 : _GEN_5323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5325 = 8'hc0 == _match_key_qbytes_5_T_2 ? phv_data_192 : _GEN_5324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5326 = 8'hc1 == _match_key_qbytes_5_T_2 ? phv_data_193 : _GEN_5325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5327 = 8'hc2 == _match_key_qbytes_5_T_2 ? phv_data_194 : _GEN_5326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5328 = 8'hc3 == _match_key_qbytes_5_T_2 ? phv_data_195 : _GEN_5327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5329 = 8'hc4 == _match_key_qbytes_5_T_2 ? phv_data_196 : _GEN_5328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5330 = 8'hc5 == _match_key_qbytes_5_T_2 ? phv_data_197 : _GEN_5329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5331 = 8'hc6 == _match_key_qbytes_5_T_2 ? phv_data_198 : _GEN_5330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5332 = 8'hc7 == _match_key_qbytes_5_T_2 ? phv_data_199 : _GEN_5331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5333 = 8'hc8 == _match_key_qbytes_5_T_2 ? phv_data_200 : _GEN_5332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5334 = 8'hc9 == _match_key_qbytes_5_T_2 ? phv_data_201 : _GEN_5333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5335 = 8'hca == _match_key_qbytes_5_T_2 ? phv_data_202 : _GEN_5334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5336 = 8'hcb == _match_key_qbytes_5_T_2 ? phv_data_203 : _GEN_5335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5337 = 8'hcc == _match_key_qbytes_5_T_2 ? phv_data_204 : _GEN_5336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5338 = 8'hcd == _match_key_qbytes_5_T_2 ? phv_data_205 : _GEN_5337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5339 = 8'hce == _match_key_qbytes_5_T_2 ? phv_data_206 : _GEN_5338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5340 = 8'hcf == _match_key_qbytes_5_T_2 ? phv_data_207 : _GEN_5339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5341 = 8'hd0 == _match_key_qbytes_5_T_2 ? phv_data_208 : _GEN_5340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5342 = 8'hd1 == _match_key_qbytes_5_T_2 ? phv_data_209 : _GEN_5341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5343 = 8'hd2 == _match_key_qbytes_5_T_2 ? phv_data_210 : _GEN_5342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5344 = 8'hd3 == _match_key_qbytes_5_T_2 ? phv_data_211 : _GEN_5343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5345 = 8'hd4 == _match_key_qbytes_5_T_2 ? phv_data_212 : _GEN_5344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5346 = 8'hd5 == _match_key_qbytes_5_T_2 ? phv_data_213 : _GEN_5345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5347 = 8'hd6 == _match_key_qbytes_5_T_2 ? phv_data_214 : _GEN_5346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5348 = 8'hd7 == _match_key_qbytes_5_T_2 ? phv_data_215 : _GEN_5347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5349 = 8'hd8 == _match_key_qbytes_5_T_2 ? phv_data_216 : _GEN_5348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5350 = 8'hd9 == _match_key_qbytes_5_T_2 ? phv_data_217 : _GEN_5349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5351 = 8'hda == _match_key_qbytes_5_T_2 ? phv_data_218 : _GEN_5350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5352 = 8'hdb == _match_key_qbytes_5_T_2 ? phv_data_219 : _GEN_5351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5353 = 8'hdc == _match_key_qbytes_5_T_2 ? phv_data_220 : _GEN_5352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5354 = 8'hdd == _match_key_qbytes_5_T_2 ? phv_data_221 : _GEN_5353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5355 = 8'hde == _match_key_qbytes_5_T_2 ? phv_data_222 : _GEN_5354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5356 = 8'hdf == _match_key_qbytes_5_T_2 ? phv_data_223 : _GEN_5355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5357 = 8'he0 == _match_key_qbytes_5_T_2 ? phv_data_224 : _GEN_5356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5358 = 8'he1 == _match_key_qbytes_5_T_2 ? phv_data_225 : _GEN_5357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5359 = 8'he2 == _match_key_qbytes_5_T_2 ? phv_data_226 : _GEN_5358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5360 = 8'he3 == _match_key_qbytes_5_T_2 ? phv_data_227 : _GEN_5359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5361 = 8'he4 == _match_key_qbytes_5_T_2 ? phv_data_228 : _GEN_5360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5362 = 8'he5 == _match_key_qbytes_5_T_2 ? phv_data_229 : _GEN_5361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5363 = 8'he6 == _match_key_qbytes_5_T_2 ? phv_data_230 : _GEN_5362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5364 = 8'he7 == _match_key_qbytes_5_T_2 ? phv_data_231 : _GEN_5363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5365 = 8'he8 == _match_key_qbytes_5_T_2 ? phv_data_232 : _GEN_5364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5366 = 8'he9 == _match_key_qbytes_5_T_2 ? phv_data_233 : _GEN_5365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5367 = 8'hea == _match_key_qbytes_5_T_2 ? phv_data_234 : _GEN_5366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5368 = 8'heb == _match_key_qbytes_5_T_2 ? phv_data_235 : _GEN_5367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5369 = 8'hec == _match_key_qbytes_5_T_2 ? phv_data_236 : _GEN_5368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5370 = 8'hed == _match_key_qbytes_5_T_2 ? phv_data_237 : _GEN_5369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5371 = 8'hee == _match_key_qbytes_5_T_2 ? phv_data_238 : _GEN_5370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5372 = 8'hef == _match_key_qbytes_5_T_2 ? phv_data_239 : _GEN_5371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5373 = 8'hf0 == _match_key_qbytes_5_T_2 ? phv_data_240 : _GEN_5372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5374 = 8'hf1 == _match_key_qbytes_5_T_2 ? phv_data_241 : _GEN_5373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5375 = 8'hf2 == _match_key_qbytes_5_T_2 ? phv_data_242 : _GEN_5374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5376 = 8'hf3 == _match_key_qbytes_5_T_2 ? phv_data_243 : _GEN_5375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5377 = 8'hf4 == _match_key_qbytes_5_T_2 ? phv_data_244 : _GEN_5376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5378 = 8'hf5 == _match_key_qbytes_5_T_2 ? phv_data_245 : _GEN_5377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5379 = 8'hf6 == _match_key_qbytes_5_T_2 ? phv_data_246 : _GEN_5378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5380 = 8'hf7 == _match_key_qbytes_5_T_2 ? phv_data_247 : _GEN_5379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5381 = 8'hf8 == _match_key_qbytes_5_T_2 ? phv_data_248 : _GEN_5380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5382 = 8'hf9 == _match_key_qbytes_5_T_2 ? phv_data_249 : _GEN_5381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5383 = 8'hfa == _match_key_qbytes_5_T_2 ? phv_data_250 : _GEN_5382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5384 = 8'hfb == _match_key_qbytes_5_T_2 ? phv_data_251 : _GEN_5383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5385 = 8'hfc == _match_key_qbytes_5_T_2 ? phv_data_252 : _GEN_5384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5386 = 8'hfd == _match_key_qbytes_5_T_2 ? phv_data_253 : _GEN_5385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5387 = 8'hfe == _match_key_qbytes_5_T_2 ? phv_data_254 : _GEN_5386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5388 = 8'hff == _match_key_qbytes_5_T_2 ? phv_data_255 : _GEN_5387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5390 = 8'h1 == local_offset_5 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5391 = 8'h2 == local_offset_5 ? phv_data_2 : _GEN_5390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5392 = 8'h3 == local_offset_5 ? phv_data_3 : _GEN_5391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5393 = 8'h4 == local_offset_5 ? phv_data_4 : _GEN_5392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5394 = 8'h5 == local_offset_5 ? phv_data_5 : _GEN_5393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5395 = 8'h6 == local_offset_5 ? phv_data_6 : _GEN_5394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5396 = 8'h7 == local_offset_5 ? phv_data_7 : _GEN_5395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5397 = 8'h8 == local_offset_5 ? phv_data_8 : _GEN_5396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5398 = 8'h9 == local_offset_5 ? phv_data_9 : _GEN_5397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5399 = 8'ha == local_offset_5 ? phv_data_10 : _GEN_5398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5400 = 8'hb == local_offset_5 ? phv_data_11 : _GEN_5399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5401 = 8'hc == local_offset_5 ? phv_data_12 : _GEN_5400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5402 = 8'hd == local_offset_5 ? phv_data_13 : _GEN_5401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5403 = 8'he == local_offset_5 ? phv_data_14 : _GEN_5402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5404 = 8'hf == local_offset_5 ? phv_data_15 : _GEN_5403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5405 = 8'h10 == local_offset_5 ? phv_data_16 : _GEN_5404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5406 = 8'h11 == local_offset_5 ? phv_data_17 : _GEN_5405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5407 = 8'h12 == local_offset_5 ? phv_data_18 : _GEN_5406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5408 = 8'h13 == local_offset_5 ? phv_data_19 : _GEN_5407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5409 = 8'h14 == local_offset_5 ? phv_data_20 : _GEN_5408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5410 = 8'h15 == local_offset_5 ? phv_data_21 : _GEN_5409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5411 = 8'h16 == local_offset_5 ? phv_data_22 : _GEN_5410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5412 = 8'h17 == local_offset_5 ? phv_data_23 : _GEN_5411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5413 = 8'h18 == local_offset_5 ? phv_data_24 : _GEN_5412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5414 = 8'h19 == local_offset_5 ? phv_data_25 : _GEN_5413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5415 = 8'h1a == local_offset_5 ? phv_data_26 : _GEN_5414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5416 = 8'h1b == local_offset_5 ? phv_data_27 : _GEN_5415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5417 = 8'h1c == local_offset_5 ? phv_data_28 : _GEN_5416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5418 = 8'h1d == local_offset_5 ? phv_data_29 : _GEN_5417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5419 = 8'h1e == local_offset_5 ? phv_data_30 : _GEN_5418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5420 = 8'h1f == local_offset_5 ? phv_data_31 : _GEN_5419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5421 = 8'h20 == local_offset_5 ? phv_data_32 : _GEN_5420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5422 = 8'h21 == local_offset_5 ? phv_data_33 : _GEN_5421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5423 = 8'h22 == local_offset_5 ? phv_data_34 : _GEN_5422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5424 = 8'h23 == local_offset_5 ? phv_data_35 : _GEN_5423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5425 = 8'h24 == local_offset_5 ? phv_data_36 : _GEN_5424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5426 = 8'h25 == local_offset_5 ? phv_data_37 : _GEN_5425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5427 = 8'h26 == local_offset_5 ? phv_data_38 : _GEN_5426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5428 = 8'h27 == local_offset_5 ? phv_data_39 : _GEN_5427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5429 = 8'h28 == local_offset_5 ? phv_data_40 : _GEN_5428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5430 = 8'h29 == local_offset_5 ? phv_data_41 : _GEN_5429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5431 = 8'h2a == local_offset_5 ? phv_data_42 : _GEN_5430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5432 = 8'h2b == local_offset_5 ? phv_data_43 : _GEN_5431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5433 = 8'h2c == local_offset_5 ? phv_data_44 : _GEN_5432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5434 = 8'h2d == local_offset_5 ? phv_data_45 : _GEN_5433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5435 = 8'h2e == local_offset_5 ? phv_data_46 : _GEN_5434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5436 = 8'h2f == local_offset_5 ? phv_data_47 : _GEN_5435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5437 = 8'h30 == local_offset_5 ? phv_data_48 : _GEN_5436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5438 = 8'h31 == local_offset_5 ? phv_data_49 : _GEN_5437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5439 = 8'h32 == local_offset_5 ? phv_data_50 : _GEN_5438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5440 = 8'h33 == local_offset_5 ? phv_data_51 : _GEN_5439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5441 = 8'h34 == local_offset_5 ? phv_data_52 : _GEN_5440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5442 = 8'h35 == local_offset_5 ? phv_data_53 : _GEN_5441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5443 = 8'h36 == local_offset_5 ? phv_data_54 : _GEN_5442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5444 = 8'h37 == local_offset_5 ? phv_data_55 : _GEN_5443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5445 = 8'h38 == local_offset_5 ? phv_data_56 : _GEN_5444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5446 = 8'h39 == local_offset_5 ? phv_data_57 : _GEN_5445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5447 = 8'h3a == local_offset_5 ? phv_data_58 : _GEN_5446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5448 = 8'h3b == local_offset_5 ? phv_data_59 : _GEN_5447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5449 = 8'h3c == local_offset_5 ? phv_data_60 : _GEN_5448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5450 = 8'h3d == local_offset_5 ? phv_data_61 : _GEN_5449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5451 = 8'h3e == local_offset_5 ? phv_data_62 : _GEN_5450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5452 = 8'h3f == local_offset_5 ? phv_data_63 : _GEN_5451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5453 = 8'h40 == local_offset_5 ? phv_data_64 : _GEN_5452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5454 = 8'h41 == local_offset_5 ? phv_data_65 : _GEN_5453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5455 = 8'h42 == local_offset_5 ? phv_data_66 : _GEN_5454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5456 = 8'h43 == local_offset_5 ? phv_data_67 : _GEN_5455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5457 = 8'h44 == local_offset_5 ? phv_data_68 : _GEN_5456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5458 = 8'h45 == local_offset_5 ? phv_data_69 : _GEN_5457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5459 = 8'h46 == local_offset_5 ? phv_data_70 : _GEN_5458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5460 = 8'h47 == local_offset_5 ? phv_data_71 : _GEN_5459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5461 = 8'h48 == local_offset_5 ? phv_data_72 : _GEN_5460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5462 = 8'h49 == local_offset_5 ? phv_data_73 : _GEN_5461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5463 = 8'h4a == local_offset_5 ? phv_data_74 : _GEN_5462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5464 = 8'h4b == local_offset_5 ? phv_data_75 : _GEN_5463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5465 = 8'h4c == local_offset_5 ? phv_data_76 : _GEN_5464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5466 = 8'h4d == local_offset_5 ? phv_data_77 : _GEN_5465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5467 = 8'h4e == local_offset_5 ? phv_data_78 : _GEN_5466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5468 = 8'h4f == local_offset_5 ? phv_data_79 : _GEN_5467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5469 = 8'h50 == local_offset_5 ? phv_data_80 : _GEN_5468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5470 = 8'h51 == local_offset_5 ? phv_data_81 : _GEN_5469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5471 = 8'h52 == local_offset_5 ? phv_data_82 : _GEN_5470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5472 = 8'h53 == local_offset_5 ? phv_data_83 : _GEN_5471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5473 = 8'h54 == local_offset_5 ? phv_data_84 : _GEN_5472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5474 = 8'h55 == local_offset_5 ? phv_data_85 : _GEN_5473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5475 = 8'h56 == local_offset_5 ? phv_data_86 : _GEN_5474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5476 = 8'h57 == local_offset_5 ? phv_data_87 : _GEN_5475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5477 = 8'h58 == local_offset_5 ? phv_data_88 : _GEN_5476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5478 = 8'h59 == local_offset_5 ? phv_data_89 : _GEN_5477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5479 = 8'h5a == local_offset_5 ? phv_data_90 : _GEN_5478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5480 = 8'h5b == local_offset_5 ? phv_data_91 : _GEN_5479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5481 = 8'h5c == local_offset_5 ? phv_data_92 : _GEN_5480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5482 = 8'h5d == local_offset_5 ? phv_data_93 : _GEN_5481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5483 = 8'h5e == local_offset_5 ? phv_data_94 : _GEN_5482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5484 = 8'h5f == local_offset_5 ? phv_data_95 : _GEN_5483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5485 = 8'h60 == local_offset_5 ? phv_data_96 : _GEN_5484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5486 = 8'h61 == local_offset_5 ? phv_data_97 : _GEN_5485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5487 = 8'h62 == local_offset_5 ? phv_data_98 : _GEN_5486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5488 = 8'h63 == local_offset_5 ? phv_data_99 : _GEN_5487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5489 = 8'h64 == local_offset_5 ? phv_data_100 : _GEN_5488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5490 = 8'h65 == local_offset_5 ? phv_data_101 : _GEN_5489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5491 = 8'h66 == local_offset_5 ? phv_data_102 : _GEN_5490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5492 = 8'h67 == local_offset_5 ? phv_data_103 : _GEN_5491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5493 = 8'h68 == local_offset_5 ? phv_data_104 : _GEN_5492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5494 = 8'h69 == local_offset_5 ? phv_data_105 : _GEN_5493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5495 = 8'h6a == local_offset_5 ? phv_data_106 : _GEN_5494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5496 = 8'h6b == local_offset_5 ? phv_data_107 : _GEN_5495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5497 = 8'h6c == local_offset_5 ? phv_data_108 : _GEN_5496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5498 = 8'h6d == local_offset_5 ? phv_data_109 : _GEN_5497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5499 = 8'h6e == local_offset_5 ? phv_data_110 : _GEN_5498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5500 = 8'h6f == local_offset_5 ? phv_data_111 : _GEN_5499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5501 = 8'h70 == local_offset_5 ? phv_data_112 : _GEN_5500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5502 = 8'h71 == local_offset_5 ? phv_data_113 : _GEN_5501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5503 = 8'h72 == local_offset_5 ? phv_data_114 : _GEN_5502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5504 = 8'h73 == local_offset_5 ? phv_data_115 : _GEN_5503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5505 = 8'h74 == local_offset_5 ? phv_data_116 : _GEN_5504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5506 = 8'h75 == local_offset_5 ? phv_data_117 : _GEN_5505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5507 = 8'h76 == local_offset_5 ? phv_data_118 : _GEN_5506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5508 = 8'h77 == local_offset_5 ? phv_data_119 : _GEN_5507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5509 = 8'h78 == local_offset_5 ? phv_data_120 : _GEN_5508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5510 = 8'h79 == local_offset_5 ? phv_data_121 : _GEN_5509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5511 = 8'h7a == local_offset_5 ? phv_data_122 : _GEN_5510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5512 = 8'h7b == local_offset_5 ? phv_data_123 : _GEN_5511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5513 = 8'h7c == local_offset_5 ? phv_data_124 : _GEN_5512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5514 = 8'h7d == local_offset_5 ? phv_data_125 : _GEN_5513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5515 = 8'h7e == local_offset_5 ? phv_data_126 : _GEN_5514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5516 = 8'h7f == local_offset_5 ? phv_data_127 : _GEN_5515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5517 = 8'h80 == local_offset_5 ? phv_data_128 : _GEN_5516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5518 = 8'h81 == local_offset_5 ? phv_data_129 : _GEN_5517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5519 = 8'h82 == local_offset_5 ? phv_data_130 : _GEN_5518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5520 = 8'h83 == local_offset_5 ? phv_data_131 : _GEN_5519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5521 = 8'h84 == local_offset_5 ? phv_data_132 : _GEN_5520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5522 = 8'h85 == local_offset_5 ? phv_data_133 : _GEN_5521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5523 = 8'h86 == local_offset_5 ? phv_data_134 : _GEN_5522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5524 = 8'h87 == local_offset_5 ? phv_data_135 : _GEN_5523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5525 = 8'h88 == local_offset_5 ? phv_data_136 : _GEN_5524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5526 = 8'h89 == local_offset_5 ? phv_data_137 : _GEN_5525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5527 = 8'h8a == local_offset_5 ? phv_data_138 : _GEN_5526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5528 = 8'h8b == local_offset_5 ? phv_data_139 : _GEN_5527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5529 = 8'h8c == local_offset_5 ? phv_data_140 : _GEN_5528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5530 = 8'h8d == local_offset_5 ? phv_data_141 : _GEN_5529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5531 = 8'h8e == local_offset_5 ? phv_data_142 : _GEN_5530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5532 = 8'h8f == local_offset_5 ? phv_data_143 : _GEN_5531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5533 = 8'h90 == local_offset_5 ? phv_data_144 : _GEN_5532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5534 = 8'h91 == local_offset_5 ? phv_data_145 : _GEN_5533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5535 = 8'h92 == local_offset_5 ? phv_data_146 : _GEN_5534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5536 = 8'h93 == local_offset_5 ? phv_data_147 : _GEN_5535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5537 = 8'h94 == local_offset_5 ? phv_data_148 : _GEN_5536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5538 = 8'h95 == local_offset_5 ? phv_data_149 : _GEN_5537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5539 = 8'h96 == local_offset_5 ? phv_data_150 : _GEN_5538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5540 = 8'h97 == local_offset_5 ? phv_data_151 : _GEN_5539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5541 = 8'h98 == local_offset_5 ? phv_data_152 : _GEN_5540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5542 = 8'h99 == local_offset_5 ? phv_data_153 : _GEN_5541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5543 = 8'h9a == local_offset_5 ? phv_data_154 : _GEN_5542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5544 = 8'h9b == local_offset_5 ? phv_data_155 : _GEN_5543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5545 = 8'h9c == local_offset_5 ? phv_data_156 : _GEN_5544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5546 = 8'h9d == local_offset_5 ? phv_data_157 : _GEN_5545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5547 = 8'h9e == local_offset_5 ? phv_data_158 : _GEN_5546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5548 = 8'h9f == local_offset_5 ? phv_data_159 : _GEN_5547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5549 = 8'ha0 == local_offset_5 ? phv_data_160 : _GEN_5548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5550 = 8'ha1 == local_offset_5 ? phv_data_161 : _GEN_5549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5551 = 8'ha2 == local_offset_5 ? phv_data_162 : _GEN_5550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5552 = 8'ha3 == local_offset_5 ? phv_data_163 : _GEN_5551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5553 = 8'ha4 == local_offset_5 ? phv_data_164 : _GEN_5552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5554 = 8'ha5 == local_offset_5 ? phv_data_165 : _GEN_5553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5555 = 8'ha6 == local_offset_5 ? phv_data_166 : _GEN_5554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5556 = 8'ha7 == local_offset_5 ? phv_data_167 : _GEN_5555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5557 = 8'ha8 == local_offset_5 ? phv_data_168 : _GEN_5556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5558 = 8'ha9 == local_offset_5 ? phv_data_169 : _GEN_5557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5559 = 8'haa == local_offset_5 ? phv_data_170 : _GEN_5558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5560 = 8'hab == local_offset_5 ? phv_data_171 : _GEN_5559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5561 = 8'hac == local_offset_5 ? phv_data_172 : _GEN_5560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5562 = 8'had == local_offset_5 ? phv_data_173 : _GEN_5561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5563 = 8'hae == local_offset_5 ? phv_data_174 : _GEN_5562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5564 = 8'haf == local_offset_5 ? phv_data_175 : _GEN_5563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5565 = 8'hb0 == local_offset_5 ? phv_data_176 : _GEN_5564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5566 = 8'hb1 == local_offset_5 ? phv_data_177 : _GEN_5565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5567 = 8'hb2 == local_offset_5 ? phv_data_178 : _GEN_5566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5568 = 8'hb3 == local_offset_5 ? phv_data_179 : _GEN_5567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5569 = 8'hb4 == local_offset_5 ? phv_data_180 : _GEN_5568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5570 = 8'hb5 == local_offset_5 ? phv_data_181 : _GEN_5569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5571 = 8'hb6 == local_offset_5 ? phv_data_182 : _GEN_5570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5572 = 8'hb7 == local_offset_5 ? phv_data_183 : _GEN_5571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5573 = 8'hb8 == local_offset_5 ? phv_data_184 : _GEN_5572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5574 = 8'hb9 == local_offset_5 ? phv_data_185 : _GEN_5573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5575 = 8'hba == local_offset_5 ? phv_data_186 : _GEN_5574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5576 = 8'hbb == local_offset_5 ? phv_data_187 : _GEN_5575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5577 = 8'hbc == local_offset_5 ? phv_data_188 : _GEN_5576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5578 = 8'hbd == local_offset_5 ? phv_data_189 : _GEN_5577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5579 = 8'hbe == local_offset_5 ? phv_data_190 : _GEN_5578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5580 = 8'hbf == local_offset_5 ? phv_data_191 : _GEN_5579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5581 = 8'hc0 == local_offset_5 ? phv_data_192 : _GEN_5580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5582 = 8'hc1 == local_offset_5 ? phv_data_193 : _GEN_5581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5583 = 8'hc2 == local_offset_5 ? phv_data_194 : _GEN_5582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5584 = 8'hc3 == local_offset_5 ? phv_data_195 : _GEN_5583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5585 = 8'hc4 == local_offset_5 ? phv_data_196 : _GEN_5584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5586 = 8'hc5 == local_offset_5 ? phv_data_197 : _GEN_5585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5587 = 8'hc6 == local_offset_5 ? phv_data_198 : _GEN_5586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5588 = 8'hc7 == local_offset_5 ? phv_data_199 : _GEN_5587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5589 = 8'hc8 == local_offset_5 ? phv_data_200 : _GEN_5588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5590 = 8'hc9 == local_offset_5 ? phv_data_201 : _GEN_5589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5591 = 8'hca == local_offset_5 ? phv_data_202 : _GEN_5590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5592 = 8'hcb == local_offset_5 ? phv_data_203 : _GEN_5591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5593 = 8'hcc == local_offset_5 ? phv_data_204 : _GEN_5592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5594 = 8'hcd == local_offset_5 ? phv_data_205 : _GEN_5593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5595 = 8'hce == local_offset_5 ? phv_data_206 : _GEN_5594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5596 = 8'hcf == local_offset_5 ? phv_data_207 : _GEN_5595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5597 = 8'hd0 == local_offset_5 ? phv_data_208 : _GEN_5596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5598 = 8'hd1 == local_offset_5 ? phv_data_209 : _GEN_5597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5599 = 8'hd2 == local_offset_5 ? phv_data_210 : _GEN_5598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5600 = 8'hd3 == local_offset_5 ? phv_data_211 : _GEN_5599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5601 = 8'hd4 == local_offset_5 ? phv_data_212 : _GEN_5600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5602 = 8'hd5 == local_offset_5 ? phv_data_213 : _GEN_5601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5603 = 8'hd6 == local_offset_5 ? phv_data_214 : _GEN_5602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5604 = 8'hd7 == local_offset_5 ? phv_data_215 : _GEN_5603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5605 = 8'hd8 == local_offset_5 ? phv_data_216 : _GEN_5604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5606 = 8'hd9 == local_offset_5 ? phv_data_217 : _GEN_5605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5607 = 8'hda == local_offset_5 ? phv_data_218 : _GEN_5606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5608 = 8'hdb == local_offset_5 ? phv_data_219 : _GEN_5607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5609 = 8'hdc == local_offset_5 ? phv_data_220 : _GEN_5608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5610 = 8'hdd == local_offset_5 ? phv_data_221 : _GEN_5609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5611 = 8'hde == local_offset_5 ? phv_data_222 : _GEN_5610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5612 = 8'hdf == local_offset_5 ? phv_data_223 : _GEN_5611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5613 = 8'he0 == local_offset_5 ? phv_data_224 : _GEN_5612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5614 = 8'he1 == local_offset_5 ? phv_data_225 : _GEN_5613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5615 = 8'he2 == local_offset_5 ? phv_data_226 : _GEN_5614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5616 = 8'he3 == local_offset_5 ? phv_data_227 : _GEN_5615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5617 = 8'he4 == local_offset_5 ? phv_data_228 : _GEN_5616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5618 = 8'he5 == local_offset_5 ? phv_data_229 : _GEN_5617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5619 = 8'he6 == local_offset_5 ? phv_data_230 : _GEN_5618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5620 = 8'he7 == local_offset_5 ? phv_data_231 : _GEN_5619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5621 = 8'he8 == local_offset_5 ? phv_data_232 : _GEN_5620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5622 = 8'he9 == local_offset_5 ? phv_data_233 : _GEN_5621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5623 = 8'hea == local_offset_5 ? phv_data_234 : _GEN_5622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5624 = 8'heb == local_offset_5 ? phv_data_235 : _GEN_5623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5625 = 8'hec == local_offset_5 ? phv_data_236 : _GEN_5624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5626 = 8'hed == local_offset_5 ? phv_data_237 : _GEN_5625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5627 = 8'hee == local_offset_5 ? phv_data_238 : _GEN_5626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5628 = 8'hef == local_offset_5 ? phv_data_239 : _GEN_5627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5629 = 8'hf0 == local_offset_5 ? phv_data_240 : _GEN_5628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5630 = 8'hf1 == local_offset_5 ? phv_data_241 : _GEN_5629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5631 = 8'hf2 == local_offset_5 ? phv_data_242 : _GEN_5630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5632 = 8'hf3 == local_offset_5 ? phv_data_243 : _GEN_5631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5633 = 8'hf4 == local_offset_5 ? phv_data_244 : _GEN_5632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5634 = 8'hf5 == local_offset_5 ? phv_data_245 : _GEN_5633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5635 = 8'hf6 == local_offset_5 ? phv_data_246 : _GEN_5634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5636 = 8'hf7 == local_offset_5 ? phv_data_247 : _GEN_5635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5637 = 8'hf8 == local_offset_5 ? phv_data_248 : _GEN_5636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5638 = 8'hf9 == local_offset_5 ? phv_data_249 : _GEN_5637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5639 = 8'hfa == local_offset_5 ? phv_data_250 : _GEN_5638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5640 = 8'hfb == local_offset_5 ? phv_data_251 : _GEN_5639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5641 = 8'hfc == local_offset_5 ? phv_data_252 : _GEN_5640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5642 = 8'hfd == local_offset_5 ? phv_data_253 : _GEN_5641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5643 = 8'hfe == local_offset_5 ? phv_data_254 : _GEN_5642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5644 = 8'hff == local_offset_5 ? phv_data_255 : _GEN_5643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5646 = 8'h1 == _match_key_qbytes_5_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5647 = 8'h2 == _match_key_qbytes_5_T ? phv_data_2 : _GEN_5646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5648 = 8'h3 == _match_key_qbytes_5_T ? phv_data_3 : _GEN_5647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5649 = 8'h4 == _match_key_qbytes_5_T ? phv_data_4 : _GEN_5648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5650 = 8'h5 == _match_key_qbytes_5_T ? phv_data_5 : _GEN_5649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5651 = 8'h6 == _match_key_qbytes_5_T ? phv_data_6 : _GEN_5650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5652 = 8'h7 == _match_key_qbytes_5_T ? phv_data_7 : _GEN_5651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5653 = 8'h8 == _match_key_qbytes_5_T ? phv_data_8 : _GEN_5652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5654 = 8'h9 == _match_key_qbytes_5_T ? phv_data_9 : _GEN_5653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5655 = 8'ha == _match_key_qbytes_5_T ? phv_data_10 : _GEN_5654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5656 = 8'hb == _match_key_qbytes_5_T ? phv_data_11 : _GEN_5655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5657 = 8'hc == _match_key_qbytes_5_T ? phv_data_12 : _GEN_5656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5658 = 8'hd == _match_key_qbytes_5_T ? phv_data_13 : _GEN_5657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5659 = 8'he == _match_key_qbytes_5_T ? phv_data_14 : _GEN_5658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5660 = 8'hf == _match_key_qbytes_5_T ? phv_data_15 : _GEN_5659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5661 = 8'h10 == _match_key_qbytes_5_T ? phv_data_16 : _GEN_5660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5662 = 8'h11 == _match_key_qbytes_5_T ? phv_data_17 : _GEN_5661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5663 = 8'h12 == _match_key_qbytes_5_T ? phv_data_18 : _GEN_5662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5664 = 8'h13 == _match_key_qbytes_5_T ? phv_data_19 : _GEN_5663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5665 = 8'h14 == _match_key_qbytes_5_T ? phv_data_20 : _GEN_5664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5666 = 8'h15 == _match_key_qbytes_5_T ? phv_data_21 : _GEN_5665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5667 = 8'h16 == _match_key_qbytes_5_T ? phv_data_22 : _GEN_5666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5668 = 8'h17 == _match_key_qbytes_5_T ? phv_data_23 : _GEN_5667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5669 = 8'h18 == _match_key_qbytes_5_T ? phv_data_24 : _GEN_5668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5670 = 8'h19 == _match_key_qbytes_5_T ? phv_data_25 : _GEN_5669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5671 = 8'h1a == _match_key_qbytes_5_T ? phv_data_26 : _GEN_5670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5672 = 8'h1b == _match_key_qbytes_5_T ? phv_data_27 : _GEN_5671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5673 = 8'h1c == _match_key_qbytes_5_T ? phv_data_28 : _GEN_5672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5674 = 8'h1d == _match_key_qbytes_5_T ? phv_data_29 : _GEN_5673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5675 = 8'h1e == _match_key_qbytes_5_T ? phv_data_30 : _GEN_5674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5676 = 8'h1f == _match_key_qbytes_5_T ? phv_data_31 : _GEN_5675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5677 = 8'h20 == _match_key_qbytes_5_T ? phv_data_32 : _GEN_5676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5678 = 8'h21 == _match_key_qbytes_5_T ? phv_data_33 : _GEN_5677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5679 = 8'h22 == _match_key_qbytes_5_T ? phv_data_34 : _GEN_5678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5680 = 8'h23 == _match_key_qbytes_5_T ? phv_data_35 : _GEN_5679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5681 = 8'h24 == _match_key_qbytes_5_T ? phv_data_36 : _GEN_5680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5682 = 8'h25 == _match_key_qbytes_5_T ? phv_data_37 : _GEN_5681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5683 = 8'h26 == _match_key_qbytes_5_T ? phv_data_38 : _GEN_5682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5684 = 8'h27 == _match_key_qbytes_5_T ? phv_data_39 : _GEN_5683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5685 = 8'h28 == _match_key_qbytes_5_T ? phv_data_40 : _GEN_5684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5686 = 8'h29 == _match_key_qbytes_5_T ? phv_data_41 : _GEN_5685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5687 = 8'h2a == _match_key_qbytes_5_T ? phv_data_42 : _GEN_5686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5688 = 8'h2b == _match_key_qbytes_5_T ? phv_data_43 : _GEN_5687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5689 = 8'h2c == _match_key_qbytes_5_T ? phv_data_44 : _GEN_5688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5690 = 8'h2d == _match_key_qbytes_5_T ? phv_data_45 : _GEN_5689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5691 = 8'h2e == _match_key_qbytes_5_T ? phv_data_46 : _GEN_5690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5692 = 8'h2f == _match_key_qbytes_5_T ? phv_data_47 : _GEN_5691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5693 = 8'h30 == _match_key_qbytes_5_T ? phv_data_48 : _GEN_5692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5694 = 8'h31 == _match_key_qbytes_5_T ? phv_data_49 : _GEN_5693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5695 = 8'h32 == _match_key_qbytes_5_T ? phv_data_50 : _GEN_5694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5696 = 8'h33 == _match_key_qbytes_5_T ? phv_data_51 : _GEN_5695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5697 = 8'h34 == _match_key_qbytes_5_T ? phv_data_52 : _GEN_5696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5698 = 8'h35 == _match_key_qbytes_5_T ? phv_data_53 : _GEN_5697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5699 = 8'h36 == _match_key_qbytes_5_T ? phv_data_54 : _GEN_5698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5700 = 8'h37 == _match_key_qbytes_5_T ? phv_data_55 : _GEN_5699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5701 = 8'h38 == _match_key_qbytes_5_T ? phv_data_56 : _GEN_5700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5702 = 8'h39 == _match_key_qbytes_5_T ? phv_data_57 : _GEN_5701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5703 = 8'h3a == _match_key_qbytes_5_T ? phv_data_58 : _GEN_5702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5704 = 8'h3b == _match_key_qbytes_5_T ? phv_data_59 : _GEN_5703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5705 = 8'h3c == _match_key_qbytes_5_T ? phv_data_60 : _GEN_5704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5706 = 8'h3d == _match_key_qbytes_5_T ? phv_data_61 : _GEN_5705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5707 = 8'h3e == _match_key_qbytes_5_T ? phv_data_62 : _GEN_5706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5708 = 8'h3f == _match_key_qbytes_5_T ? phv_data_63 : _GEN_5707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5709 = 8'h40 == _match_key_qbytes_5_T ? phv_data_64 : _GEN_5708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5710 = 8'h41 == _match_key_qbytes_5_T ? phv_data_65 : _GEN_5709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5711 = 8'h42 == _match_key_qbytes_5_T ? phv_data_66 : _GEN_5710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5712 = 8'h43 == _match_key_qbytes_5_T ? phv_data_67 : _GEN_5711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5713 = 8'h44 == _match_key_qbytes_5_T ? phv_data_68 : _GEN_5712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5714 = 8'h45 == _match_key_qbytes_5_T ? phv_data_69 : _GEN_5713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5715 = 8'h46 == _match_key_qbytes_5_T ? phv_data_70 : _GEN_5714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5716 = 8'h47 == _match_key_qbytes_5_T ? phv_data_71 : _GEN_5715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5717 = 8'h48 == _match_key_qbytes_5_T ? phv_data_72 : _GEN_5716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5718 = 8'h49 == _match_key_qbytes_5_T ? phv_data_73 : _GEN_5717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5719 = 8'h4a == _match_key_qbytes_5_T ? phv_data_74 : _GEN_5718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5720 = 8'h4b == _match_key_qbytes_5_T ? phv_data_75 : _GEN_5719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5721 = 8'h4c == _match_key_qbytes_5_T ? phv_data_76 : _GEN_5720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5722 = 8'h4d == _match_key_qbytes_5_T ? phv_data_77 : _GEN_5721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5723 = 8'h4e == _match_key_qbytes_5_T ? phv_data_78 : _GEN_5722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5724 = 8'h4f == _match_key_qbytes_5_T ? phv_data_79 : _GEN_5723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5725 = 8'h50 == _match_key_qbytes_5_T ? phv_data_80 : _GEN_5724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5726 = 8'h51 == _match_key_qbytes_5_T ? phv_data_81 : _GEN_5725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5727 = 8'h52 == _match_key_qbytes_5_T ? phv_data_82 : _GEN_5726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5728 = 8'h53 == _match_key_qbytes_5_T ? phv_data_83 : _GEN_5727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5729 = 8'h54 == _match_key_qbytes_5_T ? phv_data_84 : _GEN_5728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5730 = 8'h55 == _match_key_qbytes_5_T ? phv_data_85 : _GEN_5729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5731 = 8'h56 == _match_key_qbytes_5_T ? phv_data_86 : _GEN_5730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5732 = 8'h57 == _match_key_qbytes_5_T ? phv_data_87 : _GEN_5731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5733 = 8'h58 == _match_key_qbytes_5_T ? phv_data_88 : _GEN_5732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5734 = 8'h59 == _match_key_qbytes_5_T ? phv_data_89 : _GEN_5733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5735 = 8'h5a == _match_key_qbytes_5_T ? phv_data_90 : _GEN_5734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5736 = 8'h5b == _match_key_qbytes_5_T ? phv_data_91 : _GEN_5735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5737 = 8'h5c == _match_key_qbytes_5_T ? phv_data_92 : _GEN_5736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5738 = 8'h5d == _match_key_qbytes_5_T ? phv_data_93 : _GEN_5737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5739 = 8'h5e == _match_key_qbytes_5_T ? phv_data_94 : _GEN_5738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5740 = 8'h5f == _match_key_qbytes_5_T ? phv_data_95 : _GEN_5739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5741 = 8'h60 == _match_key_qbytes_5_T ? phv_data_96 : _GEN_5740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5742 = 8'h61 == _match_key_qbytes_5_T ? phv_data_97 : _GEN_5741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5743 = 8'h62 == _match_key_qbytes_5_T ? phv_data_98 : _GEN_5742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5744 = 8'h63 == _match_key_qbytes_5_T ? phv_data_99 : _GEN_5743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5745 = 8'h64 == _match_key_qbytes_5_T ? phv_data_100 : _GEN_5744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5746 = 8'h65 == _match_key_qbytes_5_T ? phv_data_101 : _GEN_5745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5747 = 8'h66 == _match_key_qbytes_5_T ? phv_data_102 : _GEN_5746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5748 = 8'h67 == _match_key_qbytes_5_T ? phv_data_103 : _GEN_5747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5749 = 8'h68 == _match_key_qbytes_5_T ? phv_data_104 : _GEN_5748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5750 = 8'h69 == _match_key_qbytes_5_T ? phv_data_105 : _GEN_5749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5751 = 8'h6a == _match_key_qbytes_5_T ? phv_data_106 : _GEN_5750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5752 = 8'h6b == _match_key_qbytes_5_T ? phv_data_107 : _GEN_5751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5753 = 8'h6c == _match_key_qbytes_5_T ? phv_data_108 : _GEN_5752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5754 = 8'h6d == _match_key_qbytes_5_T ? phv_data_109 : _GEN_5753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5755 = 8'h6e == _match_key_qbytes_5_T ? phv_data_110 : _GEN_5754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5756 = 8'h6f == _match_key_qbytes_5_T ? phv_data_111 : _GEN_5755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5757 = 8'h70 == _match_key_qbytes_5_T ? phv_data_112 : _GEN_5756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5758 = 8'h71 == _match_key_qbytes_5_T ? phv_data_113 : _GEN_5757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5759 = 8'h72 == _match_key_qbytes_5_T ? phv_data_114 : _GEN_5758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5760 = 8'h73 == _match_key_qbytes_5_T ? phv_data_115 : _GEN_5759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5761 = 8'h74 == _match_key_qbytes_5_T ? phv_data_116 : _GEN_5760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5762 = 8'h75 == _match_key_qbytes_5_T ? phv_data_117 : _GEN_5761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5763 = 8'h76 == _match_key_qbytes_5_T ? phv_data_118 : _GEN_5762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5764 = 8'h77 == _match_key_qbytes_5_T ? phv_data_119 : _GEN_5763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5765 = 8'h78 == _match_key_qbytes_5_T ? phv_data_120 : _GEN_5764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5766 = 8'h79 == _match_key_qbytes_5_T ? phv_data_121 : _GEN_5765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5767 = 8'h7a == _match_key_qbytes_5_T ? phv_data_122 : _GEN_5766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5768 = 8'h7b == _match_key_qbytes_5_T ? phv_data_123 : _GEN_5767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5769 = 8'h7c == _match_key_qbytes_5_T ? phv_data_124 : _GEN_5768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5770 = 8'h7d == _match_key_qbytes_5_T ? phv_data_125 : _GEN_5769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5771 = 8'h7e == _match_key_qbytes_5_T ? phv_data_126 : _GEN_5770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5772 = 8'h7f == _match_key_qbytes_5_T ? phv_data_127 : _GEN_5771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5773 = 8'h80 == _match_key_qbytes_5_T ? phv_data_128 : _GEN_5772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5774 = 8'h81 == _match_key_qbytes_5_T ? phv_data_129 : _GEN_5773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5775 = 8'h82 == _match_key_qbytes_5_T ? phv_data_130 : _GEN_5774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5776 = 8'h83 == _match_key_qbytes_5_T ? phv_data_131 : _GEN_5775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5777 = 8'h84 == _match_key_qbytes_5_T ? phv_data_132 : _GEN_5776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5778 = 8'h85 == _match_key_qbytes_5_T ? phv_data_133 : _GEN_5777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5779 = 8'h86 == _match_key_qbytes_5_T ? phv_data_134 : _GEN_5778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5780 = 8'h87 == _match_key_qbytes_5_T ? phv_data_135 : _GEN_5779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5781 = 8'h88 == _match_key_qbytes_5_T ? phv_data_136 : _GEN_5780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5782 = 8'h89 == _match_key_qbytes_5_T ? phv_data_137 : _GEN_5781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5783 = 8'h8a == _match_key_qbytes_5_T ? phv_data_138 : _GEN_5782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5784 = 8'h8b == _match_key_qbytes_5_T ? phv_data_139 : _GEN_5783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5785 = 8'h8c == _match_key_qbytes_5_T ? phv_data_140 : _GEN_5784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5786 = 8'h8d == _match_key_qbytes_5_T ? phv_data_141 : _GEN_5785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5787 = 8'h8e == _match_key_qbytes_5_T ? phv_data_142 : _GEN_5786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5788 = 8'h8f == _match_key_qbytes_5_T ? phv_data_143 : _GEN_5787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5789 = 8'h90 == _match_key_qbytes_5_T ? phv_data_144 : _GEN_5788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5790 = 8'h91 == _match_key_qbytes_5_T ? phv_data_145 : _GEN_5789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5791 = 8'h92 == _match_key_qbytes_5_T ? phv_data_146 : _GEN_5790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5792 = 8'h93 == _match_key_qbytes_5_T ? phv_data_147 : _GEN_5791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5793 = 8'h94 == _match_key_qbytes_5_T ? phv_data_148 : _GEN_5792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5794 = 8'h95 == _match_key_qbytes_5_T ? phv_data_149 : _GEN_5793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5795 = 8'h96 == _match_key_qbytes_5_T ? phv_data_150 : _GEN_5794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5796 = 8'h97 == _match_key_qbytes_5_T ? phv_data_151 : _GEN_5795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5797 = 8'h98 == _match_key_qbytes_5_T ? phv_data_152 : _GEN_5796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5798 = 8'h99 == _match_key_qbytes_5_T ? phv_data_153 : _GEN_5797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5799 = 8'h9a == _match_key_qbytes_5_T ? phv_data_154 : _GEN_5798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5800 = 8'h9b == _match_key_qbytes_5_T ? phv_data_155 : _GEN_5799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5801 = 8'h9c == _match_key_qbytes_5_T ? phv_data_156 : _GEN_5800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5802 = 8'h9d == _match_key_qbytes_5_T ? phv_data_157 : _GEN_5801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5803 = 8'h9e == _match_key_qbytes_5_T ? phv_data_158 : _GEN_5802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5804 = 8'h9f == _match_key_qbytes_5_T ? phv_data_159 : _GEN_5803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5805 = 8'ha0 == _match_key_qbytes_5_T ? phv_data_160 : _GEN_5804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5806 = 8'ha1 == _match_key_qbytes_5_T ? phv_data_161 : _GEN_5805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5807 = 8'ha2 == _match_key_qbytes_5_T ? phv_data_162 : _GEN_5806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5808 = 8'ha3 == _match_key_qbytes_5_T ? phv_data_163 : _GEN_5807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5809 = 8'ha4 == _match_key_qbytes_5_T ? phv_data_164 : _GEN_5808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5810 = 8'ha5 == _match_key_qbytes_5_T ? phv_data_165 : _GEN_5809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5811 = 8'ha6 == _match_key_qbytes_5_T ? phv_data_166 : _GEN_5810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5812 = 8'ha7 == _match_key_qbytes_5_T ? phv_data_167 : _GEN_5811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5813 = 8'ha8 == _match_key_qbytes_5_T ? phv_data_168 : _GEN_5812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5814 = 8'ha9 == _match_key_qbytes_5_T ? phv_data_169 : _GEN_5813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5815 = 8'haa == _match_key_qbytes_5_T ? phv_data_170 : _GEN_5814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5816 = 8'hab == _match_key_qbytes_5_T ? phv_data_171 : _GEN_5815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5817 = 8'hac == _match_key_qbytes_5_T ? phv_data_172 : _GEN_5816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5818 = 8'had == _match_key_qbytes_5_T ? phv_data_173 : _GEN_5817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5819 = 8'hae == _match_key_qbytes_5_T ? phv_data_174 : _GEN_5818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5820 = 8'haf == _match_key_qbytes_5_T ? phv_data_175 : _GEN_5819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5821 = 8'hb0 == _match_key_qbytes_5_T ? phv_data_176 : _GEN_5820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5822 = 8'hb1 == _match_key_qbytes_5_T ? phv_data_177 : _GEN_5821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5823 = 8'hb2 == _match_key_qbytes_5_T ? phv_data_178 : _GEN_5822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5824 = 8'hb3 == _match_key_qbytes_5_T ? phv_data_179 : _GEN_5823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5825 = 8'hb4 == _match_key_qbytes_5_T ? phv_data_180 : _GEN_5824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5826 = 8'hb5 == _match_key_qbytes_5_T ? phv_data_181 : _GEN_5825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5827 = 8'hb6 == _match_key_qbytes_5_T ? phv_data_182 : _GEN_5826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5828 = 8'hb7 == _match_key_qbytes_5_T ? phv_data_183 : _GEN_5827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5829 = 8'hb8 == _match_key_qbytes_5_T ? phv_data_184 : _GEN_5828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5830 = 8'hb9 == _match_key_qbytes_5_T ? phv_data_185 : _GEN_5829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5831 = 8'hba == _match_key_qbytes_5_T ? phv_data_186 : _GEN_5830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5832 = 8'hbb == _match_key_qbytes_5_T ? phv_data_187 : _GEN_5831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5833 = 8'hbc == _match_key_qbytes_5_T ? phv_data_188 : _GEN_5832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5834 = 8'hbd == _match_key_qbytes_5_T ? phv_data_189 : _GEN_5833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5835 = 8'hbe == _match_key_qbytes_5_T ? phv_data_190 : _GEN_5834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5836 = 8'hbf == _match_key_qbytes_5_T ? phv_data_191 : _GEN_5835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5837 = 8'hc0 == _match_key_qbytes_5_T ? phv_data_192 : _GEN_5836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5838 = 8'hc1 == _match_key_qbytes_5_T ? phv_data_193 : _GEN_5837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5839 = 8'hc2 == _match_key_qbytes_5_T ? phv_data_194 : _GEN_5838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5840 = 8'hc3 == _match_key_qbytes_5_T ? phv_data_195 : _GEN_5839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5841 = 8'hc4 == _match_key_qbytes_5_T ? phv_data_196 : _GEN_5840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5842 = 8'hc5 == _match_key_qbytes_5_T ? phv_data_197 : _GEN_5841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5843 = 8'hc6 == _match_key_qbytes_5_T ? phv_data_198 : _GEN_5842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5844 = 8'hc7 == _match_key_qbytes_5_T ? phv_data_199 : _GEN_5843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5845 = 8'hc8 == _match_key_qbytes_5_T ? phv_data_200 : _GEN_5844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5846 = 8'hc9 == _match_key_qbytes_5_T ? phv_data_201 : _GEN_5845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5847 = 8'hca == _match_key_qbytes_5_T ? phv_data_202 : _GEN_5846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5848 = 8'hcb == _match_key_qbytes_5_T ? phv_data_203 : _GEN_5847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5849 = 8'hcc == _match_key_qbytes_5_T ? phv_data_204 : _GEN_5848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5850 = 8'hcd == _match_key_qbytes_5_T ? phv_data_205 : _GEN_5849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5851 = 8'hce == _match_key_qbytes_5_T ? phv_data_206 : _GEN_5850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5852 = 8'hcf == _match_key_qbytes_5_T ? phv_data_207 : _GEN_5851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5853 = 8'hd0 == _match_key_qbytes_5_T ? phv_data_208 : _GEN_5852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5854 = 8'hd1 == _match_key_qbytes_5_T ? phv_data_209 : _GEN_5853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5855 = 8'hd2 == _match_key_qbytes_5_T ? phv_data_210 : _GEN_5854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5856 = 8'hd3 == _match_key_qbytes_5_T ? phv_data_211 : _GEN_5855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5857 = 8'hd4 == _match_key_qbytes_5_T ? phv_data_212 : _GEN_5856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5858 = 8'hd5 == _match_key_qbytes_5_T ? phv_data_213 : _GEN_5857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5859 = 8'hd6 == _match_key_qbytes_5_T ? phv_data_214 : _GEN_5858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5860 = 8'hd7 == _match_key_qbytes_5_T ? phv_data_215 : _GEN_5859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5861 = 8'hd8 == _match_key_qbytes_5_T ? phv_data_216 : _GEN_5860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5862 = 8'hd9 == _match_key_qbytes_5_T ? phv_data_217 : _GEN_5861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5863 = 8'hda == _match_key_qbytes_5_T ? phv_data_218 : _GEN_5862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5864 = 8'hdb == _match_key_qbytes_5_T ? phv_data_219 : _GEN_5863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5865 = 8'hdc == _match_key_qbytes_5_T ? phv_data_220 : _GEN_5864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5866 = 8'hdd == _match_key_qbytes_5_T ? phv_data_221 : _GEN_5865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5867 = 8'hde == _match_key_qbytes_5_T ? phv_data_222 : _GEN_5866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5868 = 8'hdf == _match_key_qbytes_5_T ? phv_data_223 : _GEN_5867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5869 = 8'he0 == _match_key_qbytes_5_T ? phv_data_224 : _GEN_5868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5870 = 8'he1 == _match_key_qbytes_5_T ? phv_data_225 : _GEN_5869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5871 = 8'he2 == _match_key_qbytes_5_T ? phv_data_226 : _GEN_5870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5872 = 8'he3 == _match_key_qbytes_5_T ? phv_data_227 : _GEN_5871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5873 = 8'he4 == _match_key_qbytes_5_T ? phv_data_228 : _GEN_5872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5874 = 8'he5 == _match_key_qbytes_5_T ? phv_data_229 : _GEN_5873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5875 = 8'he6 == _match_key_qbytes_5_T ? phv_data_230 : _GEN_5874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5876 = 8'he7 == _match_key_qbytes_5_T ? phv_data_231 : _GEN_5875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5877 = 8'he8 == _match_key_qbytes_5_T ? phv_data_232 : _GEN_5876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5878 = 8'he9 == _match_key_qbytes_5_T ? phv_data_233 : _GEN_5877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5879 = 8'hea == _match_key_qbytes_5_T ? phv_data_234 : _GEN_5878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5880 = 8'heb == _match_key_qbytes_5_T ? phv_data_235 : _GEN_5879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5881 = 8'hec == _match_key_qbytes_5_T ? phv_data_236 : _GEN_5880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5882 = 8'hed == _match_key_qbytes_5_T ? phv_data_237 : _GEN_5881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5883 = 8'hee == _match_key_qbytes_5_T ? phv_data_238 : _GEN_5882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5884 = 8'hef == _match_key_qbytes_5_T ? phv_data_239 : _GEN_5883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5885 = 8'hf0 == _match_key_qbytes_5_T ? phv_data_240 : _GEN_5884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5886 = 8'hf1 == _match_key_qbytes_5_T ? phv_data_241 : _GEN_5885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5887 = 8'hf2 == _match_key_qbytes_5_T ? phv_data_242 : _GEN_5886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5888 = 8'hf3 == _match_key_qbytes_5_T ? phv_data_243 : _GEN_5887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5889 = 8'hf4 == _match_key_qbytes_5_T ? phv_data_244 : _GEN_5888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5890 = 8'hf5 == _match_key_qbytes_5_T ? phv_data_245 : _GEN_5889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5891 = 8'hf6 == _match_key_qbytes_5_T ? phv_data_246 : _GEN_5890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5892 = 8'hf7 == _match_key_qbytes_5_T ? phv_data_247 : _GEN_5891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5893 = 8'hf8 == _match_key_qbytes_5_T ? phv_data_248 : _GEN_5892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5894 = 8'hf9 == _match_key_qbytes_5_T ? phv_data_249 : _GEN_5893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5895 = 8'hfa == _match_key_qbytes_5_T ? phv_data_250 : _GEN_5894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5896 = 8'hfb == _match_key_qbytes_5_T ? phv_data_251 : _GEN_5895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5897 = 8'hfc == _match_key_qbytes_5_T ? phv_data_252 : _GEN_5896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5898 = 8'hfd == _match_key_qbytes_5_T ? phv_data_253 : _GEN_5897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5899 = 8'hfe == _match_key_qbytes_5_T ? phv_data_254 : _GEN_5898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5900 = 8'hff == _match_key_qbytes_5_T ? phv_data_255 : _GEN_5899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5902 = 8'h1 == _match_key_qbytes_5_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5903 = 8'h2 == _match_key_qbytes_5_T_1 ? phv_data_2 : _GEN_5902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5904 = 8'h3 == _match_key_qbytes_5_T_1 ? phv_data_3 : _GEN_5903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5905 = 8'h4 == _match_key_qbytes_5_T_1 ? phv_data_4 : _GEN_5904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5906 = 8'h5 == _match_key_qbytes_5_T_1 ? phv_data_5 : _GEN_5905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5907 = 8'h6 == _match_key_qbytes_5_T_1 ? phv_data_6 : _GEN_5906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5908 = 8'h7 == _match_key_qbytes_5_T_1 ? phv_data_7 : _GEN_5907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5909 = 8'h8 == _match_key_qbytes_5_T_1 ? phv_data_8 : _GEN_5908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5910 = 8'h9 == _match_key_qbytes_5_T_1 ? phv_data_9 : _GEN_5909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5911 = 8'ha == _match_key_qbytes_5_T_1 ? phv_data_10 : _GEN_5910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5912 = 8'hb == _match_key_qbytes_5_T_1 ? phv_data_11 : _GEN_5911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5913 = 8'hc == _match_key_qbytes_5_T_1 ? phv_data_12 : _GEN_5912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5914 = 8'hd == _match_key_qbytes_5_T_1 ? phv_data_13 : _GEN_5913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5915 = 8'he == _match_key_qbytes_5_T_1 ? phv_data_14 : _GEN_5914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5916 = 8'hf == _match_key_qbytes_5_T_1 ? phv_data_15 : _GEN_5915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5917 = 8'h10 == _match_key_qbytes_5_T_1 ? phv_data_16 : _GEN_5916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5918 = 8'h11 == _match_key_qbytes_5_T_1 ? phv_data_17 : _GEN_5917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5919 = 8'h12 == _match_key_qbytes_5_T_1 ? phv_data_18 : _GEN_5918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5920 = 8'h13 == _match_key_qbytes_5_T_1 ? phv_data_19 : _GEN_5919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5921 = 8'h14 == _match_key_qbytes_5_T_1 ? phv_data_20 : _GEN_5920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5922 = 8'h15 == _match_key_qbytes_5_T_1 ? phv_data_21 : _GEN_5921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5923 = 8'h16 == _match_key_qbytes_5_T_1 ? phv_data_22 : _GEN_5922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5924 = 8'h17 == _match_key_qbytes_5_T_1 ? phv_data_23 : _GEN_5923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5925 = 8'h18 == _match_key_qbytes_5_T_1 ? phv_data_24 : _GEN_5924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5926 = 8'h19 == _match_key_qbytes_5_T_1 ? phv_data_25 : _GEN_5925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5927 = 8'h1a == _match_key_qbytes_5_T_1 ? phv_data_26 : _GEN_5926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5928 = 8'h1b == _match_key_qbytes_5_T_1 ? phv_data_27 : _GEN_5927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5929 = 8'h1c == _match_key_qbytes_5_T_1 ? phv_data_28 : _GEN_5928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5930 = 8'h1d == _match_key_qbytes_5_T_1 ? phv_data_29 : _GEN_5929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5931 = 8'h1e == _match_key_qbytes_5_T_1 ? phv_data_30 : _GEN_5930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5932 = 8'h1f == _match_key_qbytes_5_T_1 ? phv_data_31 : _GEN_5931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5933 = 8'h20 == _match_key_qbytes_5_T_1 ? phv_data_32 : _GEN_5932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5934 = 8'h21 == _match_key_qbytes_5_T_1 ? phv_data_33 : _GEN_5933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5935 = 8'h22 == _match_key_qbytes_5_T_1 ? phv_data_34 : _GEN_5934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5936 = 8'h23 == _match_key_qbytes_5_T_1 ? phv_data_35 : _GEN_5935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5937 = 8'h24 == _match_key_qbytes_5_T_1 ? phv_data_36 : _GEN_5936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5938 = 8'h25 == _match_key_qbytes_5_T_1 ? phv_data_37 : _GEN_5937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5939 = 8'h26 == _match_key_qbytes_5_T_1 ? phv_data_38 : _GEN_5938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5940 = 8'h27 == _match_key_qbytes_5_T_1 ? phv_data_39 : _GEN_5939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5941 = 8'h28 == _match_key_qbytes_5_T_1 ? phv_data_40 : _GEN_5940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5942 = 8'h29 == _match_key_qbytes_5_T_1 ? phv_data_41 : _GEN_5941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5943 = 8'h2a == _match_key_qbytes_5_T_1 ? phv_data_42 : _GEN_5942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5944 = 8'h2b == _match_key_qbytes_5_T_1 ? phv_data_43 : _GEN_5943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5945 = 8'h2c == _match_key_qbytes_5_T_1 ? phv_data_44 : _GEN_5944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5946 = 8'h2d == _match_key_qbytes_5_T_1 ? phv_data_45 : _GEN_5945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5947 = 8'h2e == _match_key_qbytes_5_T_1 ? phv_data_46 : _GEN_5946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5948 = 8'h2f == _match_key_qbytes_5_T_1 ? phv_data_47 : _GEN_5947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5949 = 8'h30 == _match_key_qbytes_5_T_1 ? phv_data_48 : _GEN_5948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5950 = 8'h31 == _match_key_qbytes_5_T_1 ? phv_data_49 : _GEN_5949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5951 = 8'h32 == _match_key_qbytes_5_T_1 ? phv_data_50 : _GEN_5950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5952 = 8'h33 == _match_key_qbytes_5_T_1 ? phv_data_51 : _GEN_5951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5953 = 8'h34 == _match_key_qbytes_5_T_1 ? phv_data_52 : _GEN_5952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5954 = 8'h35 == _match_key_qbytes_5_T_1 ? phv_data_53 : _GEN_5953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5955 = 8'h36 == _match_key_qbytes_5_T_1 ? phv_data_54 : _GEN_5954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5956 = 8'h37 == _match_key_qbytes_5_T_1 ? phv_data_55 : _GEN_5955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5957 = 8'h38 == _match_key_qbytes_5_T_1 ? phv_data_56 : _GEN_5956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5958 = 8'h39 == _match_key_qbytes_5_T_1 ? phv_data_57 : _GEN_5957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5959 = 8'h3a == _match_key_qbytes_5_T_1 ? phv_data_58 : _GEN_5958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5960 = 8'h3b == _match_key_qbytes_5_T_1 ? phv_data_59 : _GEN_5959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5961 = 8'h3c == _match_key_qbytes_5_T_1 ? phv_data_60 : _GEN_5960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5962 = 8'h3d == _match_key_qbytes_5_T_1 ? phv_data_61 : _GEN_5961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5963 = 8'h3e == _match_key_qbytes_5_T_1 ? phv_data_62 : _GEN_5962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5964 = 8'h3f == _match_key_qbytes_5_T_1 ? phv_data_63 : _GEN_5963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5965 = 8'h40 == _match_key_qbytes_5_T_1 ? phv_data_64 : _GEN_5964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5966 = 8'h41 == _match_key_qbytes_5_T_1 ? phv_data_65 : _GEN_5965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5967 = 8'h42 == _match_key_qbytes_5_T_1 ? phv_data_66 : _GEN_5966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5968 = 8'h43 == _match_key_qbytes_5_T_1 ? phv_data_67 : _GEN_5967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5969 = 8'h44 == _match_key_qbytes_5_T_1 ? phv_data_68 : _GEN_5968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5970 = 8'h45 == _match_key_qbytes_5_T_1 ? phv_data_69 : _GEN_5969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5971 = 8'h46 == _match_key_qbytes_5_T_1 ? phv_data_70 : _GEN_5970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5972 = 8'h47 == _match_key_qbytes_5_T_1 ? phv_data_71 : _GEN_5971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5973 = 8'h48 == _match_key_qbytes_5_T_1 ? phv_data_72 : _GEN_5972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5974 = 8'h49 == _match_key_qbytes_5_T_1 ? phv_data_73 : _GEN_5973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5975 = 8'h4a == _match_key_qbytes_5_T_1 ? phv_data_74 : _GEN_5974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5976 = 8'h4b == _match_key_qbytes_5_T_1 ? phv_data_75 : _GEN_5975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5977 = 8'h4c == _match_key_qbytes_5_T_1 ? phv_data_76 : _GEN_5976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5978 = 8'h4d == _match_key_qbytes_5_T_1 ? phv_data_77 : _GEN_5977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5979 = 8'h4e == _match_key_qbytes_5_T_1 ? phv_data_78 : _GEN_5978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5980 = 8'h4f == _match_key_qbytes_5_T_1 ? phv_data_79 : _GEN_5979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5981 = 8'h50 == _match_key_qbytes_5_T_1 ? phv_data_80 : _GEN_5980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5982 = 8'h51 == _match_key_qbytes_5_T_1 ? phv_data_81 : _GEN_5981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5983 = 8'h52 == _match_key_qbytes_5_T_1 ? phv_data_82 : _GEN_5982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5984 = 8'h53 == _match_key_qbytes_5_T_1 ? phv_data_83 : _GEN_5983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5985 = 8'h54 == _match_key_qbytes_5_T_1 ? phv_data_84 : _GEN_5984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5986 = 8'h55 == _match_key_qbytes_5_T_1 ? phv_data_85 : _GEN_5985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5987 = 8'h56 == _match_key_qbytes_5_T_1 ? phv_data_86 : _GEN_5986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5988 = 8'h57 == _match_key_qbytes_5_T_1 ? phv_data_87 : _GEN_5987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5989 = 8'h58 == _match_key_qbytes_5_T_1 ? phv_data_88 : _GEN_5988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5990 = 8'h59 == _match_key_qbytes_5_T_1 ? phv_data_89 : _GEN_5989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5991 = 8'h5a == _match_key_qbytes_5_T_1 ? phv_data_90 : _GEN_5990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5992 = 8'h5b == _match_key_qbytes_5_T_1 ? phv_data_91 : _GEN_5991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5993 = 8'h5c == _match_key_qbytes_5_T_1 ? phv_data_92 : _GEN_5992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5994 = 8'h5d == _match_key_qbytes_5_T_1 ? phv_data_93 : _GEN_5993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5995 = 8'h5e == _match_key_qbytes_5_T_1 ? phv_data_94 : _GEN_5994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5996 = 8'h5f == _match_key_qbytes_5_T_1 ? phv_data_95 : _GEN_5995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5997 = 8'h60 == _match_key_qbytes_5_T_1 ? phv_data_96 : _GEN_5996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5998 = 8'h61 == _match_key_qbytes_5_T_1 ? phv_data_97 : _GEN_5997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5999 = 8'h62 == _match_key_qbytes_5_T_1 ? phv_data_98 : _GEN_5998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6000 = 8'h63 == _match_key_qbytes_5_T_1 ? phv_data_99 : _GEN_5999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6001 = 8'h64 == _match_key_qbytes_5_T_1 ? phv_data_100 : _GEN_6000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6002 = 8'h65 == _match_key_qbytes_5_T_1 ? phv_data_101 : _GEN_6001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6003 = 8'h66 == _match_key_qbytes_5_T_1 ? phv_data_102 : _GEN_6002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6004 = 8'h67 == _match_key_qbytes_5_T_1 ? phv_data_103 : _GEN_6003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6005 = 8'h68 == _match_key_qbytes_5_T_1 ? phv_data_104 : _GEN_6004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6006 = 8'h69 == _match_key_qbytes_5_T_1 ? phv_data_105 : _GEN_6005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6007 = 8'h6a == _match_key_qbytes_5_T_1 ? phv_data_106 : _GEN_6006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6008 = 8'h6b == _match_key_qbytes_5_T_1 ? phv_data_107 : _GEN_6007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6009 = 8'h6c == _match_key_qbytes_5_T_1 ? phv_data_108 : _GEN_6008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6010 = 8'h6d == _match_key_qbytes_5_T_1 ? phv_data_109 : _GEN_6009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6011 = 8'h6e == _match_key_qbytes_5_T_1 ? phv_data_110 : _GEN_6010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6012 = 8'h6f == _match_key_qbytes_5_T_1 ? phv_data_111 : _GEN_6011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6013 = 8'h70 == _match_key_qbytes_5_T_1 ? phv_data_112 : _GEN_6012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6014 = 8'h71 == _match_key_qbytes_5_T_1 ? phv_data_113 : _GEN_6013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6015 = 8'h72 == _match_key_qbytes_5_T_1 ? phv_data_114 : _GEN_6014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6016 = 8'h73 == _match_key_qbytes_5_T_1 ? phv_data_115 : _GEN_6015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6017 = 8'h74 == _match_key_qbytes_5_T_1 ? phv_data_116 : _GEN_6016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6018 = 8'h75 == _match_key_qbytes_5_T_1 ? phv_data_117 : _GEN_6017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6019 = 8'h76 == _match_key_qbytes_5_T_1 ? phv_data_118 : _GEN_6018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6020 = 8'h77 == _match_key_qbytes_5_T_1 ? phv_data_119 : _GEN_6019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6021 = 8'h78 == _match_key_qbytes_5_T_1 ? phv_data_120 : _GEN_6020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6022 = 8'h79 == _match_key_qbytes_5_T_1 ? phv_data_121 : _GEN_6021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6023 = 8'h7a == _match_key_qbytes_5_T_1 ? phv_data_122 : _GEN_6022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6024 = 8'h7b == _match_key_qbytes_5_T_1 ? phv_data_123 : _GEN_6023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6025 = 8'h7c == _match_key_qbytes_5_T_1 ? phv_data_124 : _GEN_6024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6026 = 8'h7d == _match_key_qbytes_5_T_1 ? phv_data_125 : _GEN_6025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6027 = 8'h7e == _match_key_qbytes_5_T_1 ? phv_data_126 : _GEN_6026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6028 = 8'h7f == _match_key_qbytes_5_T_1 ? phv_data_127 : _GEN_6027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6029 = 8'h80 == _match_key_qbytes_5_T_1 ? phv_data_128 : _GEN_6028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6030 = 8'h81 == _match_key_qbytes_5_T_1 ? phv_data_129 : _GEN_6029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6031 = 8'h82 == _match_key_qbytes_5_T_1 ? phv_data_130 : _GEN_6030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6032 = 8'h83 == _match_key_qbytes_5_T_1 ? phv_data_131 : _GEN_6031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6033 = 8'h84 == _match_key_qbytes_5_T_1 ? phv_data_132 : _GEN_6032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6034 = 8'h85 == _match_key_qbytes_5_T_1 ? phv_data_133 : _GEN_6033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6035 = 8'h86 == _match_key_qbytes_5_T_1 ? phv_data_134 : _GEN_6034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6036 = 8'h87 == _match_key_qbytes_5_T_1 ? phv_data_135 : _GEN_6035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6037 = 8'h88 == _match_key_qbytes_5_T_1 ? phv_data_136 : _GEN_6036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6038 = 8'h89 == _match_key_qbytes_5_T_1 ? phv_data_137 : _GEN_6037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6039 = 8'h8a == _match_key_qbytes_5_T_1 ? phv_data_138 : _GEN_6038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6040 = 8'h8b == _match_key_qbytes_5_T_1 ? phv_data_139 : _GEN_6039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6041 = 8'h8c == _match_key_qbytes_5_T_1 ? phv_data_140 : _GEN_6040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6042 = 8'h8d == _match_key_qbytes_5_T_1 ? phv_data_141 : _GEN_6041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6043 = 8'h8e == _match_key_qbytes_5_T_1 ? phv_data_142 : _GEN_6042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6044 = 8'h8f == _match_key_qbytes_5_T_1 ? phv_data_143 : _GEN_6043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6045 = 8'h90 == _match_key_qbytes_5_T_1 ? phv_data_144 : _GEN_6044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6046 = 8'h91 == _match_key_qbytes_5_T_1 ? phv_data_145 : _GEN_6045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6047 = 8'h92 == _match_key_qbytes_5_T_1 ? phv_data_146 : _GEN_6046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6048 = 8'h93 == _match_key_qbytes_5_T_1 ? phv_data_147 : _GEN_6047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6049 = 8'h94 == _match_key_qbytes_5_T_1 ? phv_data_148 : _GEN_6048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6050 = 8'h95 == _match_key_qbytes_5_T_1 ? phv_data_149 : _GEN_6049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6051 = 8'h96 == _match_key_qbytes_5_T_1 ? phv_data_150 : _GEN_6050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6052 = 8'h97 == _match_key_qbytes_5_T_1 ? phv_data_151 : _GEN_6051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6053 = 8'h98 == _match_key_qbytes_5_T_1 ? phv_data_152 : _GEN_6052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6054 = 8'h99 == _match_key_qbytes_5_T_1 ? phv_data_153 : _GEN_6053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6055 = 8'h9a == _match_key_qbytes_5_T_1 ? phv_data_154 : _GEN_6054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6056 = 8'h9b == _match_key_qbytes_5_T_1 ? phv_data_155 : _GEN_6055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6057 = 8'h9c == _match_key_qbytes_5_T_1 ? phv_data_156 : _GEN_6056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6058 = 8'h9d == _match_key_qbytes_5_T_1 ? phv_data_157 : _GEN_6057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6059 = 8'h9e == _match_key_qbytes_5_T_1 ? phv_data_158 : _GEN_6058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6060 = 8'h9f == _match_key_qbytes_5_T_1 ? phv_data_159 : _GEN_6059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6061 = 8'ha0 == _match_key_qbytes_5_T_1 ? phv_data_160 : _GEN_6060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6062 = 8'ha1 == _match_key_qbytes_5_T_1 ? phv_data_161 : _GEN_6061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6063 = 8'ha2 == _match_key_qbytes_5_T_1 ? phv_data_162 : _GEN_6062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6064 = 8'ha3 == _match_key_qbytes_5_T_1 ? phv_data_163 : _GEN_6063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6065 = 8'ha4 == _match_key_qbytes_5_T_1 ? phv_data_164 : _GEN_6064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6066 = 8'ha5 == _match_key_qbytes_5_T_1 ? phv_data_165 : _GEN_6065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6067 = 8'ha6 == _match_key_qbytes_5_T_1 ? phv_data_166 : _GEN_6066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6068 = 8'ha7 == _match_key_qbytes_5_T_1 ? phv_data_167 : _GEN_6067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6069 = 8'ha8 == _match_key_qbytes_5_T_1 ? phv_data_168 : _GEN_6068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6070 = 8'ha9 == _match_key_qbytes_5_T_1 ? phv_data_169 : _GEN_6069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6071 = 8'haa == _match_key_qbytes_5_T_1 ? phv_data_170 : _GEN_6070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6072 = 8'hab == _match_key_qbytes_5_T_1 ? phv_data_171 : _GEN_6071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6073 = 8'hac == _match_key_qbytes_5_T_1 ? phv_data_172 : _GEN_6072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6074 = 8'had == _match_key_qbytes_5_T_1 ? phv_data_173 : _GEN_6073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6075 = 8'hae == _match_key_qbytes_5_T_1 ? phv_data_174 : _GEN_6074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6076 = 8'haf == _match_key_qbytes_5_T_1 ? phv_data_175 : _GEN_6075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6077 = 8'hb0 == _match_key_qbytes_5_T_1 ? phv_data_176 : _GEN_6076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6078 = 8'hb1 == _match_key_qbytes_5_T_1 ? phv_data_177 : _GEN_6077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6079 = 8'hb2 == _match_key_qbytes_5_T_1 ? phv_data_178 : _GEN_6078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6080 = 8'hb3 == _match_key_qbytes_5_T_1 ? phv_data_179 : _GEN_6079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6081 = 8'hb4 == _match_key_qbytes_5_T_1 ? phv_data_180 : _GEN_6080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6082 = 8'hb5 == _match_key_qbytes_5_T_1 ? phv_data_181 : _GEN_6081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6083 = 8'hb6 == _match_key_qbytes_5_T_1 ? phv_data_182 : _GEN_6082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6084 = 8'hb7 == _match_key_qbytes_5_T_1 ? phv_data_183 : _GEN_6083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6085 = 8'hb8 == _match_key_qbytes_5_T_1 ? phv_data_184 : _GEN_6084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6086 = 8'hb9 == _match_key_qbytes_5_T_1 ? phv_data_185 : _GEN_6085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6087 = 8'hba == _match_key_qbytes_5_T_1 ? phv_data_186 : _GEN_6086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6088 = 8'hbb == _match_key_qbytes_5_T_1 ? phv_data_187 : _GEN_6087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6089 = 8'hbc == _match_key_qbytes_5_T_1 ? phv_data_188 : _GEN_6088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6090 = 8'hbd == _match_key_qbytes_5_T_1 ? phv_data_189 : _GEN_6089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6091 = 8'hbe == _match_key_qbytes_5_T_1 ? phv_data_190 : _GEN_6090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6092 = 8'hbf == _match_key_qbytes_5_T_1 ? phv_data_191 : _GEN_6091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6093 = 8'hc0 == _match_key_qbytes_5_T_1 ? phv_data_192 : _GEN_6092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6094 = 8'hc1 == _match_key_qbytes_5_T_1 ? phv_data_193 : _GEN_6093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6095 = 8'hc2 == _match_key_qbytes_5_T_1 ? phv_data_194 : _GEN_6094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6096 = 8'hc3 == _match_key_qbytes_5_T_1 ? phv_data_195 : _GEN_6095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6097 = 8'hc4 == _match_key_qbytes_5_T_1 ? phv_data_196 : _GEN_6096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6098 = 8'hc5 == _match_key_qbytes_5_T_1 ? phv_data_197 : _GEN_6097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6099 = 8'hc6 == _match_key_qbytes_5_T_1 ? phv_data_198 : _GEN_6098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6100 = 8'hc7 == _match_key_qbytes_5_T_1 ? phv_data_199 : _GEN_6099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6101 = 8'hc8 == _match_key_qbytes_5_T_1 ? phv_data_200 : _GEN_6100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6102 = 8'hc9 == _match_key_qbytes_5_T_1 ? phv_data_201 : _GEN_6101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6103 = 8'hca == _match_key_qbytes_5_T_1 ? phv_data_202 : _GEN_6102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6104 = 8'hcb == _match_key_qbytes_5_T_1 ? phv_data_203 : _GEN_6103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6105 = 8'hcc == _match_key_qbytes_5_T_1 ? phv_data_204 : _GEN_6104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6106 = 8'hcd == _match_key_qbytes_5_T_1 ? phv_data_205 : _GEN_6105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6107 = 8'hce == _match_key_qbytes_5_T_1 ? phv_data_206 : _GEN_6106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6108 = 8'hcf == _match_key_qbytes_5_T_1 ? phv_data_207 : _GEN_6107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6109 = 8'hd0 == _match_key_qbytes_5_T_1 ? phv_data_208 : _GEN_6108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6110 = 8'hd1 == _match_key_qbytes_5_T_1 ? phv_data_209 : _GEN_6109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6111 = 8'hd2 == _match_key_qbytes_5_T_1 ? phv_data_210 : _GEN_6110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6112 = 8'hd3 == _match_key_qbytes_5_T_1 ? phv_data_211 : _GEN_6111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6113 = 8'hd4 == _match_key_qbytes_5_T_1 ? phv_data_212 : _GEN_6112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6114 = 8'hd5 == _match_key_qbytes_5_T_1 ? phv_data_213 : _GEN_6113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6115 = 8'hd6 == _match_key_qbytes_5_T_1 ? phv_data_214 : _GEN_6114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6116 = 8'hd7 == _match_key_qbytes_5_T_1 ? phv_data_215 : _GEN_6115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6117 = 8'hd8 == _match_key_qbytes_5_T_1 ? phv_data_216 : _GEN_6116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6118 = 8'hd9 == _match_key_qbytes_5_T_1 ? phv_data_217 : _GEN_6117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6119 = 8'hda == _match_key_qbytes_5_T_1 ? phv_data_218 : _GEN_6118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6120 = 8'hdb == _match_key_qbytes_5_T_1 ? phv_data_219 : _GEN_6119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6121 = 8'hdc == _match_key_qbytes_5_T_1 ? phv_data_220 : _GEN_6120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6122 = 8'hdd == _match_key_qbytes_5_T_1 ? phv_data_221 : _GEN_6121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6123 = 8'hde == _match_key_qbytes_5_T_1 ? phv_data_222 : _GEN_6122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6124 = 8'hdf == _match_key_qbytes_5_T_1 ? phv_data_223 : _GEN_6123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6125 = 8'he0 == _match_key_qbytes_5_T_1 ? phv_data_224 : _GEN_6124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6126 = 8'he1 == _match_key_qbytes_5_T_1 ? phv_data_225 : _GEN_6125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6127 = 8'he2 == _match_key_qbytes_5_T_1 ? phv_data_226 : _GEN_6126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6128 = 8'he3 == _match_key_qbytes_5_T_1 ? phv_data_227 : _GEN_6127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6129 = 8'he4 == _match_key_qbytes_5_T_1 ? phv_data_228 : _GEN_6128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6130 = 8'he5 == _match_key_qbytes_5_T_1 ? phv_data_229 : _GEN_6129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6131 = 8'he6 == _match_key_qbytes_5_T_1 ? phv_data_230 : _GEN_6130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6132 = 8'he7 == _match_key_qbytes_5_T_1 ? phv_data_231 : _GEN_6131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6133 = 8'he8 == _match_key_qbytes_5_T_1 ? phv_data_232 : _GEN_6132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6134 = 8'he9 == _match_key_qbytes_5_T_1 ? phv_data_233 : _GEN_6133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6135 = 8'hea == _match_key_qbytes_5_T_1 ? phv_data_234 : _GEN_6134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6136 = 8'heb == _match_key_qbytes_5_T_1 ? phv_data_235 : _GEN_6135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6137 = 8'hec == _match_key_qbytes_5_T_1 ? phv_data_236 : _GEN_6136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6138 = 8'hed == _match_key_qbytes_5_T_1 ? phv_data_237 : _GEN_6137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6139 = 8'hee == _match_key_qbytes_5_T_1 ? phv_data_238 : _GEN_6138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6140 = 8'hef == _match_key_qbytes_5_T_1 ? phv_data_239 : _GEN_6139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6141 = 8'hf0 == _match_key_qbytes_5_T_1 ? phv_data_240 : _GEN_6140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6142 = 8'hf1 == _match_key_qbytes_5_T_1 ? phv_data_241 : _GEN_6141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6143 = 8'hf2 == _match_key_qbytes_5_T_1 ? phv_data_242 : _GEN_6142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6144 = 8'hf3 == _match_key_qbytes_5_T_1 ? phv_data_243 : _GEN_6143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6145 = 8'hf4 == _match_key_qbytes_5_T_1 ? phv_data_244 : _GEN_6144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6146 = 8'hf5 == _match_key_qbytes_5_T_1 ? phv_data_245 : _GEN_6145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6147 = 8'hf6 == _match_key_qbytes_5_T_1 ? phv_data_246 : _GEN_6146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6148 = 8'hf7 == _match_key_qbytes_5_T_1 ? phv_data_247 : _GEN_6147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6149 = 8'hf8 == _match_key_qbytes_5_T_1 ? phv_data_248 : _GEN_6148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6150 = 8'hf9 == _match_key_qbytes_5_T_1 ? phv_data_249 : _GEN_6149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6151 = 8'hfa == _match_key_qbytes_5_T_1 ? phv_data_250 : _GEN_6150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6152 = 8'hfb == _match_key_qbytes_5_T_1 ? phv_data_251 : _GEN_6151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6153 = 8'hfc == _match_key_qbytes_5_T_1 ? phv_data_252 : _GEN_6152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6154 = 8'hfd == _match_key_qbytes_5_T_1 ? phv_data_253 : _GEN_6153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6155 = 8'hfe == _match_key_qbytes_5_T_1 ? phv_data_254 : _GEN_6154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6156 = 8'hff == _match_key_qbytes_5_T_1 ? phv_data_255 : _GEN_6155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_5_T_3 = {_GEN_5900,_GEN_6156,_GEN_5388,_GEN_5644}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_5 = local_offset_5 < end_offset ? _match_key_qbytes_5_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 69:29]
  assign io_bias_out = key_offset[1:0]; // @[matcher.scala 79:38]
  assign io_match_key_bytes_0 = phv_is_valid_processor ? match_key_qbytes_0[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_1 = phv_is_valid_processor ? match_key_qbytes_0[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_2 = phv_is_valid_processor ? match_key_qbytes_0[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_3 = phv_is_valid_processor ? match_key_qbytes_0[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_4 = phv_is_valid_processor ? match_key_qbytes_1[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_5 = phv_is_valid_processor ? match_key_qbytes_1[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_6 = phv_is_valid_processor ? match_key_qbytes_1[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_7 = phv_is_valid_processor ? match_key_qbytes_1[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_8 = phv_is_valid_processor ? match_key_qbytes_2[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_9 = phv_is_valid_processor ? match_key_qbytes_2[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_10 = phv_is_valid_processor ? match_key_qbytes_2[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_11 = phv_is_valid_processor ? match_key_qbytes_2[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_12 = phv_is_valid_processor ? match_key_qbytes_3[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_13 = phv_is_valid_processor ? match_key_qbytes_3[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_14 = phv_is_valid_processor ? match_key_qbytes_3[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_15 = phv_is_valid_processor ? match_key_qbytes_3[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_16 = phv_is_valid_processor ? match_key_qbytes_4[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_17 = phv_is_valid_processor ? match_key_qbytes_4[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_18 = phv_is_valid_processor ? match_key_qbytes_4[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_19 = phv_is_valid_processor ? match_key_qbytes_4[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_20 = phv_is_valid_processor ? match_key_qbytes_5[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_21 = phv_is_valid_processor ? match_key_qbytes_5[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_22 = phv_is_valid_processor ? match_key_qbytes_5[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_23 = phv_is_valid_processor ? match_key_qbytes_5[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 68:17]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 68:17]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 68:17]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 68:17]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 68:17]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 68:17]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 68:17]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 68:17]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 68:17]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 68:17]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 68:17]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 68:17]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 68:17]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 68:17]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 68:17]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 68:17]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 68:17]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 68:17]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 68:17]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 68:17]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 68:17]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 68:17]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 68:17]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 68:17]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 68:17]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 68:17]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 68:17]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 68:17]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 68:17]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 68:17]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 68:17]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 68:17]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 68:17]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 68:17]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 68:17]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 68:17]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 68:17]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 68:17]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 68:17]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 68:17]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 68:17]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 68:17]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 68:17]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 68:17]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 68:17]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 68:17]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 68:17]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 68:17]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 68:17]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 68:17]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 68:17]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 68:17]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 68:17]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 68:17]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 68:17]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 68:17]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 68:17]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 68:17]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 68:17]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 68:17]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 68:17]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 68:17]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 68:17]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 68:17]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 68:17]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 68:17]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 68:17]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 68:17]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 68:17]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 68:17]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 68:17]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 68:17]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 68:17]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 68:17]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 68:17]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 68:17]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 68:17]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 68:17]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 68:17]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 68:17]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 68:17]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 68:17]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 68:17]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 68:17]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 68:17]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 68:17]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 68:17]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 68:17]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 68:17]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 68:17]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 68:17]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 68:17]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 68:17]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 68:17]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 68:17]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 68:17]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher.scala 68:17]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher.scala 68:17]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher.scala 68:17]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher.scala 68:17]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher.scala 68:17]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher.scala 68:17]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher.scala 68:17]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher.scala 68:17]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher.scala 68:17]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher.scala 68:17]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher.scala 68:17]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher.scala 68:17]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher.scala 68:17]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher.scala 68:17]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher.scala 68:17]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher.scala 68:17]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher.scala 68:17]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher.scala 68:17]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher.scala 68:17]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher.scala 68:17]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher.scala 68:17]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher.scala 68:17]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher.scala 68:17]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher.scala 68:17]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher.scala 68:17]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher.scala 68:17]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher.scala 68:17]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher.scala 68:17]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher.scala 68:17]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher.scala 68:17]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher.scala 68:17]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher.scala 68:17]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher.scala 68:17]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher.scala 68:17]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher.scala 68:17]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher.scala 68:17]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher.scala 68:17]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher.scala 68:17]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher.scala 68:17]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher.scala 68:17]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher.scala 68:17]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher.scala 68:17]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher.scala 68:17]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher.scala 68:17]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher.scala 68:17]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher.scala 68:17]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher.scala 68:17]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher.scala 68:17]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher.scala 68:17]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher.scala 68:17]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher.scala 68:17]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher.scala 68:17]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher.scala 68:17]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher.scala 68:17]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher.scala 68:17]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher.scala 68:17]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher.scala 68:17]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher.scala 68:17]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher.scala 68:17]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher.scala 68:17]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher.scala 68:17]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher.scala 68:17]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher.scala 68:17]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher.scala 68:17]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[matcher.scala 68:17]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[matcher.scala 68:17]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[matcher.scala 68:17]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[matcher.scala 68:17]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[matcher.scala 68:17]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[matcher.scala 68:17]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[matcher.scala 68:17]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[matcher.scala 68:17]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[matcher.scala 68:17]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[matcher.scala 68:17]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[matcher.scala 68:17]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[matcher.scala 68:17]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[matcher.scala 68:17]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[matcher.scala 68:17]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[matcher.scala 68:17]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[matcher.scala 68:17]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[matcher.scala 68:17]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[matcher.scala 68:17]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[matcher.scala 68:17]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[matcher.scala 68:17]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[matcher.scala 68:17]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[matcher.scala 68:17]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[matcher.scala 68:17]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[matcher.scala 68:17]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[matcher.scala 68:17]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[matcher.scala 68:17]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[matcher.scala 68:17]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[matcher.scala 68:17]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[matcher.scala 68:17]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[matcher.scala 68:17]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[matcher.scala 68:17]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[matcher.scala 68:17]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[matcher.scala 68:17]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[matcher.scala 68:17]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[matcher.scala 68:17]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[matcher.scala 68:17]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[matcher.scala 68:17]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[matcher.scala 68:17]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[matcher.scala 68:17]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[matcher.scala 68:17]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[matcher.scala 68:17]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[matcher.scala 68:17]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[matcher.scala 68:17]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[matcher.scala 68:17]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[matcher.scala 68:17]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[matcher.scala 68:17]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[matcher.scala 68:17]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[matcher.scala 68:17]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[matcher.scala 68:17]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[matcher.scala 68:17]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[matcher.scala 68:17]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[matcher.scala 68:17]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[matcher.scala 68:17]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[matcher.scala 68:17]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[matcher.scala 68:17]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[matcher.scala 68:17]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[matcher.scala 68:17]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[matcher.scala 68:17]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[matcher.scala 68:17]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[matcher.scala 68:17]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[matcher.scala 68:17]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[matcher.scala 68:17]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[matcher.scala 68:17]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[matcher.scala 68:17]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[matcher.scala 68:17]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[matcher.scala 68:17]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[matcher.scala 68:17]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[matcher.scala 68:17]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[matcher.scala 68:17]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[matcher.scala 68:17]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[matcher.scala 68:17]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[matcher.scala 68:17]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[matcher.scala 68:17]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[matcher.scala 68:17]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[matcher.scala 68:17]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[matcher.scala 68:17]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[matcher.scala 68:17]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[matcher.scala 68:17]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[matcher.scala 68:17]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[matcher.scala 68:17]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[matcher.scala 68:17]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[matcher.scala 68:17]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[matcher.scala 68:17]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[matcher.scala 68:17]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[matcher.scala 68:17]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[matcher.scala 68:17]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[matcher.scala 68:17]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[matcher.scala 68:17]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[matcher.scala 68:17]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[matcher.scala 68:17]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[matcher.scala 68:17]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[matcher.scala 68:17]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[matcher.scala 68:17]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[matcher.scala 68:17]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[matcher.scala 68:17]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[matcher.scala 68:17]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 68:17]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 68:17]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 68:17]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 68:17]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 68:17]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 68:17]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 68:17]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 68:17]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 68:17]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 68:17]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 68:17]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 68:17]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 68:17]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 68:17]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 68:17]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 68:17]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 68:17]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 68:17]
    key_offset <= io_key_offset_in; // @[matcher.scala 72:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_header_0 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  phv_header_1 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  phv_header_2 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  phv_header_3 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  phv_header_4 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  phv_header_5 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  phv_header_6 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  phv_header_7 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  phv_header_8 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  phv_header_9 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  phv_header_10 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  phv_header_11 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  phv_header_12 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  phv_header_13 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  phv_header_14 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  phv_header_15 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  phv_next_config_id = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  key_offset = _RAND_274[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
