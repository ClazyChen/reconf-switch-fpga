module MatchGetKeyRaw(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [7:0]  io_key_config_0_key_length,
  input  [7:0]  io_key_config_1_key_length,
  input  [7:0]  io_key_offset_in,
  output [1:0]  io_bias_out,
  output [7:0]  io_match_key_bytes_0,
  output [7:0]  io_match_key_bytes_1,
  output [7:0]  io_match_key_bytes_2,
  output [7:0]  io_match_key_bytes_3,
  output [7:0]  io_match_key_bytes_4,
  output [7:0]  io_match_key_bytes_5,
  output [7:0]  io_match_key_bytes_6,
  output [7:0]  io_match_key_bytes_7,
  output [7:0]  io_match_key_bytes_8,
  output [7:0]  io_match_key_bytes_9,
  output [7:0]  io_match_key_bytes_10,
  output [7:0]  io_match_key_bytes_11,
  output [7:0]  io_match_key_bytes_12,
  output [7:0]  io_match_key_bytes_13,
  output [7:0]  io_match_key_bytes_14,
  output [7:0]  io_match_key_bytes_15,
  output [7:0]  io_match_key_bytes_16,
  output [7:0]  io_match_key_bytes_17,
  output [7:0]  io_match_key_bytes_18,
  output [7:0]  io_match_key_bytes_19,
  output [7:0]  io_match_key_bytes_20,
  output [7:0]  io_match_key_bytes_21,
  output [7:0]  io_match_key_bytes_22,
  output [7:0]  io_match_key_bytes_23
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher.scala 67:26]
  reg [7:0] phv_data_1; // @[matcher.scala 67:26]
  reg [7:0] phv_data_2; // @[matcher.scala 67:26]
  reg [7:0] phv_data_3; // @[matcher.scala 67:26]
  reg [7:0] phv_data_4; // @[matcher.scala 67:26]
  reg [7:0] phv_data_5; // @[matcher.scala 67:26]
  reg [7:0] phv_data_6; // @[matcher.scala 67:26]
  reg [7:0] phv_data_7; // @[matcher.scala 67:26]
  reg [7:0] phv_data_8; // @[matcher.scala 67:26]
  reg [7:0] phv_data_9; // @[matcher.scala 67:26]
  reg [7:0] phv_data_10; // @[matcher.scala 67:26]
  reg [7:0] phv_data_11; // @[matcher.scala 67:26]
  reg [7:0] phv_data_12; // @[matcher.scala 67:26]
  reg [7:0] phv_data_13; // @[matcher.scala 67:26]
  reg [7:0] phv_data_14; // @[matcher.scala 67:26]
  reg [7:0] phv_data_15; // @[matcher.scala 67:26]
  reg [7:0] phv_data_16; // @[matcher.scala 67:26]
  reg [7:0] phv_data_17; // @[matcher.scala 67:26]
  reg [7:0] phv_data_18; // @[matcher.scala 67:26]
  reg [7:0] phv_data_19; // @[matcher.scala 67:26]
  reg [7:0] phv_data_20; // @[matcher.scala 67:26]
  reg [7:0] phv_data_21; // @[matcher.scala 67:26]
  reg [7:0] phv_data_22; // @[matcher.scala 67:26]
  reg [7:0] phv_data_23; // @[matcher.scala 67:26]
  reg [7:0] phv_data_24; // @[matcher.scala 67:26]
  reg [7:0] phv_data_25; // @[matcher.scala 67:26]
  reg [7:0] phv_data_26; // @[matcher.scala 67:26]
  reg [7:0] phv_data_27; // @[matcher.scala 67:26]
  reg [7:0] phv_data_28; // @[matcher.scala 67:26]
  reg [7:0] phv_data_29; // @[matcher.scala 67:26]
  reg [7:0] phv_data_30; // @[matcher.scala 67:26]
  reg [7:0] phv_data_31; // @[matcher.scala 67:26]
  reg [7:0] phv_data_32; // @[matcher.scala 67:26]
  reg [7:0] phv_data_33; // @[matcher.scala 67:26]
  reg [7:0] phv_data_34; // @[matcher.scala 67:26]
  reg [7:0] phv_data_35; // @[matcher.scala 67:26]
  reg [7:0] phv_data_36; // @[matcher.scala 67:26]
  reg [7:0] phv_data_37; // @[matcher.scala 67:26]
  reg [7:0] phv_data_38; // @[matcher.scala 67:26]
  reg [7:0] phv_data_39; // @[matcher.scala 67:26]
  reg [7:0] phv_data_40; // @[matcher.scala 67:26]
  reg [7:0] phv_data_41; // @[matcher.scala 67:26]
  reg [7:0] phv_data_42; // @[matcher.scala 67:26]
  reg [7:0] phv_data_43; // @[matcher.scala 67:26]
  reg [7:0] phv_data_44; // @[matcher.scala 67:26]
  reg [7:0] phv_data_45; // @[matcher.scala 67:26]
  reg [7:0] phv_data_46; // @[matcher.scala 67:26]
  reg [7:0] phv_data_47; // @[matcher.scala 67:26]
  reg [7:0] phv_data_48; // @[matcher.scala 67:26]
  reg [7:0] phv_data_49; // @[matcher.scala 67:26]
  reg [7:0] phv_data_50; // @[matcher.scala 67:26]
  reg [7:0] phv_data_51; // @[matcher.scala 67:26]
  reg [7:0] phv_data_52; // @[matcher.scala 67:26]
  reg [7:0] phv_data_53; // @[matcher.scala 67:26]
  reg [7:0] phv_data_54; // @[matcher.scala 67:26]
  reg [7:0] phv_data_55; // @[matcher.scala 67:26]
  reg [7:0] phv_data_56; // @[matcher.scala 67:26]
  reg [7:0] phv_data_57; // @[matcher.scala 67:26]
  reg [7:0] phv_data_58; // @[matcher.scala 67:26]
  reg [7:0] phv_data_59; // @[matcher.scala 67:26]
  reg [7:0] phv_data_60; // @[matcher.scala 67:26]
  reg [7:0] phv_data_61; // @[matcher.scala 67:26]
  reg [7:0] phv_data_62; // @[matcher.scala 67:26]
  reg [7:0] phv_data_63; // @[matcher.scala 67:26]
  reg [7:0] phv_data_64; // @[matcher.scala 67:26]
  reg [7:0] phv_data_65; // @[matcher.scala 67:26]
  reg [7:0] phv_data_66; // @[matcher.scala 67:26]
  reg [7:0] phv_data_67; // @[matcher.scala 67:26]
  reg [7:0] phv_data_68; // @[matcher.scala 67:26]
  reg [7:0] phv_data_69; // @[matcher.scala 67:26]
  reg [7:0] phv_data_70; // @[matcher.scala 67:26]
  reg [7:0] phv_data_71; // @[matcher.scala 67:26]
  reg [7:0] phv_data_72; // @[matcher.scala 67:26]
  reg [7:0] phv_data_73; // @[matcher.scala 67:26]
  reg [7:0] phv_data_74; // @[matcher.scala 67:26]
  reg [7:0] phv_data_75; // @[matcher.scala 67:26]
  reg [7:0] phv_data_76; // @[matcher.scala 67:26]
  reg [7:0] phv_data_77; // @[matcher.scala 67:26]
  reg [7:0] phv_data_78; // @[matcher.scala 67:26]
  reg [7:0] phv_data_79; // @[matcher.scala 67:26]
  reg [7:0] phv_data_80; // @[matcher.scala 67:26]
  reg [7:0] phv_data_81; // @[matcher.scala 67:26]
  reg [7:0] phv_data_82; // @[matcher.scala 67:26]
  reg [7:0] phv_data_83; // @[matcher.scala 67:26]
  reg [7:0] phv_data_84; // @[matcher.scala 67:26]
  reg [7:0] phv_data_85; // @[matcher.scala 67:26]
  reg [7:0] phv_data_86; // @[matcher.scala 67:26]
  reg [7:0] phv_data_87; // @[matcher.scala 67:26]
  reg [7:0] phv_data_88; // @[matcher.scala 67:26]
  reg [7:0] phv_data_89; // @[matcher.scala 67:26]
  reg [7:0] phv_data_90; // @[matcher.scala 67:26]
  reg [7:0] phv_data_91; // @[matcher.scala 67:26]
  reg [7:0] phv_data_92; // @[matcher.scala 67:26]
  reg [7:0] phv_data_93; // @[matcher.scala 67:26]
  reg [7:0] phv_data_94; // @[matcher.scala 67:26]
  reg [7:0] phv_data_95; // @[matcher.scala 67:26]
  reg [7:0] phv_data_96; // @[matcher.scala 67:26]
  reg [7:0] phv_data_97; // @[matcher.scala 67:26]
  reg [7:0] phv_data_98; // @[matcher.scala 67:26]
  reg [7:0] phv_data_99; // @[matcher.scala 67:26]
  reg [7:0] phv_data_100; // @[matcher.scala 67:26]
  reg [7:0] phv_data_101; // @[matcher.scala 67:26]
  reg [7:0] phv_data_102; // @[matcher.scala 67:26]
  reg [7:0] phv_data_103; // @[matcher.scala 67:26]
  reg [7:0] phv_data_104; // @[matcher.scala 67:26]
  reg [7:0] phv_data_105; // @[matcher.scala 67:26]
  reg [7:0] phv_data_106; // @[matcher.scala 67:26]
  reg [7:0] phv_data_107; // @[matcher.scala 67:26]
  reg [7:0] phv_data_108; // @[matcher.scala 67:26]
  reg [7:0] phv_data_109; // @[matcher.scala 67:26]
  reg [7:0] phv_data_110; // @[matcher.scala 67:26]
  reg [7:0] phv_data_111; // @[matcher.scala 67:26]
  reg [7:0] phv_data_112; // @[matcher.scala 67:26]
  reg [7:0] phv_data_113; // @[matcher.scala 67:26]
  reg [7:0] phv_data_114; // @[matcher.scala 67:26]
  reg [7:0] phv_data_115; // @[matcher.scala 67:26]
  reg [7:0] phv_data_116; // @[matcher.scala 67:26]
  reg [7:0] phv_data_117; // @[matcher.scala 67:26]
  reg [7:0] phv_data_118; // @[matcher.scala 67:26]
  reg [7:0] phv_data_119; // @[matcher.scala 67:26]
  reg [7:0] phv_data_120; // @[matcher.scala 67:26]
  reg [7:0] phv_data_121; // @[matcher.scala 67:26]
  reg [7:0] phv_data_122; // @[matcher.scala 67:26]
  reg [7:0] phv_data_123; // @[matcher.scala 67:26]
  reg [7:0] phv_data_124; // @[matcher.scala 67:26]
  reg [7:0] phv_data_125; // @[matcher.scala 67:26]
  reg [7:0] phv_data_126; // @[matcher.scala 67:26]
  reg [7:0] phv_data_127; // @[matcher.scala 67:26]
  reg [7:0] phv_data_128; // @[matcher.scala 67:26]
  reg [7:0] phv_data_129; // @[matcher.scala 67:26]
  reg [7:0] phv_data_130; // @[matcher.scala 67:26]
  reg [7:0] phv_data_131; // @[matcher.scala 67:26]
  reg [7:0] phv_data_132; // @[matcher.scala 67:26]
  reg [7:0] phv_data_133; // @[matcher.scala 67:26]
  reg [7:0] phv_data_134; // @[matcher.scala 67:26]
  reg [7:0] phv_data_135; // @[matcher.scala 67:26]
  reg [7:0] phv_data_136; // @[matcher.scala 67:26]
  reg [7:0] phv_data_137; // @[matcher.scala 67:26]
  reg [7:0] phv_data_138; // @[matcher.scala 67:26]
  reg [7:0] phv_data_139; // @[matcher.scala 67:26]
  reg [7:0] phv_data_140; // @[matcher.scala 67:26]
  reg [7:0] phv_data_141; // @[matcher.scala 67:26]
  reg [7:0] phv_data_142; // @[matcher.scala 67:26]
  reg [7:0] phv_data_143; // @[matcher.scala 67:26]
  reg [7:0] phv_data_144; // @[matcher.scala 67:26]
  reg [7:0] phv_data_145; // @[matcher.scala 67:26]
  reg [7:0] phv_data_146; // @[matcher.scala 67:26]
  reg [7:0] phv_data_147; // @[matcher.scala 67:26]
  reg [7:0] phv_data_148; // @[matcher.scala 67:26]
  reg [7:0] phv_data_149; // @[matcher.scala 67:26]
  reg [7:0] phv_data_150; // @[matcher.scala 67:26]
  reg [7:0] phv_data_151; // @[matcher.scala 67:26]
  reg [7:0] phv_data_152; // @[matcher.scala 67:26]
  reg [7:0] phv_data_153; // @[matcher.scala 67:26]
  reg [7:0] phv_data_154; // @[matcher.scala 67:26]
  reg [7:0] phv_data_155; // @[matcher.scala 67:26]
  reg [7:0] phv_data_156; // @[matcher.scala 67:26]
  reg [7:0] phv_data_157; // @[matcher.scala 67:26]
  reg [7:0] phv_data_158; // @[matcher.scala 67:26]
  reg [7:0] phv_data_159; // @[matcher.scala 67:26]
  reg [7:0] phv_data_160; // @[matcher.scala 67:26]
  reg [7:0] phv_data_161; // @[matcher.scala 67:26]
  reg [7:0] phv_data_162; // @[matcher.scala 67:26]
  reg [7:0] phv_data_163; // @[matcher.scala 67:26]
  reg [7:0] phv_data_164; // @[matcher.scala 67:26]
  reg [7:0] phv_data_165; // @[matcher.scala 67:26]
  reg [7:0] phv_data_166; // @[matcher.scala 67:26]
  reg [7:0] phv_data_167; // @[matcher.scala 67:26]
  reg [7:0] phv_data_168; // @[matcher.scala 67:26]
  reg [7:0] phv_data_169; // @[matcher.scala 67:26]
  reg [7:0] phv_data_170; // @[matcher.scala 67:26]
  reg [7:0] phv_data_171; // @[matcher.scala 67:26]
  reg [7:0] phv_data_172; // @[matcher.scala 67:26]
  reg [7:0] phv_data_173; // @[matcher.scala 67:26]
  reg [7:0] phv_data_174; // @[matcher.scala 67:26]
  reg [7:0] phv_data_175; // @[matcher.scala 67:26]
  reg [7:0] phv_data_176; // @[matcher.scala 67:26]
  reg [7:0] phv_data_177; // @[matcher.scala 67:26]
  reg [7:0] phv_data_178; // @[matcher.scala 67:26]
  reg [7:0] phv_data_179; // @[matcher.scala 67:26]
  reg [7:0] phv_data_180; // @[matcher.scala 67:26]
  reg [7:0] phv_data_181; // @[matcher.scala 67:26]
  reg [7:0] phv_data_182; // @[matcher.scala 67:26]
  reg [7:0] phv_data_183; // @[matcher.scala 67:26]
  reg [7:0] phv_data_184; // @[matcher.scala 67:26]
  reg [7:0] phv_data_185; // @[matcher.scala 67:26]
  reg [7:0] phv_data_186; // @[matcher.scala 67:26]
  reg [7:0] phv_data_187; // @[matcher.scala 67:26]
  reg [7:0] phv_data_188; // @[matcher.scala 67:26]
  reg [7:0] phv_data_189; // @[matcher.scala 67:26]
  reg [7:0] phv_data_190; // @[matcher.scala 67:26]
  reg [7:0] phv_data_191; // @[matcher.scala 67:26]
  reg [7:0] phv_data_192; // @[matcher.scala 67:26]
  reg [7:0] phv_data_193; // @[matcher.scala 67:26]
  reg [7:0] phv_data_194; // @[matcher.scala 67:26]
  reg [7:0] phv_data_195; // @[matcher.scala 67:26]
  reg [7:0] phv_data_196; // @[matcher.scala 67:26]
  reg [7:0] phv_data_197; // @[matcher.scala 67:26]
  reg [7:0] phv_data_198; // @[matcher.scala 67:26]
  reg [7:0] phv_data_199; // @[matcher.scala 67:26]
  reg [7:0] phv_data_200; // @[matcher.scala 67:26]
  reg [7:0] phv_data_201; // @[matcher.scala 67:26]
  reg [7:0] phv_data_202; // @[matcher.scala 67:26]
  reg [7:0] phv_data_203; // @[matcher.scala 67:26]
  reg [7:0] phv_data_204; // @[matcher.scala 67:26]
  reg [7:0] phv_data_205; // @[matcher.scala 67:26]
  reg [7:0] phv_data_206; // @[matcher.scala 67:26]
  reg [7:0] phv_data_207; // @[matcher.scala 67:26]
  reg [7:0] phv_data_208; // @[matcher.scala 67:26]
  reg [7:0] phv_data_209; // @[matcher.scala 67:26]
  reg [7:0] phv_data_210; // @[matcher.scala 67:26]
  reg [7:0] phv_data_211; // @[matcher.scala 67:26]
  reg [7:0] phv_data_212; // @[matcher.scala 67:26]
  reg [7:0] phv_data_213; // @[matcher.scala 67:26]
  reg [7:0] phv_data_214; // @[matcher.scala 67:26]
  reg [7:0] phv_data_215; // @[matcher.scala 67:26]
  reg [7:0] phv_data_216; // @[matcher.scala 67:26]
  reg [7:0] phv_data_217; // @[matcher.scala 67:26]
  reg [7:0] phv_data_218; // @[matcher.scala 67:26]
  reg [7:0] phv_data_219; // @[matcher.scala 67:26]
  reg [7:0] phv_data_220; // @[matcher.scala 67:26]
  reg [7:0] phv_data_221; // @[matcher.scala 67:26]
  reg [7:0] phv_data_222; // @[matcher.scala 67:26]
  reg [7:0] phv_data_223; // @[matcher.scala 67:26]
  reg [7:0] phv_data_224; // @[matcher.scala 67:26]
  reg [7:0] phv_data_225; // @[matcher.scala 67:26]
  reg [7:0] phv_data_226; // @[matcher.scala 67:26]
  reg [7:0] phv_data_227; // @[matcher.scala 67:26]
  reg [7:0] phv_data_228; // @[matcher.scala 67:26]
  reg [7:0] phv_data_229; // @[matcher.scala 67:26]
  reg [7:0] phv_data_230; // @[matcher.scala 67:26]
  reg [7:0] phv_data_231; // @[matcher.scala 67:26]
  reg [7:0] phv_data_232; // @[matcher.scala 67:26]
  reg [7:0] phv_data_233; // @[matcher.scala 67:26]
  reg [7:0] phv_data_234; // @[matcher.scala 67:26]
  reg [7:0] phv_data_235; // @[matcher.scala 67:26]
  reg [7:0] phv_data_236; // @[matcher.scala 67:26]
  reg [7:0] phv_data_237; // @[matcher.scala 67:26]
  reg [7:0] phv_data_238; // @[matcher.scala 67:26]
  reg [7:0] phv_data_239; // @[matcher.scala 67:26]
  reg [7:0] phv_data_240; // @[matcher.scala 67:26]
  reg [7:0] phv_data_241; // @[matcher.scala 67:26]
  reg [7:0] phv_data_242; // @[matcher.scala 67:26]
  reg [7:0] phv_data_243; // @[matcher.scala 67:26]
  reg [7:0] phv_data_244; // @[matcher.scala 67:26]
  reg [7:0] phv_data_245; // @[matcher.scala 67:26]
  reg [7:0] phv_data_246; // @[matcher.scala 67:26]
  reg [7:0] phv_data_247; // @[matcher.scala 67:26]
  reg [7:0] phv_data_248; // @[matcher.scala 67:26]
  reg [7:0] phv_data_249; // @[matcher.scala 67:26]
  reg [7:0] phv_data_250; // @[matcher.scala 67:26]
  reg [7:0] phv_data_251; // @[matcher.scala 67:26]
  reg [7:0] phv_data_252; // @[matcher.scala 67:26]
  reg [7:0] phv_data_253; // @[matcher.scala 67:26]
  reg [7:0] phv_data_254; // @[matcher.scala 67:26]
  reg [7:0] phv_data_255; // @[matcher.scala 67:26]
  reg [7:0] phv_data_256; // @[matcher.scala 67:26]
  reg [7:0] phv_data_257; // @[matcher.scala 67:26]
  reg [7:0] phv_data_258; // @[matcher.scala 67:26]
  reg [7:0] phv_data_259; // @[matcher.scala 67:26]
  reg [7:0] phv_data_260; // @[matcher.scala 67:26]
  reg [7:0] phv_data_261; // @[matcher.scala 67:26]
  reg [7:0] phv_data_262; // @[matcher.scala 67:26]
  reg [7:0] phv_data_263; // @[matcher.scala 67:26]
  reg [7:0] phv_data_264; // @[matcher.scala 67:26]
  reg [7:0] phv_data_265; // @[matcher.scala 67:26]
  reg [7:0] phv_data_266; // @[matcher.scala 67:26]
  reg [7:0] phv_data_267; // @[matcher.scala 67:26]
  reg [7:0] phv_data_268; // @[matcher.scala 67:26]
  reg [7:0] phv_data_269; // @[matcher.scala 67:26]
  reg [7:0] phv_data_270; // @[matcher.scala 67:26]
  reg [7:0] phv_data_271; // @[matcher.scala 67:26]
  reg [7:0] phv_data_272; // @[matcher.scala 67:26]
  reg [7:0] phv_data_273; // @[matcher.scala 67:26]
  reg [7:0] phv_data_274; // @[matcher.scala 67:26]
  reg [7:0] phv_data_275; // @[matcher.scala 67:26]
  reg [7:0] phv_data_276; // @[matcher.scala 67:26]
  reg [7:0] phv_data_277; // @[matcher.scala 67:26]
  reg [7:0] phv_data_278; // @[matcher.scala 67:26]
  reg [7:0] phv_data_279; // @[matcher.scala 67:26]
  reg [7:0] phv_data_280; // @[matcher.scala 67:26]
  reg [7:0] phv_data_281; // @[matcher.scala 67:26]
  reg [7:0] phv_data_282; // @[matcher.scala 67:26]
  reg [7:0] phv_data_283; // @[matcher.scala 67:26]
  reg [7:0] phv_data_284; // @[matcher.scala 67:26]
  reg [7:0] phv_data_285; // @[matcher.scala 67:26]
  reg [7:0] phv_data_286; // @[matcher.scala 67:26]
  reg [7:0] phv_data_287; // @[matcher.scala 67:26]
  reg [7:0] phv_data_288; // @[matcher.scala 67:26]
  reg [7:0] phv_data_289; // @[matcher.scala 67:26]
  reg [7:0] phv_data_290; // @[matcher.scala 67:26]
  reg [7:0] phv_data_291; // @[matcher.scala 67:26]
  reg [7:0] phv_data_292; // @[matcher.scala 67:26]
  reg [7:0] phv_data_293; // @[matcher.scala 67:26]
  reg [7:0] phv_data_294; // @[matcher.scala 67:26]
  reg [7:0] phv_data_295; // @[matcher.scala 67:26]
  reg [7:0] phv_data_296; // @[matcher.scala 67:26]
  reg [7:0] phv_data_297; // @[matcher.scala 67:26]
  reg [7:0] phv_data_298; // @[matcher.scala 67:26]
  reg [7:0] phv_data_299; // @[matcher.scala 67:26]
  reg [7:0] phv_data_300; // @[matcher.scala 67:26]
  reg [7:0] phv_data_301; // @[matcher.scala 67:26]
  reg [7:0] phv_data_302; // @[matcher.scala 67:26]
  reg [7:0] phv_data_303; // @[matcher.scala 67:26]
  reg [7:0] phv_data_304; // @[matcher.scala 67:26]
  reg [7:0] phv_data_305; // @[matcher.scala 67:26]
  reg [7:0] phv_data_306; // @[matcher.scala 67:26]
  reg [7:0] phv_data_307; // @[matcher.scala 67:26]
  reg [7:0] phv_data_308; // @[matcher.scala 67:26]
  reg [7:0] phv_data_309; // @[matcher.scala 67:26]
  reg [7:0] phv_data_310; // @[matcher.scala 67:26]
  reg [7:0] phv_data_311; // @[matcher.scala 67:26]
  reg [7:0] phv_data_312; // @[matcher.scala 67:26]
  reg [7:0] phv_data_313; // @[matcher.scala 67:26]
  reg [7:0] phv_data_314; // @[matcher.scala 67:26]
  reg [7:0] phv_data_315; // @[matcher.scala 67:26]
  reg [7:0] phv_data_316; // @[matcher.scala 67:26]
  reg [7:0] phv_data_317; // @[matcher.scala 67:26]
  reg [7:0] phv_data_318; // @[matcher.scala 67:26]
  reg [7:0] phv_data_319; // @[matcher.scala 67:26]
  reg [7:0] phv_data_320; // @[matcher.scala 67:26]
  reg [7:0] phv_data_321; // @[matcher.scala 67:26]
  reg [7:0] phv_data_322; // @[matcher.scala 67:26]
  reg [7:0] phv_data_323; // @[matcher.scala 67:26]
  reg [7:0] phv_data_324; // @[matcher.scala 67:26]
  reg [7:0] phv_data_325; // @[matcher.scala 67:26]
  reg [7:0] phv_data_326; // @[matcher.scala 67:26]
  reg [7:0] phv_data_327; // @[matcher.scala 67:26]
  reg [7:0] phv_data_328; // @[matcher.scala 67:26]
  reg [7:0] phv_data_329; // @[matcher.scala 67:26]
  reg [7:0] phv_data_330; // @[matcher.scala 67:26]
  reg [7:0] phv_data_331; // @[matcher.scala 67:26]
  reg [7:0] phv_data_332; // @[matcher.scala 67:26]
  reg [7:0] phv_data_333; // @[matcher.scala 67:26]
  reg [7:0] phv_data_334; // @[matcher.scala 67:26]
  reg [7:0] phv_data_335; // @[matcher.scala 67:26]
  reg [7:0] phv_data_336; // @[matcher.scala 67:26]
  reg [7:0] phv_data_337; // @[matcher.scala 67:26]
  reg [7:0] phv_data_338; // @[matcher.scala 67:26]
  reg [7:0] phv_data_339; // @[matcher.scala 67:26]
  reg [7:0] phv_data_340; // @[matcher.scala 67:26]
  reg [7:0] phv_data_341; // @[matcher.scala 67:26]
  reg [7:0] phv_data_342; // @[matcher.scala 67:26]
  reg [7:0] phv_data_343; // @[matcher.scala 67:26]
  reg [7:0] phv_data_344; // @[matcher.scala 67:26]
  reg [7:0] phv_data_345; // @[matcher.scala 67:26]
  reg [7:0] phv_data_346; // @[matcher.scala 67:26]
  reg [7:0] phv_data_347; // @[matcher.scala 67:26]
  reg [7:0] phv_data_348; // @[matcher.scala 67:26]
  reg [7:0] phv_data_349; // @[matcher.scala 67:26]
  reg [7:0] phv_data_350; // @[matcher.scala 67:26]
  reg [7:0] phv_data_351; // @[matcher.scala 67:26]
  reg [7:0] phv_data_352; // @[matcher.scala 67:26]
  reg [7:0] phv_data_353; // @[matcher.scala 67:26]
  reg [7:0] phv_data_354; // @[matcher.scala 67:26]
  reg [7:0] phv_data_355; // @[matcher.scala 67:26]
  reg [7:0] phv_data_356; // @[matcher.scala 67:26]
  reg [7:0] phv_data_357; // @[matcher.scala 67:26]
  reg [7:0] phv_data_358; // @[matcher.scala 67:26]
  reg [7:0] phv_data_359; // @[matcher.scala 67:26]
  reg [7:0] phv_data_360; // @[matcher.scala 67:26]
  reg [7:0] phv_data_361; // @[matcher.scala 67:26]
  reg [7:0] phv_data_362; // @[matcher.scala 67:26]
  reg [7:0] phv_data_363; // @[matcher.scala 67:26]
  reg [7:0] phv_data_364; // @[matcher.scala 67:26]
  reg [7:0] phv_data_365; // @[matcher.scala 67:26]
  reg [7:0] phv_data_366; // @[matcher.scala 67:26]
  reg [7:0] phv_data_367; // @[matcher.scala 67:26]
  reg [7:0] phv_data_368; // @[matcher.scala 67:26]
  reg [7:0] phv_data_369; // @[matcher.scala 67:26]
  reg [7:0] phv_data_370; // @[matcher.scala 67:26]
  reg [7:0] phv_data_371; // @[matcher.scala 67:26]
  reg [7:0] phv_data_372; // @[matcher.scala 67:26]
  reg [7:0] phv_data_373; // @[matcher.scala 67:26]
  reg [7:0] phv_data_374; // @[matcher.scala 67:26]
  reg [7:0] phv_data_375; // @[matcher.scala 67:26]
  reg [7:0] phv_data_376; // @[matcher.scala 67:26]
  reg [7:0] phv_data_377; // @[matcher.scala 67:26]
  reg [7:0] phv_data_378; // @[matcher.scala 67:26]
  reg [7:0] phv_data_379; // @[matcher.scala 67:26]
  reg [7:0] phv_data_380; // @[matcher.scala 67:26]
  reg [7:0] phv_data_381; // @[matcher.scala 67:26]
  reg [7:0] phv_data_382; // @[matcher.scala 67:26]
  reg [7:0] phv_data_383; // @[matcher.scala 67:26]
  reg [7:0] phv_data_384; // @[matcher.scala 67:26]
  reg [7:0] phv_data_385; // @[matcher.scala 67:26]
  reg [7:0] phv_data_386; // @[matcher.scala 67:26]
  reg [7:0] phv_data_387; // @[matcher.scala 67:26]
  reg [7:0] phv_data_388; // @[matcher.scala 67:26]
  reg [7:0] phv_data_389; // @[matcher.scala 67:26]
  reg [7:0] phv_data_390; // @[matcher.scala 67:26]
  reg [7:0] phv_data_391; // @[matcher.scala 67:26]
  reg [7:0] phv_data_392; // @[matcher.scala 67:26]
  reg [7:0] phv_data_393; // @[matcher.scala 67:26]
  reg [7:0] phv_data_394; // @[matcher.scala 67:26]
  reg [7:0] phv_data_395; // @[matcher.scala 67:26]
  reg [7:0] phv_data_396; // @[matcher.scala 67:26]
  reg [7:0] phv_data_397; // @[matcher.scala 67:26]
  reg [7:0] phv_data_398; // @[matcher.scala 67:26]
  reg [7:0] phv_data_399; // @[matcher.scala 67:26]
  reg [7:0] phv_data_400; // @[matcher.scala 67:26]
  reg [7:0] phv_data_401; // @[matcher.scala 67:26]
  reg [7:0] phv_data_402; // @[matcher.scala 67:26]
  reg [7:0] phv_data_403; // @[matcher.scala 67:26]
  reg [7:0] phv_data_404; // @[matcher.scala 67:26]
  reg [7:0] phv_data_405; // @[matcher.scala 67:26]
  reg [7:0] phv_data_406; // @[matcher.scala 67:26]
  reg [7:0] phv_data_407; // @[matcher.scala 67:26]
  reg [7:0] phv_data_408; // @[matcher.scala 67:26]
  reg [7:0] phv_data_409; // @[matcher.scala 67:26]
  reg [7:0] phv_data_410; // @[matcher.scala 67:26]
  reg [7:0] phv_data_411; // @[matcher.scala 67:26]
  reg [7:0] phv_data_412; // @[matcher.scala 67:26]
  reg [7:0] phv_data_413; // @[matcher.scala 67:26]
  reg [7:0] phv_data_414; // @[matcher.scala 67:26]
  reg [7:0] phv_data_415; // @[matcher.scala 67:26]
  reg [7:0] phv_data_416; // @[matcher.scala 67:26]
  reg [7:0] phv_data_417; // @[matcher.scala 67:26]
  reg [7:0] phv_data_418; // @[matcher.scala 67:26]
  reg [7:0] phv_data_419; // @[matcher.scala 67:26]
  reg [7:0] phv_data_420; // @[matcher.scala 67:26]
  reg [7:0] phv_data_421; // @[matcher.scala 67:26]
  reg [7:0] phv_data_422; // @[matcher.scala 67:26]
  reg [7:0] phv_data_423; // @[matcher.scala 67:26]
  reg [7:0] phv_data_424; // @[matcher.scala 67:26]
  reg [7:0] phv_data_425; // @[matcher.scala 67:26]
  reg [7:0] phv_data_426; // @[matcher.scala 67:26]
  reg [7:0] phv_data_427; // @[matcher.scala 67:26]
  reg [7:0] phv_data_428; // @[matcher.scala 67:26]
  reg [7:0] phv_data_429; // @[matcher.scala 67:26]
  reg [7:0] phv_data_430; // @[matcher.scala 67:26]
  reg [7:0] phv_data_431; // @[matcher.scala 67:26]
  reg [7:0] phv_data_432; // @[matcher.scala 67:26]
  reg [7:0] phv_data_433; // @[matcher.scala 67:26]
  reg [7:0] phv_data_434; // @[matcher.scala 67:26]
  reg [7:0] phv_data_435; // @[matcher.scala 67:26]
  reg [7:0] phv_data_436; // @[matcher.scala 67:26]
  reg [7:0] phv_data_437; // @[matcher.scala 67:26]
  reg [7:0] phv_data_438; // @[matcher.scala 67:26]
  reg [7:0] phv_data_439; // @[matcher.scala 67:26]
  reg [7:0] phv_data_440; // @[matcher.scala 67:26]
  reg [7:0] phv_data_441; // @[matcher.scala 67:26]
  reg [7:0] phv_data_442; // @[matcher.scala 67:26]
  reg [7:0] phv_data_443; // @[matcher.scala 67:26]
  reg [7:0] phv_data_444; // @[matcher.scala 67:26]
  reg [7:0] phv_data_445; // @[matcher.scala 67:26]
  reg [7:0] phv_data_446; // @[matcher.scala 67:26]
  reg [7:0] phv_data_447; // @[matcher.scala 67:26]
  reg [7:0] phv_data_448; // @[matcher.scala 67:26]
  reg [7:0] phv_data_449; // @[matcher.scala 67:26]
  reg [7:0] phv_data_450; // @[matcher.scala 67:26]
  reg [7:0] phv_data_451; // @[matcher.scala 67:26]
  reg [7:0] phv_data_452; // @[matcher.scala 67:26]
  reg [7:0] phv_data_453; // @[matcher.scala 67:26]
  reg [7:0] phv_data_454; // @[matcher.scala 67:26]
  reg [7:0] phv_data_455; // @[matcher.scala 67:26]
  reg [7:0] phv_data_456; // @[matcher.scala 67:26]
  reg [7:0] phv_data_457; // @[matcher.scala 67:26]
  reg [7:0] phv_data_458; // @[matcher.scala 67:26]
  reg [7:0] phv_data_459; // @[matcher.scala 67:26]
  reg [7:0] phv_data_460; // @[matcher.scala 67:26]
  reg [7:0] phv_data_461; // @[matcher.scala 67:26]
  reg [7:0] phv_data_462; // @[matcher.scala 67:26]
  reg [7:0] phv_data_463; // @[matcher.scala 67:26]
  reg [7:0] phv_data_464; // @[matcher.scala 67:26]
  reg [7:0] phv_data_465; // @[matcher.scala 67:26]
  reg [7:0] phv_data_466; // @[matcher.scala 67:26]
  reg [7:0] phv_data_467; // @[matcher.scala 67:26]
  reg [7:0] phv_data_468; // @[matcher.scala 67:26]
  reg [7:0] phv_data_469; // @[matcher.scala 67:26]
  reg [7:0] phv_data_470; // @[matcher.scala 67:26]
  reg [7:0] phv_data_471; // @[matcher.scala 67:26]
  reg [7:0] phv_data_472; // @[matcher.scala 67:26]
  reg [7:0] phv_data_473; // @[matcher.scala 67:26]
  reg [7:0] phv_data_474; // @[matcher.scala 67:26]
  reg [7:0] phv_data_475; // @[matcher.scala 67:26]
  reg [7:0] phv_data_476; // @[matcher.scala 67:26]
  reg [7:0] phv_data_477; // @[matcher.scala 67:26]
  reg [7:0] phv_data_478; // @[matcher.scala 67:26]
  reg [7:0] phv_data_479; // @[matcher.scala 67:26]
  reg [7:0] phv_data_480; // @[matcher.scala 67:26]
  reg [7:0] phv_data_481; // @[matcher.scala 67:26]
  reg [7:0] phv_data_482; // @[matcher.scala 67:26]
  reg [7:0] phv_data_483; // @[matcher.scala 67:26]
  reg [7:0] phv_data_484; // @[matcher.scala 67:26]
  reg [7:0] phv_data_485; // @[matcher.scala 67:26]
  reg [7:0] phv_data_486; // @[matcher.scala 67:26]
  reg [7:0] phv_data_487; // @[matcher.scala 67:26]
  reg [7:0] phv_data_488; // @[matcher.scala 67:26]
  reg [7:0] phv_data_489; // @[matcher.scala 67:26]
  reg [7:0] phv_data_490; // @[matcher.scala 67:26]
  reg [7:0] phv_data_491; // @[matcher.scala 67:26]
  reg [7:0] phv_data_492; // @[matcher.scala 67:26]
  reg [7:0] phv_data_493; // @[matcher.scala 67:26]
  reg [7:0] phv_data_494; // @[matcher.scala 67:26]
  reg [7:0] phv_data_495; // @[matcher.scala 67:26]
  reg [7:0] phv_data_496; // @[matcher.scala 67:26]
  reg [7:0] phv_data_497; // @[matcher.scala 67:26]
  reg [7:0] phv_data_498; // @[matcher.scala 67:26]
  reg [7:0] phv_data_499; // @[matcher.scala 67:26]
  reg [7:0] phv_data_500; // @[matcher.scala 67:26]
  reg [7:0] phv_data_501; // @[matcher.scala 67:26]
  reg [7:0] phv_data_502; // @[matcher.scala 67:26]
  reg [7:0] phv_data_503; // @[matcher.scala 67:26]
  reg [7:0] phv_data_504; // @[matcher.scala 67:26]
  reg [7:0] phv_data_505; // @[matcher.scala 67:26]
  reg [7:0] phv_data_506; // @[matcher.scala 67:26]
  reg [7:0] phv_data_507; // @[matcher.scala 67:26]
  reg [7:0] phv_data_508; // @[matcher.scala 67:26]
  reg [7:0] phv_data_509; // @[matcher.scala 67:26]
  reg [7:0] phv_data_510; // @[matcher.scala 67:26]
  reg [7:0] phv_data_511; // @[matcher.scala 67:26]
  reg [15:0] phv_header_0; // @[matcher.scala 67:26]
  reg [15:0] phv_header_1; // @[matcher.scala 67:26]
  reg [15:0] phv_header_2; // @[matcher.scala 67:26]
  reg [15:0] phv_header_3; // @[matcher.scala 67:26]
  reg [15:0] phv_header_4; // @[matcher.scala 67:26]
  reg [15:0] phv_header_5; // @[matcher.scala 67:26]
  reg [15:0] phv_header_6; // @[matcher.scala 67:26]
  reg [15:0] phv_header_7; // @[matcher.scala 67:26]
  reg [15:0] phv_header_8; // @[matcher.scala 67:26]
  reg [15:0] phv_header_9; // @[matcher.scala 67:26]
  reg [15:0] phv_header_10; // @[matcher.scala 67:26]
  reg [15:0] phv_header_11; // @[matcher.scala 67:26]
  reg [15:0] phv_header_12; // @[matcher.scala 67:26]
  reg [15:0] phv_header_13; // @[matcher.scala 67:26]
  reg [15:0] phv_header_14; // @[matcher.scala 67:26]
  reg [15:0] phv_header_15; // @[matcher.scala 67:26]
  reg [7:0] phv_parse_current_state; // @[matcher.scala 67:26]
  reg [7:0] phv_parse_current_offset; // @[matcher.scala 67:26]
  reg [15:0] phv_parse_transition_field; // @[matcher.scala 67:26]
  reg [3:0] phv_next_processor_id; // @[matcher.scala 67:26]
  reg  phv_next_config_id; // @[matcher.scala 67:26]
  reg  phv_is_valid_processor; // @[matcher.scala 67:26]
  reg [7:0] key_offset; // @[matcher.scala 71:33]
  wire [5:0] read_key_offset_hi = key_offset[7:2]; // @[matcher.scala 73:49]
  wire [7:0] read_key_offset = {read_key_offset_hi,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_6 = phv_next_config_id ? io_key_config_1_key_length : io_key_config_0_key_length; // @[matcher.scala 84:85 matcher.scala 84:85]
  wire [7:0] end_offset = _GEN_6 + key_offset; // @[matcher.scala 84:85]
  wire [8:0] _local_offset_T = {{1'd0}, read_key_offset}; // @[matcher.scala 87:77]
  wire [7:0] local_offset = _local_offset_T[7:0]; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_0_hi = local_offset[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_0_T = {match_key_qbytes_0_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_0_T_1 = {match_key_qbytes_0_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_0_T_2 = {match_key_qbytes_0_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_9 = 8'h1 == _match_key_qbytes_0_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10 = 8'h2 == _match_key_qbytes_0_T_2 ? phv_data_2 : _GEN_9; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11 = 8'h3 == _match_key_qbytes_0_T_2 ? phv_data_3 : _GEN_10; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12 = 8'h4 == _match_key_qbytes_0_T_2 ? phv_data_4 : _GEN_11; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_13 = 8'h5 == _match_key_qbytes_0_T_2 ? phv_data_5 : _GEN_12; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_14 = 8'h6 == _match_key_qbytes_0_T_2 ? phv_data_6 : _GEN_13; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_15 = 8'h7 == _match_key_qbytes_0_T_2 ? phv_data_7 : _GEN_14; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_16 = 8'h8 == _match_key_qbytes_0_T_2 ? phv_data_8 : _GEN_15; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_17 = 8'h9 == _match_key_qbytes_0_T_2 ? phv_data_9 : _GEN_16; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_18 = 8'ha == _match_key_qbytes_0_T_2 ? phv_data_10 : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_19 = 8'hb == _match_key_qbytes_0_T_2 ? phv_data_11 : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_20 = 8'hc == _match_key_qbytes_0_T_2 ? phv_data_12 : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_21 = 8'hd == _match_key_qbytes_0_T_2 ? phv_data_13 : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_22 = 8'he == _match_key_qbytes_0_T_2 ? phv_data_14 : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_23 = 8'hf == _match_key_qbytes_0_T_2 ? phv_data_15 : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_24 = 8'h10 == _match_key_qbytes_0_T_2 ? phv_data_16 : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_25 = 8'h11 == _match_key_qbytes_0_T_2 ? phv_data_17 : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_26 = 8'h12 == _match_key_qbytes_0_T_2 ? phv_data_18 : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_27 = 8'h13 == _match_key_qbytes_0_T_2 ? phv_data_19 : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_28 = 8'h14 == _match_key_qbytes_0_T_2 ? phv_data_20 : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_29 = 8'h15 == _match_key_qbytes_0_T_2 ? phv_data_21 : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_30 = 8'h16 == _match_key_qbytes_0_T_2 ? phv_data_22 : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_31 = 8'h17 == _match_key_qbytes_0_T_2 ? phv_data_23 : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_32 = 8'h18 == _match_key_qbytes_0_T_2 ? phv_data_24 : _GEN_31; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_33 = 8'h19 == _match_key_qbytes_0_T_2 ? phv_data_25 : _GEN_32; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_34 = 8'h1a == _match_key_qbytes_0_T_2 ? phv_data_26 : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_35 = 8'h1b == _match_key_qbytes_0_T_2 ? phv_data_27 : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_36 = 8'h1c == _match_key_qbytes_0_T_2 ? phv_data_28 : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_37 = 8'h1d == _match_key_qbytes_0_T_2 ? phv_data_29 : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_38 = 8'h1e == _match_key_qbytes_0_T_2 ? phv_data_30 : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_39 = 8'h1f == _match_key_qbytes_0_T_2 ? phv_data_31 : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_40 = 8'h20 == _match_key_qbytes_0_T_2 ? phv_data_32 : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_41 = 8'h21 == _match_key_qbytes_0_T_2 ? phv_data_33 : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_42 = 8'h22 == _match_key_qbytes_0_T_2 ? phv_data_34 : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_43 = 8'h23 == _match_key_qbytes_0_T_2 ? phv_data_35 : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_44 = 8'h24 == _match_key_qbytes_0_T_2 ? phv_data_36 : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_45 = 8'h25 == _match_key_qbytes_0_T_2 ? phv_data_37 : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_46 = 8'h26 == _match_key_qbytes_0_T_2 ? phv_data_38 : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_47 = 8'h27 == _match_key_qbytes_0_T_2 ? phv_data_39 : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_48 = 8'h28 == _match_key_qbytes_0_T_2 ? phv_data_40 : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_49 = 8'h29 == _match_key_qbytes_0_T_2 ? phv_data_41 : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_50 = 8'h2a == _match_key_qbytes_0_T_2 ? phv_data_42 : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 8'h2b == _match_key_qbytes_0_T_2 ? phv_data_43 : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 8'h2c == _match_key_qbytes_0_T_2 ? phv_data_44 : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 8'h2d == _match_key_qbytes_0_T_2 ? phv_data_45 : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 8'h2e == _match_key_qbytes_0_T_2 ? phv_data_46 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 8'h2f == _match_key_qbytes_0_T_2 ? phv_data_47 : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 8'h30 == _match_key_qbytes_0_T_2 ? phv_data_48 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 8'h31 == _match_key_qbytes_0_T_2 ? phv_data_49 : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 8'h32 == _match_key_qbytes_0_T_2 ? phv_data_50 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 8'h33 == _match_key_qbytes_0_T_2 ? phv_data_51 : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 8'h34 == _match_key_qbytes_0_T_2 ? phv_data_52 : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 8'h35 == _match_key_qbytes_0_T_2 ? phv_data_53 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 8'h36 == _match_key_qbytes_0_T_2 ? phv_data_54 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 8'h37 == _match_key_qbytes_0_T_2 ? phv_data_55 : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_64 = 8'h38 == _match_key_qbytes_0_T_2 ? phv_data_56 : _GEN_63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_65 = 8'h39 == _match_key_qbytes_0_T_2 ? phv_data_57 : _GEN_64; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_66 = 8'h3a == _match_key_qbytes_0_T_2 ? phv_data_58 : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_67 = 8'h3b == _match_key_qbytes_0_T_2 ? phv_data_59 : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_68 = 8'h3c == _match_key_qbytes_0_T_2 ? phv_data_60 : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_69 = 8'h3d == _match_key_qbytes_0_T_2 ? phv_data_61 : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_70 = 8'h3e == _match_key_qbytes_0_T_2 ? phv_data_62 : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_71 = 8'h3f == _match_key_qbytes_0_T_2 ? phv_data_63 : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_72 = 8'h40 == _match_key_qbytes_0_T_2 ? phv_data_64 : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_73 = 8'h41 == _match_key_qbytes_0_T_2 ? phv_data_65 : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_74 = 8'h42 == _match_key_qbytes_0_T_2 ? phv_data_66 : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_75 = 8'h43 == _match_key_qbytes_0_T_2 ? phv_data_67 : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_76 = 8'h44 == _match_key_qbytes_0_T_2 ? phv_data_68 : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_77 = 8'h45 == _match_key_qbytes_0_T_2 ? phv_data_69 : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_78 = 8'h46 == _match_key_qbytes_0_T_2 ? phv_data_70 : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_79 = 8'h47 == _match_key_qbytes_0_T_2 ? phv_data_71 : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_80 = 8'h48 == _match_key_qbytes_0_T_2 ? phv_data_72 : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_81 = 8'h49 == _match_key_qbytes_0_T_2 ? phv_data_73 : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_82 = 8'h4a == _match_key_qbytes_0_T_2 ? phv_data_74 : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_83 = 8'h4b == _match_key_qbytes_0_T_2 ? phv_data_75 : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_84 = 8'h4c == _match_key_qbytes_0_T_2 ? phv_data_76 : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_85 = 8'h4d == _match_key_qbytes_0_T_2 ? phv_data_77 : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_86 = 8'h4e == _match_key_qbytes_0_T_2 ? phv_data_78 : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_87 = 8'h4f == _match_key_qbytes_0_T_2 ? phv_data_79 : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_88 = 8'h50 == _match_key_qbytes_0_T_2 ? phv_data_80 : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_89 = 8'h51 == _match_key_qbytes_0_T_2 ? phv_data_81 : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_90 = 8'h52 == _match_key_qbytes_0_T_2 ? phv_data_82 : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_91 = 8'h53 == _match_key_qbytes_0_T_2 ? phv_data_83 : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_92 = 8'h54 == _match_key_qbytes_0_T_2 ? phv_data_84 : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_93 = 8'h55 == _match_key_qbytes_0_T_2 ? phv_data_85 : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_94 = 8'h56 == _match_key_qbytes_0_T_2 ? phv_data_86 : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_95 = 8'h57 == _match_key_qbytes_0_T_2 ? phv_data_87 : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_96 = 8'h58 == _match_key_qbytes_0_T_2 ? phv_data_88 : _GEN_95; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_97 = 8'h59 == _match_key_qbytes_0_T_2 ? phv_data_89 : _GEN_96; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_98 = 8'h5a == _match_key_qbytes_0_T_2 ? phv_data_90 : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_99 = 8'h5b == _match_key_qbytes_0_T_2 ? phv_data_91 : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_100 = 8'h5c == _match_key_qbytes_0_T_2 ? phv_data_92 : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_101 = 8'h5d == _match_key_qbytes_0_T_2 ? phv_data_93 : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_102 = 8'h5e == _match_key_qbytes_0_T_2 ? phv_data_94 : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_103 = 8'h5f == _match_key_qbytes_0_T_2 ? phv_data_95 : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_104 = 8'h60 == _match_key_qbytes_0_T_2 ? phv_data_96 : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_105 = 8'h61 == _match_key_qbytes_0_T_2 ? phv_data_97 : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_106 = 8'h62 == _match_key_qbytes_0_T_2 ? phv_data_98 : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_107 = 8'h63 == _match_key_qbytes_0_T_2 ? phv_data_99 : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_108 = 8'h64 == _match_key_qbytes_0_T_2 ? phv_data_100 : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_109 = 8'h65 == _match_key_qbytes_0_T_2 ? phv_data_101 : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_110 = 8'h66 == _match_key_qbytes_0_T_2 ? phv_data_102 : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_111 = 8'h67 == _match_key_qbytes_0_T_2 ? phv_data_103 : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_112 = 8'h68 == _match_key_qbytes_0_T_2 ? phv_data_104 : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_113 = 8'h69 == _match_key_qbytes_0_T_2 ? phv_data_105 : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_114 = 8'h6a == _match_key_qbytes_0_T_2 ? phv_data_106 : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_115 = 8'h6b == _match_key_qbytes_0_T_2 ? phv_data_107 : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_116 = 8'h6c == _match_key_qbytes_0_T_2 ? phv_data_108 : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_117 = 8'h6d == _match_key_qbytes_0_T_2 ? phv_data_109 : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_118 = 8'h6e == _match_key_qbytes_0_T_2 ? phv_data_110 : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_119 = 8'h6f == _match_key_qbytes_0_T_2 ? phv_data_111 : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_120 = 8'h70 == _match_key_qbytes_0_T_2 ? phv_data_112 : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_121 = 8'h71 == _match_key_qbytes_0_T_2 ? phv_data_113 : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_122 = 8'h72 == _match_key_qbytes_0_T_2 ? phv_data_114 : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_123 = 8'h73 == _match_key_qbytes_0_T_2 ? phv_data_115 : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_124 = 8'h74 == _match_key_qbytes_0_T_2 ? phv_data_116 : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_125 = 8'h75 == _match_key_qbytes_0_T_2 ? phv_data_117 : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_126 = 8'h76 == _match_key_qbytes_0_T_2 ? phv_data_118 : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_127 = 8'h77 == _match_key_qbytes_0_T_2 ? phv_data_119 : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_128 = 8'h78 == _match_key_qbytes_0_T_2 ? phv_data_120 : _GEN_127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_129 = 8'h79 == _match_key_qbytes_0_T_2 ? phv_data_121 : _GEN_128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_130 = 8'h7a == _match_key_qbytes_0_T_2 ? phv_data_122 : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_131 = 8'h7b == _match_key_qbytes_0_T_2 ? phv_data_123 : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_132 = 8'h7c == _match_key_qbytes_0_T_2 ? phv_data_124 : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_133 = 8'h7d == _match_key_qbytes_0_T_2 ? phv_data_125 : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_134 = 8'h7e == _match_key_qbytes_0_T_2 ? phv_data_126 : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_135 = 8'h7f == _match_key_qbytes_0_T_2 ? phv_data_127 : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_136 = 8'h80 == _match_key_qbytes_0_T_2 ? phv_data_128 : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_137 = 8'h81 == _match_key_qbytes_0_T_2 ? phv_data_129 : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_138 = 8'h82 == _match_key_qbytes_0_T_2 ? phv_data_130 : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_139 = 8'h83 == _match_key_qbytes_0_T_2 ? phv_data_131 : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_140 = 8'h84 == _match_key_qbytes_0_T_2 ? phv_data_132 : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_141 = 8'h85 == _match_key_qbytes_0_T_2 ? phv_data_133 : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_142 = 8'h86 == _match_key_qbytes_0_T_2 ? phv_data_134 : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_143 = 8'h87 == _match_key_qbytes_0_T_2 ? phv_data_135 : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_144 = 8'h88 == _match_key_qbytes_0_T_2 ? phv_data_136 : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_145 = 8'h89 == _match_key_qbytes_0_T_2 ? phv_data_137 : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_146 = 8'h8a == _match_key_qbytes_0_T_2 ? phv_data_138 : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_147 = 8'h8b == _match_key_qbytes_0_T_2 ? phv_data_139 : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_148 = 8'h8c == _match_key_qbytes_0_T_2 ? phv_data_140 : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_149 = 8'h8d == _match_key_qbytes_0_T_2 ? phv_data_141 : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_150 = 8'h8e == _match_key_qbytes_0_T_2 ? phv_data_142 : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_151 = 8'h8f == _match_key_qbytes_0_T_2 ? phv_data_143 : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_152 = 8'h90 == _match_key_qbytes_0_T_2 ? phv_data_144 : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_153 = 8'h91 == _match_key_qbytes_0_T_2 ? phv_data_145 : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_154 = 8'h92 == _match_key_qbytes_0_T_2 ? phv_data_146 : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_155 = 8'h93 == _match_key_qbytes_0_T_2 ? phv_data_147 : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_156 = 8'h94 == _match_key_qbytes_0_T_2 ? phv_data_148 : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_157 = 8'h95 == _match_key_qbytes_0_T_2 ? phv_data_149 : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_158 = 8'h96 == _match_key_qbytes_0_T_2 ? phv_data_150 : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_159 = 8'h97 == _match_key_qbytes_0_T_2 ? phv_data_151 : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_160 = 8'h98 == _match_key_qbytes_0_T_2 ? phv_data_152 : _GEN_159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_161 = 8'h99 == _match_key_qbytes_0_T_2 ? phv_data_153 : _GEN_160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_162 = 8'h9a == _match_key_qbytes_0_T_2 ? phv_data_154 : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_163 = 8'h9b == _match_key_qbytes_0_T_2 ? phv_data_155 : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_164 = 8'h9c == _match_key_qbytes_0_T_2 ? phv_data_156 : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_165 = 8'h9d == _match_key_qbytes_0_T_2 ? phv_data_157 : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_166 = 8'h9e == _match_key_qbytes_0_T_2 ? phv_data_158 : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_167 = 8'h9f == _match_key_qbytes_0_T_2 ? phv_data_159 : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_168 = 8'ha0 == _match_key_qbytes_0_T_2 ? phv_data_160 : _GEN_167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_169 = 8'ha1 == _match_key_qbytes_0_T_2 ? phv_data_161 : _GEN_168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_170 = 8'ha2 == _match_key_qbytes_0_T_2 ? phv_data_162 : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_171 = 8'ha3 == _match_key_qbytes_0_T_2 ? phv_data_163 : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_172 = 8'ha4 == _match_key_qbytes_0_T_2 ? phv_data_164 : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_173 = 8'ha5 == _match_key_qbytes_0_T_2 ? phv_data_165 : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_174 = 8'ha6 == _match_key_qbytes_0_T_2 ? phv_data_166 : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_175 = 8'ha7 == _match_key_qbytes_0_T_2 ? phv_data_167 : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_176 = 8'ha8 == _match_key_qbytes_0_T_2 ? phv_data_168 : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_177 = 8'ha9 == _match_key_qbytes_0_T_2 ? phv_data_169 : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_178 = 8'haa == _match_key_qbytes_0_T_2 ? phv_data_170 : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_179 = 8'hab == _match_key_qbytes_0_T_2 ? phv_data_171 : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_180 = 8'hac == _match_key_qbytes_0_T_2 ? phv_data_172 : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_181 = 8'had == _match_key_qbytes_0_T_2 ? phv_data_173 : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_182 = 8'hae == _match_key_qbytes_0_T_2 ? phv_data_174 : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_183 = 8'haf == _match_key_qbytes_0_T_2 ? phv_data_175 : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_184 = 8'hb0 == _match_key_qbytes_0_T_2 ? phv_data_176 : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_185 = 8'hb1 == _match_key_qbytes_0_T_2 ? phv_data_177 : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_186 = 8'hb2 == _match_key_qbytes_0_T_2 ? phv_data_178 : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_187 = 8'hb3 == _match_key_qbytes_0_T_2 ? phv_data_179 : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_188 = 8'hb4 == _match_key_qbytes_0_T_2 ? phv_data_180 : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_189 = 8'hb5 == _match_key_qbytes_0_T_2 ? phv_data_181 : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_190 = 8'hb6 == _match_key_qbytes_0_T_2 ? phv_data_182 : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_191 = 8'hb7 == _match_key_qbytes_0_T_2 ? phv_data_183 : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_192 = 8'hb8 == _match_key_qbytes_0_T_2 ? phv_data_184 : _GEN_191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_193 = 8'hb9 == _match_key_qbytes_0_T_2 ? phv_data_185 : _GEN_192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_194 = 8'hba == _match_key_qbytes_0_T_2 ? phv_data_186 : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_195 = 8'hbb == _match_key_qbytes_0_T_2 ? phv_data_187 : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_196 = 8'hbc == _match_key_qbytes_0_T_2 ? phv_data_188 : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_197 = 8'hbd == _match_key_qbytes_0_T_2 ? phv_data_189 : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_198 = 8'hbe == _match_key_qbytes_0_T_2 ? phv_data_190 : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_199 = 8'hbf == _match_key_qbytes_0_T_2 ? phv_data_191 : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_200 = 8'hc0 == _match_key_qbytes_0_T_2 ? phv_data_192 : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_201 = 8'hc1 == _match_key_qbytes_0_T_2 ? phv_data_193 : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_202 = 8'hc2 == _match_key_qbytes_0_T_2 ? phv_data_194 : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_203 = 8'hc3 == _match_key_qbytes_0_T_2 ? phv_data_195 : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_204 = 8'hc4 == _match_key_qbytes_0_T_2 ? phv_data_196 : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_205 = 8'hc5 == _match_key_qbytes_0_T_2 ? phv_data_197 : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_206 = 8'hc6 == _match_key_qbytes_0_T_2 ? phv_data_198 : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_207 = 8'hc7 == _match_key_qbytes_0_T_2 ? phv_data_199 : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_208 = 8'hc8 == _match_key_qbytes_0_T_2 ? phv_data_200 : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_209 = 8'hc9 == _match_key_qbytes_0_T_2 ? phv_data_201 : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_210 = 8'hca == _match_key_qbytes_0_T_2 ? phv_data_202 : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_211 = 8'hcb == _match_key_qbytes_0_T_2 ? phv_data_203 : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_212 = 8'hcc == _match_key_qbytes_0_T_2 ? phv_data_204 : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_213 = 8'hcd == _match_key_qbytes_0_T_2 ? phv_data_205 : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_214 = 8'hce == _match_key_qbytes_0_T_2 ? phv_data_206 : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_215 = 8'hcf == _match_key_qbytes_0_T_2 ? phv_data_207 : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_216 = 8'hd0 == _match_key_qbytes_0_T_2 ? phv_data_208 : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_217 = 8'hd1 == _match_key_qbytes_0_T_2 ? phv_data_209 : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_218 = 8'hd2 == _match_key_qbytes_0_T_2 ? phv_data_210 : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_219 = 8'hd3 == _match_key_qbytes_0_T_2 ? phv_data_211 : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_220 = 8'hd4 == _match_key_qbytes_0_T_2 ? phv_data_212 : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_221 = 8'hd5 == _match_key_qbytes_0_T_2 ? phv_data_213 : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_222 = 8'hd6 == _match_key_qbytes_0_T_2 ? phv_data_214 : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_223 = 8'hd7 == _match_key_qbytes_0_T_2 ? phv_data_215 : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_224 = 8'hd8 == _match_key_qbytes_0_T_2 ? phv_data_216 : _GEN_223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_225 = 8'hd9 == _match_key_qbytes_0_T_2 ? phv_data_217 : _GEN_224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_226 = 8'hda == _match_key_qbytes_0_T_2 ? phv_data_218 : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_227 = 8'hdb == _match_key_qbytes_0_T_2 ? phv_data_219 : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_228 = 8'hdc == _match_key_qbytes_0_T_2 ? phv_data_220 : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_229 = 8'hdd == _match_key_qbytes_0_T_2 ? phv_data_221 : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_230 = 8'hde == _match_key_qbytes_0_T_2 ? phv_data_222 : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_231 = 8'hdf == _match_key_qbytes_0_T_2 ? phv_data_223 : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_232 = 8'he0 == _match_key_qbytes_0_T_2 ? phv_data_224 : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_233 = 8'he1 == _match_key_qbytes_0_T_2 ? phv_data_225 : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_234 = 8'he2 == _match_key_qbytes_0_T_2 ? phv_data_226 : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_235 = 8'he3 == _match_key_qbytes_0_T_2 ? phv_data_227 : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_236 = 8'he4 == _match_key_qbytes_0_T_2 ? phv_data_228 : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_237 = 8'he5 == _match_key_qbytes_0_T_2 ? phv_data_229 : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_238 = 8'he6 == _match_key_qbytes_0_T_2 ? phv_data_230 : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_239 = 8'he7 == _match_key_qbytes_0_T_2 ? phv_data_231 : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_240 = 8'he8 == _match_key_qbytes_0_T_2 ? phv_data_232 : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_241 = 8'he9 == _match_key_qbytes_0_T_2 ? phv_data_233 : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_242 = 8'hea == _match_key_qbytes_0_T_2 ? phv_data_234 : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_243 = 8'heb == _match_key_qbytes_0_T_2 ? phv_data_235 : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_244 = 8'hec == _match_key_qbytes_0_T_2 ? phv_data_236 : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_245 = 8'hed == _match_key_qbytes_0_T_2 ? phv_data_237 : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_246 = 8'hee == _match_key_qbytes_0_T_2 ? phv_data_238 : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_247 = 8'hef == _match_key_qbytes_0_T_2 ? phv_data_239 : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_248 = 8'hf0 == _match_key_qbytes_0_T_2 ? phv_data_240 : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_249 = 8'hf1 == _match_key_qbytes_0_T_2 ? phv_data_241 : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_250 = 8'hf2 == _match_key_qbytes_0_T_2 ? phv_data_242 : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_251 = 8'hf3 == _match_key_qbytes_0_T_2 ? phv_data_243 : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_252 = 8'hf4 == _match_key_qbytes_0_T_2 ? phv_data_244 : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_253 = 8'hf5 == _match_key_qbytes_0_T_2 ? phv_data_245 : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_254 = 8'hf6 == _match_key_qbytes_0_T_2 ? phv_data_246 : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_255 = 8'hf7 == _match_key_qbytes_0_T_2 ? phv_data_247 : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_256 = 8'hf8 == _match_key_qbytes_0_T_2 ? phv_data_248 : _GEN_255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_257 = 8'hf9 == _match_key_qbytes_0_T_2 ? phv_data_249 : _GEN_256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_258 = 8'hfa == _match_key_qbytes_0_T_2 ? phv_data_250 : _GEN_257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_259 = 8'hfb == _match_key_qbytes_0_T_2 ? phv_data_251 : _GEN_258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_260 = 8'hfc == _match_key_qbytes_0_T_2 ? phv_data_252 : _GEN_259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_261 = 8'hfd == _match_key_qbytes_0_T_2 ? phv_data_253 : _GEN_260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_262 = 8'hfe == _match_key_qbytes_0_T_2 ? phv_data_254 : _GEN_261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_263 = 8'hff == _match_key_qbytes_0_T_2 ? phv_data_255 : _GEN_262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_12326 = {{1'd0}, _match_key_qbytes_0_T_2}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_264 = 9'h100 == _GEN_12326 ? phv_data_256 : _GEN_263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_265 = 9'h101 == _GEN_12326 ? phv_data_257 : _GEN_264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_266 = 9'h102 == _GEN_12326 ? phv_data_258 : _GEN_265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_267 = 9'h103 == _GEN_12326 ? phv_data_259 : _GEN_266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_268 = 9'h104 == _GEN_12326 ? phv_data_260 : _GEN_267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_269 = 9'h105 == _GEN_12326 ? phv_data_261 : _GEN_268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_270 = 9'h106 == _GEN_12326 ? phv_data_262 : _GEN_269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_271 = 9'h107 == _GEN_12326 ? phv_data_263 : _GEN_270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_272 = 9'h108 == _GEN_12326 ? phv_data_264 : _GEN_271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_273 = 9'h109 == _GEN_12326 ? phv_data_265 : _GEN_272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_274 = 9'h10a == _GEN_12326 ? phv_data_266 : _GEN_273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_275 = 9'h10b == _GEN_12326 ? phv_data_267 : _GEN_274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_276 = 9'h10c == _GEN_12326 ? phv_data_268 : _GEN_275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_277 = 9'h10d == _GEN_12326 ? phv_data_269 : _GEN_276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_278 = 9'h10e == _GEN_12326 ? phv_data_270 : _GEN_277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_279 = 9'h10f == _GEN_12326 ? phv_data_271 : _GEN_278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_280 = 9'h110 == _GEN_12326 ? phv_data_272 : _GEN_279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_281 = 9'h111 == _GEN_12326 ? phv_data_273 : _GEN_280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_282 = 9'h112 == _GEN_12326 ? phv_data_274 : _GEN_281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_283 = 9'h113 == _GEN_12326 ? phv_data_275 : _GEN_282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_284 = 9'h114 == _GEN_12326 ? phv_data_276 : _GEN_283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_285 = 9'h115 == _GEN_12326 ? phv_data_277 : _GEN_284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_286 = 9'h116 == _GEN_12326 ? phv_data_278 : _GEN_285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_287 = 9'h117 == _GEN_12326 ? phv_data_279 : _GEN_286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_288 = 9'h118 == _GEN_12326 ? phv_data_280 : _GEN_287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_289 = 9'h119 == _GEN_12326 ? phv_data_281 : _GEN_288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_290 = 9'h11a == _GEN_12326 ? phv_data_282 : _GEN_289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_291 = 9'h11b == _GEN_12326 ? phv_data_283 : _GEN_290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_292 = 9'h11c == _GEN_12326 ? phv_data_284 : _GEN_291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_293 = 9'h11d == _GEN_12326 ? phv_data_285 : _GEN_292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_294 = 9'h11e == _GEN_12326 ? phv_data_286 : _GEN_293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_295 = 9'h11f == _GEN_12326 ? phv_data_287 : _GEN_294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_296 = 9'h120 == _GEN_12326 ? phv_data_288 : _GEN_295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_297 = 9'h121 == _GEN_12326 ? phv_data_289 : _GEN_296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_298 = 9'h122 == _GEN_12326 ? phv_data_290 : _GEN_297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_299 = 9'h123 == _GEN_12326 ? phv_data_291 : _GEN_298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_300 = 9'h124 == _GEN_12326 ? phv_data_292 : _GEN_299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_301 = 9'h125 == _GEN_12326 ? phv_data_293 : _GEN_300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_302 = 9'h126 == _GEN_12326 ? phv_data_294 : _GEN_301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_303 = 9'h127 == _GEN_12326 ? phv_data_295 : _GEN_302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_304 = 9'h128 == _GEN_12326 ? phv_data_296 : _GEN_303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_305 = 9'h129 == _GEN_12326 ? phv_data_297 : _GEN_304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_306 = 9'h12a == _GEN_12326 ? phv_data_298 : _GEN_305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_307 = 9'h12b == _GEN_12326 ? phv_data_299 : _GEN_306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_308 = 9'h12c == _GEN_12326 ? phv_data_300 : _GEN_307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_309 = 9'h12d == _GEN_12326 ? phv_data_301 : _GEN_308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_310 = 9'h12e == _GEN_12326 ? phv_data_302 : _GEN_309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_311 = 9'h12f == _GEN_12326 ? phv_data_303 : _GEN_310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_312 = 9'h130 == _GEN_12326 ? phv_data_304 : _GEN_311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_313 = 9'h131 == _GEN_12326 ? phv_data_305 : _GEN_312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_314 = 9'h132 == _GEN_12326 ? phv_data_306 : _GEN_313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_315 = 9'h133 == _GEN_12326 ? phv_data_307 : _GEN_314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_316 = 9'h134 == _GEN_12326 ? phv_data_308 : _GEN_315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_317 = 9'h135 == _GEN_12326 ? phv_data_309 : _GEN_316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_318 = 9'h136 == _GEN_12326 ? phv_data_310 : _GEN_317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_319 = 9'h137 == _GEN_12326 ? phv_data_311 : _GEN_318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_320 = 9'h138 == _GEN_12326 ? phv_data_312 : _GEN_319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_321 = 9'h139 == _GEN_12326 ? phv_data_313 : _GEN_320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_322 = 9'h13a == _GEN_12326 ? phv_data_314 : _GEN_321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_323 = 9'h13b == _GEN_12326 ? phv_data_315 : _GEN_322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_324 = 9'h13c == _GEN_12326 ? phv_data_316 : _GEN_323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_325 = 9'h13d == _GEN_12326 ? phv_data_317 : _GEN_324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_326 = 9'h13e == _GEN_12326 ? phv_data_318 : _GEN_325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_327 = 9'h13f == _GEN_12326 ? phv_data_319 : _GEN_326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_328 = 9'h140 == _GEN_12326 ? phv_data_320 : _GEN_327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_329 = 9'h141 == _GEN_12326 ? phv_data_321 : _GEN_328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_330 = 9'h142 == _GEN_12326 ? phv_data_322 : _GEN_329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_331 = 9'h143 == _GEN_12326 ? phv_data_323 : _GEN_330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_332 = 9'h144 == _GEN_12326 ? phv_data_324 : _GEN_331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_333 = 9'h145 == _GEN_12326 ? phv_data_325 : _GEN_332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_334 = 9'h146 == _GEN_12326 ? phv_data_326 : _GEN_333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_335 = 9'h147 == _GEN_12326 ? phv_data_327 : _GEN_334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_336 = 9'h148 == _GEN_12326 ? phv_data_328 : _GEN_335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_337 = 9'h149 == _GEN_12326 ? phv_data_329 : _GEN_336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_338 = 9'h14a == _GEN_12326 ? phv_data_330 : _GEN_337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_339 = 9'h14b == _GEN_12326 ? phv_data_331 : _GEN_338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_340 = 9'h14c == _GEN_12326 ? phv_data_332 : _GEN_339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_341 = 9'h14d == _GEN_12326 ? phv_data_333 : _GEN_340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_342 = 9'h14e == _GEN_12326 ? phv_data_334 : _GEN_341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_343 = 9'h14f == _GEN_12326 ? phv_data_335 : _GEN_342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_344 = 9'h150 == _GEN_12326 ? phv_data_336 : _GEN_343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_345 = 9'h151 == _GEN_12326 ? phv_data_337 : _GEN_344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_346 = 9'h152 == _GEN_12326 ? phv_data_338 : _GEN_345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_347 = 9'h153 == _GEN_12326 ? phv_data_339 : _GEN_346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_348 = 9'h154 == _GEN_12326 ? phv_data_340 : _GEN_347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_349 = 9'h155 == _GEN_12326 ? phv_data_341 : _GEN_348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_350 = 9'h156 == _GEN_12326 ? phv_data_342 : _GEN_349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_351 = 9'h157 == _GEN_12326 ? phv_data_343 : _GEN_350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_352 = 9'h158 == _GEN_12326 ? phv_data_344 : _GEN_351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_353 = 9'h159 == _GEN_12326 ? phv_data_345 : _GEN_352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_354 = 9'h15a == _GEN_12326 ? phv_data_346 : _GEN_353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_355 = 9'h15b == _GEN_12326 ? phv_data_347 : _GEN_354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_356 = 9'h15c == _GEN_12326 ? phv_data_348 : _GEN_355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_357 = 9'h15d == _GEN_12326 ? phv_data_349 : _GEN_356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_358 = 9'h15e == _GEN_12326 ? phv_data_350 : _GEN_357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_359 = 9'h15f == _GEN_12326 ? phv_data_351 : _GEN_358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_360 = 9'h160 == _GEN_12326 ? phv_data_352 : _GEN_359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_361 = 9'h161 == _GEN_12326 ? phv_data_353 : _GEN_360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_362 = 9'h162 == _GEN_12326 ? phv_data_354 : _GEN_361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_363 = 9'h163 == _GEN_12326 ? phv_data_355 : _GEN_362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_364 = 9'h164 == _GEN_12326 ? phv_data_356 : _GEN_363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_365 = 9'h165 == _GEN_12326 ? phv_data_357 : _GEN_364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_366 = 9'h166 == _GEN_12326 ? phv_data_358 : _GEN_365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_367 = 9'h167 == _GEN_12326 ? phv_data_359 : _GEN_366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_368 = 9'h168 == _GEN_12326 ? phv_data_360 : _GEN_367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_369 = 9'h169 == _GEN_12326 ? phv_data_361 : _GEN_368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_370 = 9'h16a == _GEN_12326 ? phv_data_362 : _GEN_369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_371 = 9'h16b == _GEN_12326 ? phv_data_363 : _GEN_370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_372 = 9'h16c == _GEN_12326 ? phv_data_364 : _GEN_371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_373 = 9'h16d == _GEN_12326 ? phv_data_365 : _GEN_372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_374 = 9'h16e == _GEN_12326 ? phv_data_366 : _GEN_373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_375 = 9'h16f == _GEN_12326 ? phv_data_367 : _GEN_374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_376 = 9'h170 == _GEN_12326 ? phv_data_368 : _GEN_375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_377 = 9'h171 == _GEN_12326 ? phv_data_369 : _GEN_376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_378 = 9'h172 == _GEN_12326 ? phv_data_370 : _GEN_377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_379 = 9'h173 == _GEN_12326 ? phv_data_371 : _GEN_378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_380 = 9'h174 == _GEN_12326 ? phv_data_372 : _GEN_379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_381 = 9'h175 == _GEN_12326 ? phv_data_373 : _GEN_380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_382 = 9'h176 == _GEN_12326 ? phv_data_374 : _GEN_381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_383 = 9'h177 == _GEN_12326 ? phv_data_375 : _GEN_382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_384 = 9'h178 == _GEN_12326 ? phv_data_376 : _GEN_383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_385 = 9'h179 == _GEN_12326 ? phv_data_377 : _GEN_384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_386 = 9'h17a == _GEN_12326 ? phv_data_378 : _GEN_385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_387 = 9'h17b == _GEN_12326 ? phv_data_379 : _GEN_386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_388 = 9'h17c == _GEN_12326 ? phv_data_380 : _GEN_387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_389 = 9'h17d == _GEN_12326 ? phv_data_381 : _GEN_388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_390 = 9'h17e == _GEN_12326 ? phv_data_382 : _GEN_389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_391 = 9'h17f == _GEN_12326 ? phv_data_383 : _GEN_390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_392 = 9'h180 == _GEN_12326 ? phv_data_384 : _GEN_391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_393 = 9'h181 == _GEN_12326 ? phv_data_385 : _GEN_392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_394 = 9'h182 == _GEN_12326 ? phv_data_386 : _GEN_393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_395 = 9'h183 == _GEN_12326 ? phv_data_387 : _GEN_394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_396 = 9'h184 == _GEN_12326 ? phv_data_388 : _GEN_395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_397 = 9'h185 == _GEN_12326 ? phv_data_389 : _GEN_396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_398 = 9'h186 == _GEN_12326 ? phv_data_390 : _GEN_397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_399 = 9'h187 == _GEN_12326 ? phv_data_391 : _GEN_398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_400 = 9'h188 == _GEN_12326 ? phv_data_392 : _GEN_399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_401 = 9'h189 == _GEN_12326 ? phv_data_393 : _GEN_400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_402 = 9'h18a == _GEN_12326 ? phv_data_394 : _GEN_401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_403 = 9'h18b == _GEN_12326 ? phv_data_395 : _GEN_402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_404 = 9'h18c == _GEN_12326 ? phv_data_396 : _GEN_403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_405 = 9'h18d == _GEN_12326 ? phv_data_397 : _GEN_404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_406 = 9'h18e == _GEN_12326 ? phv_data_398 : _GEN_405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_407 = 9'h18f == _GEN_12326 ? phv_data_399 : _GEN_406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_408 = 9'h190 == _GEN_12326 ? phv_data_400 : _GEN_407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_409 = 9'h191 == _GEN_12326 ? phv_data_401 : _GEN_408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_410 = 9'h192 == _GEN_12326 ? phv_data_402 : _GEN_409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_411 = 9'h193 == _GEN_12326 ? phv_data_403 : _GEN_410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_412 = 9'h194 == _GEN_12326 ? phv_data_404 : _GEN_411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_413 = 9'h195 == _GEN_12326 ? phv_data_405 : _GEN_412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_414 = 9'h196 == _GEN_12326 ? phv_data_406 : _GEN_413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_415 = 9'h197 == _GEN_12326 ? phv_data_407 : _GEN_414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_416 = 9'h198 == _GEN_12326 ? phv_data_408 : _GEN_415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_417 = 9'h199 == _GEN_12326 ? phv_data_409 : _GEN_416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_418 = 9'h19a == _GEN_12326 ? phv_data_410 : _GEN_417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_419 = 9'h19b == _GEN_12326 ? phv_data_411 : _GEN_418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_420 = 9'h19c == _GEN_12326 ? phv_data_412 : _GEN_419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_421 = 9'h19d == _GEN_12326 ? phv_data_413 : _GEN_420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_422 = 9'h19e == _GEN_12326 ? phv_data_414 : _GEN_421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_423 = 9'h19f == _GEN_12326 ? phv_data_415 : _GEN_422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_424 = 9'h1a0 == _GEN_12326 ? phv_data_416 : _GEN_423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_425 = 9'h1a1 == _GEN_12326 ? phv_data_417 : _GEN_424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_426 = 9'h1a2 == _GEN_12326 ? phv_data_418 : _GEN_425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_427 = 9'h1a3 == _GEN_12326 ? phv_data_419 : _GEN_426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_428 = 9'h1a4 == _GEN_12326 ? phv_data_420 : _GEN_427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_429 = 9'h1a5 == _GEN_12326 ? phv_data_421 : _GEN_428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_430 = 9'h1a6 == _GEN_12326 ? phv_data_422 : _GEN_429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_431 = 9'h1a7 == _GEN_12326 ? phv_data_423 : _GEN_430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_432 = 9'h1a8 == _GEN_12326 ? phv_data_424 : _GEN_431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_433 = 9'h1a9 == _GEN_12326 ? phv_data_425 : _GEN_432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_434 = 9'h1aa == _GEN_12326 ? phv_data_426 : _GEN_433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_435 = 9'h1ab == _GEN_12326 ? phv_data_427 : _GEN_434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_436 = 9'h1ac == _GEN_12326 ? phv_data_428 : _GEN_435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_437 = 9'h1ad == _GEN_12326 ? phv_data_429 : _GEN_436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_438 = 9'h1ae == _GEN_12326 ? phv_data_430 : _GEN_437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_439 = 9'h1af == _GEN_12326 ? phv_data_431 : _GEN_438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_440 = 9'h1b0 == _GEN_12326 ? phv_data_432 : _GEN_439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_441 = 9'h1b1 == _GEN_12326 ? phv_data_433 : _GEN_440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_442 = 9'h1b2 == _GEN_12326 ? phv_data_434 : _GEN_441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_443 = 9'h1b3 == _GEN_12326 ? phv_data_435 : _GEN_442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_444 = 9'h1b4 == _GEN_12326 ? phv_data_436 : _GEN_443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_445 = 9'h1b5 == _GEN_12326 ? phv_data_437 : _GEN_444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_446 = 9'h1b6 == _GEN_12326 ? phv_data_438 : _GEN_445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_447 = 9'h1b7 == _GEN_12326 ? phv_data_439 : _GEN_446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_448 = 9'h1b8 == _GEN_12326 ? phv_data_440 : _GEN_447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_449 = 9'h1b9 == _GEN_12326 ? phv_data_441 : _GEN_448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_450 = 9'h1ba == _GEN_12326 ? phv_data_442 : _GEN_449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_451 = 9'h1bb == _GEN_12326 ? phv_data_443 : _GEN_450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_452 = 9'h1bc == _GEN_12326 ? phv_data_444 : _GEN_451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_453 = 9'h1bd == _GEN_12326 ? phv_data_445 : _GEN_452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_454 = 9'h1be == _GEN_12326 ? phv_data_446 : _GEN_453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_455 = 9'h1bf == _GEN_12326 ? phv_data_447 : _GEN_454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_456 = 9'h1c0 == _GEN_12326 ? phv_data_448 : _GEN_455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_457 = 9'h1c1 == _GEN_12326 ? phv_data_449 : _GEN_456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_458 = 9'h1c2 == _GEN_12326 ? phv_data_450 : _GEN_457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_459 = 9'h1c3 == _GEN_12326 ? phv_data_451 : _GEN_458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_460 = 9'h1c4 == _GEN_12326 ? phv_data_452 : _GEN_459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_461 = 9'h1c5 == _GEN_12326 ? phv_data_453 : _GEN_460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_462 = 9'h1c6 == _GEN_12326 ? phv_data_454 : _GEN_461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_463 = 9'h1c7 == _GEN_12326 ? phv_data_455 : _GEN_462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_464 = 9'h1c8 == _GEN_12326 ? phv_data_456 : _GEN_463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_465 = 9'h1c9 == _GEN_12326 ? phv_data_457 : _GEN_464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_466 = 9'h1ca == _GEN_12326 ? phv_data_458 : _GEN_465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_467 = 9'h1cb == _GEN_12326 ? phv_data_459 : _GEN_466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_468 = 9'h1cc == _GEN_12326 ? phv_data_460 : _GEN_467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_469 = 9'h1cd == _GEN_12326 ? phv_data_461 : _GEN_468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_470 = 9'h1ce == _GEN_12326 ? phv_data_462 : _GEN_469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_471 = 9'h1cf == _GEN_12326 ? phv_data_463 : _GEN_470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_472 = 9'h1d0 == _GEN_12326 ? phv_data_464 : _GEN_471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_473 = 9'h1d1 == _GEN_12326 ? phv_data_465 : _GEN_472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_474 = 9'h1d2 == _GEN_12326 ? phv_data_466 : _GEN_473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_475 = 9'h1d3 == _GEN_12326 ? phv_data_467 : _GEN_474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_476 = 9'h1d4 == _GEN_12326 ? phv_data_468 : _GEN_475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_477 = 9'h1d5 == _GEN_12326 ? phv_data_469 : _GEN_476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_478 = 9'h1d6 == _GEN_12326 ? phv_data_470 : _GEN_477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_479 = 9'h1d7 == _GEN_12326 ? phv_data_471 : _GEN_478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_480 = 9'h1d8 == _GEN_12326 ? phv_data_472 : _GEN_479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_481 = 9'h1d9 == _GEN_12326 ? phv_data_473 : _GEN_480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_482 = 9'h1da == _GEN_12326 ? phv_data_474 : _GEN_481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_483 = 9'h1db == _GEN_12326 ? phv_data_475 : _GEN_482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_484 = 9'h1dc == _GEN_12326 ? phv_data_476 : _GEN_483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_485 = 9'h1dd == _GEN_12326 ? phv_data_477 : _GEN_484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_486 = 9'h1de == _GEN_12326 ? phv_data_478 : _GEN_485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_487 = 9'h1df == _GEN_12326 ? phv_data_479 : _GEN_486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_488 = 9'h1e0 == _GEN_12326 ? phv_data_480 : _GEN_487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_489 = 9'h1e1 == _GEN_12326 ? phv_data_481 : _GEN_488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_490 = 9'h1e2 == _GEN_12326 ? phv_data_482 : _GEN_489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_491 = 9'h1e3 == _GEN_12326 ? phv_data_483 : _GEN_490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_492 = 9'h1e4 == _GEN_12326 ? phv_data_484 : _GEN_491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_493 = 9'h1e5 == _GEN_12326 ? phv_data_485 : _GEN_492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_494 = 9'h1e6 == _GEN_12326 ? phv_data_486 : _GEN_493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_495 = 9'h1e7 == _GEN_12326 ? phv_data_487 : _GEN_494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_496 = 9'h1e8 == _GEN_12326 ? phv_data_488 : _GEN_495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_497 = 9'h1e9 == _GEN_12326 ? phv_data_489 : _GEN_496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_498 = 9'h1ea == _GEN_12326 ? phv_data_490 : _GEN_497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_499 = 9'h1eb == _GEN_12326 ? phv_data_491 : _GEN_498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_500 = 9'h1ec == _GEN_12326 ? phv_data_492 : _GEN_499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_501 = 9'h1ed == _GEN_12326 ? phv_data_493 : _GEN_500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_502 = 9'h1ee == _GEN_12326 ? phv_data_494 : _GEN_501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_503 = 9'h1ef == _GEN_12326 ? phv_data_495 : _GEN_502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_504 = 9'h1f0 == _GEN_12326 ? phv_data_496 : _GEN_503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_505 = 9'h1f1 == _GEN_12326 ? phv_data_497 : _GEN_504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_506 = 9'h1f2 == _GEN_12326 ? phv_data_498 : _GEN_505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_507 = 9'h1f3 == _GEN_12326 ? phv_data_499 : _GEN_506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_508 = 9'h1f4 == _GEN_12326 ? phv_data_500 : _GEN_507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_509 = 9'h1f5 == _GEN_12326 ? phv_data_501 : _GEN_508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_510 = 9'h1f6 == _GEN_12326 ? phv_data_502 : _GEN_509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_511 = 9'h1f7 == _GEN_12326 ? phv_data_503 : _GEN_510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_512 = 9'h1f8 == _GEN_12326 ? phv_data_504 : _GEN_511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_513 = 9'h1f9 == _GEN_12326 ? phv_data_505 : _GEN_512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_514 = 9'h1fa == _GEN_12326 ? phv_data_506 : _GEN_513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_515 = 9'h1fb == _GEN_12326 ? phv_data_507 : _GEN_514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_516 = 9'h1fc == _GEN_12326 ? phv_data_508 : _GEN_515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_517 = 9'h1fd == _GEN_12326 ? phv_data_509 : _GEN_516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_518 = 9'h1fe == _GEN_12326 ? phv_data_510 : _GEN_517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_519 = 9'h1ff == _GEN_12326 ? phv_data_511 : _GEN_518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_521 = 8'h1 == local_offset ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_522 = 8'h2 == local_offset ? phv_data_2 : _GEN_521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_523 = 8'h3 == local_offset ? phv_data_3 : _GEN_522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_524 = 8'h4 == local_offset ? phv_data_4 : _GEN_523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_525 = 8'h5 == local_offset ? phv_data_5 : _GEN_524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_526 = 8'h6 == local_offset ? phv_data_6 : _GEN_525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_527 = 8'h7 == local_offset ? phv_data_7 : _GEN_526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_528 = 8'h8 == local_offset ? phv_data_8 : _GEN_527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_529 = 8'h9 == local_offset ? phv_data_9 : _GEN_528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_530 = 8'ha == local_offset ? phv_data_10 : _GEN_529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_531 = 8'hb == local_offset ? phv_data_11 : _GEN_530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_532 = 8'hc == local_offset ? phv_data_12 : _GEN_531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_533 = 8'hd == local_offset ? phv_data_13 : _GEN_532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_534 = 8'he == local_offset ? phv_data_14 : _GEN_533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_535 = 8'hf == local_offset ? phv_data_15 : _GEN_534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_536 = 8'h10 == local_offset ? phv_data_16 : _GEN_535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_537 = 8'h11 == local_offset ? phv_data_17 : _GEN_536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_538 = 8'h12 == local_offset ? phv_data_18 : _GEN_537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_539 = 8'h13 == local_offset ? phv_data_19 : _GEN_538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_540 = 8'h14 == local_offset ? phv_data_20 : _GEN_539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_541 = 8'h15 == local_offset ? phv_data_21 : _GEN_540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_542 = 8'h16 == local_offset ? phv_data_22 : _GEN_541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_543 = 8'h17 == local_offset ? phv_data_23 : _GEN_542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_544 = 8'h18 == local_offset ? phv_data_24 : _GEN_543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_545 = 8'h19 == local_offset ? phv_data_25 : _GEN_544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_546 = 8'h1a == local_offset ? phv_data_26 : _GEN_545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_547 = 8'h1b == local_offset ? phv_data_27 : _GEN_546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_548 = 8'h1c == local_offset ? phv_data_28 : _GEN_547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_549 = 8'h1d == local_offset ? phv_data_29 : _GEN_548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_550 = 8'h1e == local_offset ? phv_data_30 : _GEN_549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_551 = 8'h1f == local_offset ? phv_data_31 : _GEN_550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_552 = 8'h20 == local_offset ? phv_data_32 : _GEN_551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_553 = 8'h21 == local_offset ? phv_data_33 : _GEN_552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_554 = 8'h22 == local_offset ? phv_data_34 : _GEN_553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_555 = 8'h23 == local_offset ? phv_data_35 : _GEN_554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_556 = 8'h24 == local_offset ? phv_data_36 : _GEN_555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_557 = 8'h25 == local_offset ? phv_data_37 : _GEN_556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_558 = 8'h26 == local_offset ? phv_data_38 : _GEN_557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_559 = 8'h27 == local_offset ? phv_data_39 : _GEN_558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_560 = 8'h28 == local_offset ? phv_data_40 : _GEN_559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_561 = 8'h29 == local_offset ? phv_data_41 : _GEN_560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_562 = 8'h2a == local_offset ? phv_data_42 : _GEN_561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_563 = 8'h2b == local_offset ? phv_data_43 : _GEN_562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_564 = 8'h2c == local_offset ? phv_data_44 : _GEN_563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_565 = 8'h2d == local_offset ? phv_data_45 : _GEN_564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_566 = 8'h2e == local_offset ? phv_data_46 : _GEN_565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_567 = 8'h2f == local_offset ? phv_data_47 : _GEN_566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_568 = 8'h30 == local_offset ? phv_data_48 : _GEN_567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_569 = 8'h31 == local_offset ? phv_data_49 : _GEN_568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_570 = 8'h32 == local_offset ? phv_data_50 : _GEN_569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_571 = 8'h33 == local_offset ? phv_data_51 : _GEN_570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_572 = 8'h34 == local_offset ? phv_data_52 : _GEN_571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_573 = 8'h35 == local_offset ? phv_data_53 : _GEN_572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_574 = 8'h36 == local_offset ? phv_data_54 : _GEN_573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_575 = 8'h37 == local_offset ? phv_data_55 : _GEN_574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_576 = 8'h38 == local_offset ? phv_data_56 : _GEN_575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_577 = 8'h39 == local_offset ? phv_data_57 : _GEN_576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_578 = 8'h3a == local_offset ? phv_data_58 : _GEN_577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_579 = 8'h3b == local_offset ? phv_data_59 : _GEN_578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_580 = 8'h3c == local_offset ? phv_data_60 : _GEN_579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_581 = 8'h3d == local_offset ? phv_data_61 : _GEN_580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_582 = 8'h3e == local_offset ? phv_data_62 : _GEN_581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_583 = 8'h3f == local_offset ? phv_data_63 : _GEN_582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_584 = 8'h40 == local_offset ? phv_data_64 : _GEN_583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_585 = 8'h41 == local_offset ? phv_data_65 : _GEN_584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_586 = 8'h42 == local_offset ? phv_data_66 : _GEN_585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_587 = 8'h43 == local_offset ? phv_data_67 : _GEN_586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_588 = 8'h44 == local_offset ? phv_data_68 : _GEN_587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_589 = 8'h45 == local_offset ? phv_data_69 : _GEN_588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_590 = 8'h46 == local_offset ? phv_data_70 : _GEN_589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_591 = 8'h47 == local_offset ? phv_data_71 : _GEN_590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_592 = 8'h48 == local_offset ? phv_data_72 : _GEN_591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_593 = 8'h49 == local_offset ? phv_data_73 : _GEN_592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_594 = 8'h4a == local_offset ? phv_data_74 : _GEN_593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_595 = 8'h4b == local_offset ? phv_data_75 : _GEN_594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_596 = 8'h4c == local_offset ? phv_data_76 : _GEN_595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_597 = 8'h4d == local_offset ? phv_data_77 : _GEN_596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_598 = 8'h4e == local_offset ? phv_data_78 : _GEN_597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_599 = 8'h4f == local_offset ? phv_data_79 : _GEN_598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_600 = 8'h50 == local_offset ? phv_data_80 : _GEN_599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_601 = 8'h51 == local_offset ? phv_data_81 : _GEN_600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_602 = 8'h52 == local_offset ? phv_data_82 : _GEN_601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_603 = 8'h53 == local_offset ? phv_data_83 : _GEN_602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_604 = 8'h54 == local_offset ? phv_data_84 : _GEN_603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_605 = 8'h55 == local_offset ? phv_data_85 : _GEN_604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_606 = 8'h56 == local_offset ? phv_data_86 : _GEN_605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_607 = 8'h57 == local_offset ? phv_data_87 : _GEN_606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_608 = 8'h58 == local_offset ? phv_data_88 : _GEN_607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_609 = 8'h59 == local_offset ? phv_data_89 : _GEN_608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_610 = 8'h5a == local_offset ? phv_data_90 : _GEN_609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_611 = 8'h5b == local_offset ? phv_data_91 : _GEN_610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_612 = 8'h5c == local_offset ? phv_data_92 : _GEN_611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_613 = 8'h5d == local_offset ? phv_data_93 : _GEN_612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_614 = 8'h5e == local_offset ? phv_data_94 : _GEN_613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_615 = 8'h5f == local_offset ? phv_data_95 : _GEN_614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_616 = 8'h60 == local_offset ? phv_data_96 : _GEN_615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_617 = 8'h61 == local_offset ? phv_data_97 : _GEN_616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_618 = 8'h62 == local_offset ? phv_data_98 : _GEN_617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_619 = 8'h63 == local_offset ? phv_data_99 : _GEN_618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_620 = 8'h64 == local_offset ? phv_data_100 : _GEN_619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_621 = 8'h65 == local_offset ? phv_data_101 : _GEN_620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_622 = 8'h66 == local_offset ? phv_data_102 : _GEN_621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_623 = 8'h67 == local_offset ? phv_data_103 : _GEN_622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_624 = 8'h68 == local_offset ? phv_data_104 : _GEN_623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_625 = 8'h69 == local_offset ? phv_data_105 : _GEN_624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_626 = 8'h6a == local_offset ? phv_data_106 : _GEN_625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_627 = 8'h6b == local_offset ? phv_data_107 : _GEN_626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_628 = 8'h6c == local_offset ? phv_data_108 : _GEN_627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_629 = 8'h6d == local_offset ? phv_data_109 : _GEN_628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_630 = 8'h6e == local_offset ? phv_data_110 : _GEN_629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_631 = 8'h6f == local_offset ? phv_data_111 : _GEN_630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_632 = 8'h70 == local_offset ? phv_data_112 : _GEN_631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_633 = 8'h71 == local_offset ? phv_data_113 : _GEN_632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_634 = 8'h72 == local_offset ? phv_data_114 : _GEN_633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_635 = 8'h73 == local_offset ? phv_data_115 : _GEN_634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_636 = 8'h74 == local_offset ? phv_data_116 : _GEN_635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_637 = 8'h75 == local_offset ? phv_data_117 : _GEN_636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_638 = 8'h76 == local_offset ? phv_data_118 : _GEN_637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_639 = 8'h77 == local_offset ? phv_data_119 : _GEN_638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_640 = 8'h78 == local_offset ? phv_data_120 : _GEN_639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_641 = 8'h79 == local_offset ? phv_data_121 : _GEN_640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_642 = 8'h7a == local_offset ? phv_data_122 : _GEN_641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_643 = 8'h7b == local_offset ? phv_data_123 : _GEN_642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_644 = 8'h7c == local_offset ? phv_data_124 : _GEN_643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_645 = 8'h7d == local_offset ? phv_data_125 : _GEN_644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_646 = 8'h7e == local_offset ? phv_data_126 : _GEN_645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_647 = 8'h7f == local_offset ? phv_data_127 : _GEN_646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_648 = 8'h80 == local_offset ? phv_data_128 : _GEN_647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_649 = 8'h81 == local_offset ? phv_data_129 : _GEN_648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_650 = 8'h82 == local_offset ? phv_data_130 : _GEN_649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_651 = 8'h83 == local_offset ? phv_data_131 : _GEN_650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_652 = 8'h84 == local_offset ? phv_data_132 : _GEN_651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_653 = 8'h85 == local_offset ? phv_data_133 : _GEN_652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_654 = 8'h86 == local_offset ? phv_data_134 : _GEN_653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_655 = 8'h87 == local_offset ? phv_data_135 : _GEN_654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_656 = 8'h88 == local_offset ? phv_data_136 : _GEN_655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_657 = 8'h89 == local_offset ? phv_data_137 : _GEN_656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_658 = 8'h8a == local_offset ? phv_data_138 : _GEN_657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_659 = 8'h8b == local_offset ? phv_data_139 : _GEN_658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_660 = 8'h8c == local_offset ? phv_data_140 : _GEN_659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_661 = 8'h8d == local_offset ? phv_data_141 : _GEN_660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_662 = 8'h8e == local_offset ? phv_data_142 : _GEN_661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_663 = 8'h8f == local_offset ? phv_data_143 : _GEN_662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_664 = 8'h90 == local_offset ? phv_data_144 : _GEN_663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_665 = 8'h91 == local_offset ? phv_data_145 : _GEN_664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_666 = 8'h92 == local_offset ? phv_data_146 : _GEN_665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_667 = 8'h93 == local_offset ? phv_data_147 : _GEN_666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_668 = 8'h94 == local_offset ? phv_data_148 : _GEN_667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_669 = 8'h95 == local_offset ? phv_data_149 : _GEN_668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_670 = 8'h96 == local_offset ? phv_data_150 : _GEN_669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_671 = 8'h97 == local_offset ? phv_data_151 : _GEN_670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_672 = 8'h98 == local_offset ? phv_data_152 : _GEN_671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_673 = 8'h99 == local_offset ? phv_data_153 : _GEN_672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_674 = 8'h9a == local_offset ? phv_data_154 : _GEN_673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_675 = 8'h9b == local_offset ? phv_data_155 : _GEN_674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_676 = 8'h9c == local_offset ? phv_data_156 : _GEN_675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_677 = 8'h9d == local_offset ? phv_data_157 : _GEN_676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_678 = 8'h9e == local_offset ? phv_data_158 : _GEN_677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_679 = 8'h9f == local_offset ? phv_data_159 : _GEN_678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_680 = 8'ha0 == local_offset ? phv_data_160 : _GEN_679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_681 = 8'ha1 == local_offset ? phv_data_161 : _GEN_680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_682 = 8'ha2 == local_offset ? phv_data_162 : _GEN_681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_683 = 8'ha3 == local_offset ? phv_data_163 : _GEN_682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_684 = 8'ha4 == local_offset ? phv_data_164 : _GEN_683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_685 = 8'ha5 == local_offset ? phv_data_165 : _GEN_684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_686 = 8'ha6 == local_offset ? phv_data_166 : _GEN_685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_687 = 8'ha7 == local_offset ? phv_data_167 : _GEN_686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_688 = 8'ha8 == local_offset ? phv_data_168 : _GEN_687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_689 = 8'ha9 == local_offset ? phv_data_169 : _GEN_688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_690 = 8'haa == local_offset ? phv_data_170 : _GEN_689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_691 = 8'hab == local_offset ? phv_data_171 : _GEN_690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_692 = 8'hac == local_offset ? phv_data_172 : _GEN_691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_693 = 8'had == local_offset ? phv_data_173 : _GEN_692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_694 = 8'hae == local_offset ? phv_data_174 : _GEN_693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_695 = 8'haf == local_offset ? phv_data_175 : _GEN_694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_696 = 8'hb0 == local_offset ? phv_data_176 : _GEN_695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_697 = 8'hb1 == local_offset ? phv_data_177 : _GEN_696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_698 = 8'hb2 == local_offset ? phv_data_178 : _GEN_697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_699 = 8'hb3 == local_offset ? phv_data_179 : _GEN_698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_700 = 8'hb4 == local_offset ? phv_data_180 : _GEN_699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_701 = 8'hb5 == local_offset ? phv_data_181 : _GEN_700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_702 = 8'hb6 == local_offset ? phv_data_182 : _GEN_701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_703 = 8'hb7 == local_offset ? phv_data_183 : _GEN_702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_704 = 8'hb8 == local_offset ? phv_data_184 : _GEN_703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_705 = 8'hb9 == local_offset ? phv_data_185 : _GEN_704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_706 = 8'hba == local_offset ? phv_data_186 : _GEN_705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_707 = 8'hbb == local_offset ? phv_data_187 : _GEN_706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_708 = 8'hbc == local_offset ? phv_data_188 : _GEN_707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_709 = 8'hbd == local_offset ? phv_data_189 : _GEN_708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_710 = 8'hbe == local_offset ? phv_data_190 : _GEN_709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_711 = 8'hbf == local_offset ? phv_data_191 : _GEN_710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_712 = 8'hc0 == local_offset ? phv_data_192 : _GEN_711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_713 = 8'hc1 == local_offset ? phv_data_193 : _GEN_712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_714 = 8'hc2 == local_offset ? phv_data_194 : _GEN_713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_715 = 8'hc3 == local_offset ? phv_data_195 : _GEN_714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_716 = 8'hc4 == local_offset ? phv_data_196 : _GEN_715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_717 = 8'hc5 == local_offset ? phv_data_197 : _GEN_716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_718 = 8'hc6 == local_offset ? phv_data_198 : _GEN_717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_719 = 8'hc7 == local_offset ? phv_data_199 : _GEN_718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_720 = 8'hc8 == local_offset ? phv_data_200 : _GEN_719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_721 = 8'hc9 == local_offset ? phv_data_201 : _GEN_720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_722 = 8'hca == local_offset ? phv_data_202 : _GEN_721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_723 = 8'hcb == local_offset ? phv_data_203 : _GEN_722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_724 = 8'hcc == local_offset ? phv_data_204 : _GEN_723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_725 = 8'hcd == local_offset ? phv_data_205 : _GEN_724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_726 = 8'hce == local_offset ? phv_data_206 : _GEN_725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_727 = 8'hcf == local_offset ? phv_data_207 : _GEN_726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_728 = 8'hd0 == local_offset ? phv_data_208 : _GEN_727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_729 = 8'hd1 == local_offset ? phv_data_209 : _GEN_728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_730 = 8'hd2 == local_offset ? phv_data_210 : _GEN_729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_731 = 8'hd3 == local_offset ? phv_data_211 : _GEN_730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_732 = 8'hd4 == local_offset ? phv_data_212 : _GEN_731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_733 = 8'hd5 == local_offset ? phv_data_213 : _GEN_732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_734 = 8'hd6 == local_offset ? phv_data_214 : _GEN_733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_735 = 8'hd7 == local_offset ? phv_data_215 : _GEN_734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_736 = 8'hd8 == local_offset ? phv_data_216 : _GEN_735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_737 = 8'hd9 == local_offset ? phv_data_217 : _GEN_736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_738 = 8'hda == local_offset ? phv_data_218 : _GEN_737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_739 = 8'hdb == local_offset ? phv_data_219 : _GEN_738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_740 = 8'hdc == local_offset ? phv_data_220 : _GEN_739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_741 = 8'hdd == local_offset ? phv_data_221 : _GEN_740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_742 = 8'hde == local_offset ? phv_data_222 : _GEN_741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_743 = 8'hdf == local_offset ? phv_data_223 : _GEN_742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_744 = 8'he0 == local_offset ? phv_data_224 : _GEN_743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_745 = 8'he1 == local_offset ? phv_data_225 : _GEN_744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_746 = 8'he2 == local_offset ? phv_data_226 : _GEN_745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_747 = 8'he3 == local_offset ? phv_data_227 : _GEN_746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_748 = 8'he4 == local_offset ? phv_data_228 : _GEN_747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_749 = 8'he5 == local_offset ? phv_data_229 : _GEN_748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_750 = 8'he6 == local_offset ? phv_data_230 : _GEN_749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_751 = 8'he7 == local_offset ? phv_data_231 : _GEN_750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_752 = 8'he8 == local_offset ? phv_data_232 : _GEN_751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_753 = 8'he9 == local_offset ? phv_data_233 : _GEN_752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_754 = 8'hea == local_offset ? phv_data_234 : _GEN_753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_755 = 8'heb == local_offset ? phv_data_235 : _GEN_754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_756 = 8'hec == local_offset ? phv_data_236 : _GEN_755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_757 = 8'hed == local_offset ? phv_data_237 : _GEN_756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_758 = 8'hee == local_offset ? phv_data_238 : _GEN_757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_759 = 8'hef == local_offset ? phv_data_239 : _GEN_758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_760 = 8'hf0 == local_offset ? phv_data_240 : _GEN_759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_761 = 8'hf1 == local_offset ? phv_data_241 : _GEN_760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_762 = 8'hf2 == local_offset ? phv_data_242 : _GEN_761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_763 = 8'hf3 == local_offset ? phv_data_243 : _GEN_762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_764 = 8'hf4 == local_offset ? phv_data_244 : _GEN_763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_765 = 8'hf5 == local_offset ? phv_data_245 : _GEN_764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_766 = 8'hf6 == local_offset ? phv_data_246 : _GEN_765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_767 = 8'hf7 == local_offset ? phv_data_247 : _GEN_766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_768 = 8'hf8 == local_offset ? phv_data_248 : _GEN_767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_769 = 8'hf9 == local_offset ? phv_data_249 : _GEN_768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_770 = 8'hfa == local_offset ? phv_data_250 : _GEN_769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_771 = 8'hfb == local_offset ? phv_data_251 : _GEN_770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_772 = 8'hfc == local_offset ? phv_data_252 : _GEN_771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_773 = 8'hfd == local_offset ? phv_data_253 : _GEN_772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_774 = 8'hfe == local_offset ? phv_data_254 : _GEN_773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_775 = 8'hff == local_offset ? phv_data_255 : _GEN_774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_12582 = {{1'd0}, local_offset}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_776 = 9'h100 == _GEN_12582 ? phv_data_256 : _GEN_775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_777 = 9'h101 == _GEN_12582 ? phv_data_257 : _GEN_776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_778 = 9'h102 == _GEN_12582 ? phv_data_258 : _GEN_777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_779 = 9'h103 == _GEN_12582 ? phv_data_259 : _GEN_778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_780 = 9'h104 == _GEN_12582 ? phv_data_260 : _GEN_779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_781 = 9'h105 == _GEN_12582 ? phv_data_261 : _GEN_780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_782 = 9'h106 == _GEN_12582 ? phv_data_262 : _GEN_781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_783 = 9'h107 == _GEN_12582 ? phv_data_263 : _GEN_782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_784 = 9'h108 == _GEN_12582 ? phv_data_264 : _GEN_783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_785 = 9'h109 == _GEN_12582 ? phv_data_265 : _GEN_784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_786 = 9'h10a == _GEN_12582 ? phv_data_266 : _GEN_785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_787 = 9'h10b == _GEN_12582 ? phv_data_267 : _GEN_786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_788 = 9'h10c == _GEN_12582 ? phv_data_268 : _GEN_787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_789 = 9'h10d == _GEN_12582 ? phv_data_269 : _GEN_788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_790 = 9'h10e == _GEN_12582 ? phv_data_270 : _GEN_789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_791 = 9'h10f == _GEN_12582 ? phv_data_271 : _GEN_790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_792 = 9'h110 == _GEN_12582 ? phv_data_272 : _GEN_791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_793 = 9'h111 == _GEN_12582 ? phv_data_273 : _GEN_792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_794 = 9'h112 == _GEN_12582 ? phv_data_274 : _GEN_793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_795 = 9'h113 == _GEN_12582 ? phv_data_275 : _GEN_794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_796 = 9'h114 == _GEN_12582 ? phv_data_276 : _GEN_795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_797 = 9'h115 == _GEN_12582 ? phv_data_277 : _GEN_796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_798 = 9'h116 == _GEN_12582 ? phv_data_278 : _GEN_797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_799 = 9'h117 == _GEN_12582 ? phv_data_279 : _GEN_798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_800 = 9'h118 == _GEN_12582 ? phv_data_280 : _GEN_799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_801 = 9'h119 == _GEN_12582 ? phv_data_281 : _GEN_800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_802 = 9'h11a == _GEN_12582 ? phv_data_282 : _GEN_801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_803 = 9'h11b == _GEN_12582 ? phv_data_283 : _GEN_802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_804 = 9'h11c == _GEN_12582 ? phv_data_284 : _GEN_803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_805 = 9'h11d == _GEN_12582 ? phv_data_285 : _GEN_804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_806 = 9'h11e == _GEN_12582 ? phv_data_286 : _GEN_805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_807 = 9'h11f == _GEN_12582 ? phv_data_287 : _GEN_806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_808 = 9'h120 == _GEN_12582 ? phv_data_288 : _GEN_807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_809 = 9'h121 == _GEN_12582 ? phv_data_289 : _GEN_808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_810 = 9'h122 == _GEN_12582 ? phv_data_290 : _GEN_809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_811 = 9'h123 == _GEN_12582 ? phv_data_291 : _GEN_810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_812 = 9'h124 == _GEN_12582 ? phv_data_292 : _GEN_811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_813 = 9'h125 == _GEN_12582 ? phv_data_293 : _GEN_812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_814 = 9'h126 == _GEN_12582 ? phv_data_294 : _GEN_813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_815 = 9'h127 == _GEN_12582 ? phv_data_295 : _GEN_814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_816 = 9'h128 == _GEN_12582 ? phv_data_296 : _GEN_815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_817 = 9'h129 == _GEN_12582 ? phv_data_297 : _GEN_816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_818 = 9'h12a == _GEN_12582 ? phv_data_298 : _GEN_817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_819 = 9'h12b == _GEN_12582 ? phv_data_299 : _GEN_818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_820 = 9'h12c == _GEN_12582 ? phv_data_300 : _GEN_819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_821 = 9'h12d == _GEN_12582 ? phv_data_301 : _GEN_820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_822 = 9'h12e == _GEN_12582 ? phv_data_302 : _GEN_821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_823 = 9'h12f == _GEN_12582 ? phv_data_303 : _GEN_822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_824 = 9'h130 == _GEN_12582 ? phv_data_304 : _GEN_823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_825 = 9'h131 == _GEN_12582 ? phv_data_305 : _GEN_824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_826 = 9'h132 == _GEN_12582 ? phv_data_306 : _GEN_825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_827 = 9'h133 == _GEN_12582 ? phv_data_307 : _GEN_826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_828 = 9'h134 == _GEN_12582 ? phv_data_308 : _GEN_827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_829 = 9'h135 == _GEN_12582 ? phv_data_309 : _GEN_828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_830 = 9'h136 == _GEN_12582 ? phv_data_310 : _GEN_829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_831 = 9'h137 == _GEN_12582 ? phv_data_311 : _GEN_830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_832 = 9'h138 == _GEN_12582 ? phv_data_312 : _GEN_831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_833 = 9'h139 == _GEN_12582 ? phv_data_313 : _GEN_832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_834 = 9'h13a == _GEN_12582 ? phv_data_314 : _GEN_833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_835 = 9'h13b == _GEN_12582 ? phv_data_315 : _GEN_834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_836 = 9'h13c == _GEN_12582 ? phv_data_316 : _GEN_835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_837 = 9'h13d == _GEN_12582 ? phv_data_317 : _GEN_836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_838 = 9'h13e == _GEN_12582 ? phv_data_318 : _GEN_837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_839 = 9'h13f == _GEN_12582 ? phv_data_319 : _GEN_838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_840 = 9'h140 == _GEN_12582 ? phv_data_320 : _GEN_839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_841 = 9'h141 == _GEN_12582 ? phv_data_321 : _GEN_840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_842 = 9'h142 == _GEN_12582 ? phv_data_322 : _GEN_841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_843 = 9'h143 == _GEN_12582 ? phv_data_323 : _GEN_842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_844 = 9'h144 == _GEN_12582 ? phv_data_324 : _GEN_843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_845 = 9'h145 == _GEN_12582 ? phv_data_325 : _GEN_844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_846 = 9'h146 == _GEN_12582 ? phv_data_326 : _GEN_845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_847 = 9'h147 == _GEN_12582 ? phv_data_327 : _GEN_846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_848 = 9'h148 == _GEN_12582 ? phv_data_328 : _GEN_847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_849 = 9'h149 == _GEN_12582 ? phv_data_329 : _GEN_848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_850 = 9'h14a == _GEN_12582 ? phv_data_330 : _GEN_849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_851 = 9'h14b == _GEN_12582 ? phv_data_331 : _GEN_850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_852 = 9'h14c == _GEN_12582 ? phv_data_332 : _GEN_851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_853 = 9'h14d == _GEN_12582 ? phv_data_333 : _GEN_852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_854 = 9'h14e == _GEN_12582 ? phv_data_334 : _GEN_853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_855 = 9'h14f == _GEN_12582 ? phv_data_335 : _GEN_854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_856 = 9'h150 == _GEN_12582 ? phv_data_336 : _GEN_855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_857 = 9'h151 == _GEN_12582 ? phv_data_337 : _GEN_856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_858 = 9'h152 == _GEN_12582 ? phv_data_338 : _GEN_857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_859 = 9'h153 == _GEN_12582 ? phv_data_339 : _GEN_858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_860 = 9'h154 == _GEN_12582 ? phv_data_340 : _GEN_859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_861 = 9'h155 == _GEN_12582 ? phv_data_341 : _GEN_860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_862 = 9'h156 == _GEN_12582 ? phv_data_342 : _GEN_861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_863 = 9'h157 == _GEN_12582 ? phv_data_343 : _GEN_862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_864 = 9'h158 == _GEN_12582 ? phv_data_344 : _GEN_863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_865 = 9'h159 == _GEN_12582 ? phv_data_345 : _GEN_864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_866 = 9'h15a == _GEN_12582 ? phv_data_346 : _GEN_865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_867 = 9'h15b == _GEN_12582 ? phv_data_347 : _GEN_866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_868 = 9'h15c == _GEN_12582 ? phv_data_348 : _GEN_867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_869 = 9'h15d == _GEN_12582 ? phv_data_349 : _GEN_868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_870 = 9'h15e == _GEN_12582 ? phv_data_350 : _GEN_869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_871 = 9'h15f == _GEN_12582 ? phv_data_351 : _GEN_870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_872 = 9'h160 == _GEN_12582 ? phv_data_352 : _GEN_871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_873 = 9'h161 == _GEN_12582 ? phv_data_353 : _GEN_872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_874 = 9'h162 == _GEN_12582 ? phv_data_354 : _GEN_873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_875 = 9'h163 == _GEN_12582 ? phv_data_355 : _GEN_874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_876 = 9'h164 == _GEN_12582 ? phv_data_356 : _GEN_875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_877 = 9'h165 == _GEN_12582 ? phv_data_357 : _GEN_876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_878 = 9'h166 == _GEN_12582 ? phv_data_358 : _GEN_877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_879 = 9'h167 == _GEN_12582 ? phv_data_359 : _GEN_878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_880 = 9'h168 == _GEN_12582 ? phv_data_360 : _GEN_879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_881 = 9'h169 == _GEN_12582 ? phv_data_361 : _GEN_880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_882 = 9'h16a == _GEN_12582 ? phv_data_362 : _GEN_881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_883 = 9'h16b == _GEN_12582 ? phv_data_363 : _GEN_882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_884 = 9'h16c == _GEN_12582 ? phv_data_364 : _GEN_883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_885 = 9'h16d == _GEN_12582 ? phv_data_365 : _GEN_884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_886 = 9'h16e == _GEN_12582 ? phv_data_366 : _GEN_885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_887 = 9'h16f == _GEN_12582 ? phv_data_367 : _GEN_886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_888 = 9'h170 == _GEN_12582 ? phv_data_368 : _GEN_887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_889 = 9'h171 == _GEN_12582 ? phv_data_369 : _GEN_888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_890 = 9'h172 == _GEN_12582 ? phv_data_370 : _GEN_889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_891 = 9'h173 == _GEN_12582 ? phv_data_371 : _GEN_890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_892 = 9'h174 == _GEN_12582 ? phv_data_372 : _GEN_891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_893 = 9'h175 == _GEN_12582 ? phv_data_373 : _GEN_892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_894 = 9'h176 == _GEN_12582 ? phv_data_374 : _GEN_893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_895 = 9'h177 == _GEN_12582 ? phv_data_375 : _GEN_894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_896 = 9'h178 == _GEN_12582 ? phv_data_376 : _GEN_895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_897 = 9'h179 == _GEN_12582 ? phv_data_377 : _GEN_896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_898 = 9'h17a == _GEN_12582 ? phv_data_378 : _GEN_897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_899 = 9'h17b == _GEN_12582 ? phv_data_379 : _GEN_898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_900 = 9'h17c == _GEN_12582 ? phv_data_380 : _GEN_899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_901 = 9'h17d == _GEN_12582 ? phv_data_381 : _GEN_900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_902 = 9'h17e == _GEN_12582 ? phv_data_382 : _GEN_901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_903 = 9'h17f == _GEN_12582 ? phv_data_383 : _GEN_902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_904 = 9'h180 == _GEN_12582 ? phv_data_384 : _GEN_903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_905 = 9'h181 == _GEN_12582 ? phv_data_385 : _GEN_904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_906 = 9'h182 == _GEN_12582 ? phv_data_386 : _GEN_905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_907 = 9'h183 == _GEN_12582 ? phv_data_387 : _GEN_906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_908 = 9'h184 == _GEN_12582 ? phv_data_388 : _GEN_907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_909 = 9'h185 == _GEN_12582 ? phv_data_389 : _GEN_908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_910 = 9'h186 == _GEN_12582 ? phv_data_390 : _GEN_909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_911 = 9'h187 == _GEN_12582 ? phv_data_391 : _GEN_910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_912 = 9'h188 == _GEN_12582 ? phv_data_392 : _GEN_911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_913 = 9'h189 == _GEN_12582 ? phv_data_393 : _GEN_912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_914 = 9'h18a == _GEN_12582 ? phv_data_394 : _GEN_913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_915 = 9'h18b == _GEN_12582 ? phv_data_395 : _GEN_914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_916 = 9'h18c == _GEN_12582 ? phv_data_396 : _GEN_915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_917 = 9'h18d == _GEN_12582 ? phv_data_397 : _GEN_916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_918 = 9'h18e == _GEN_12582 ? phv_data_398 : _GEN_917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_919 = 9'h18f == _GEN_12582 ? phv_data_399 : _GEN_918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_920 = 9'h190 == _GEN_12582 ? phv_data_400 : _GEN_919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_921 = 9'h191 == _GEN_12582 ? phv_data_401 : _GEN_920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_922 = 9'h192 == _GEN_12582 ? phv_data_402 : _GEN_921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_923 = 9'h193 == _GEN_12582 ? phv_data_403 : _GEN_922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_924 = 9'h194 == _GEN_12582 ? phv_data_404 : _GEN_923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_925 = 9'h195 == _GEN_12582 ? phv_data_405 : _GEN_924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_926 = 9'h196 == _GEN_12582 ? phv_data_406 : _GEN_925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_927 = 9'h197 == _GEN_12582 ? phv_data_407 : _GEN_926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_928 = 9'h198 == _GEN_12582 ? phv_data_408 : _GEN_927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_929 = 9'h199 == _GEN_12582 ? phv_data_409 : _GEN_928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_930 = 9'h19a == _GEN_12582 ? phv_data_410 : _GEN_929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_931 = 9'h19b == _GEN_12582 ? phv_data_411 : _GEN_930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_932 = 9'h19c == _GEN_12582 ? phv_data_412 : _GEN_931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_933 = 9'h19d == _GEN_12582 ? phv_data_413 : _GEN_932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_934 = 9'h19e == _GEN_12582 ? phv_data_414 : _GEN_933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_935 = 9'h19f == _GEN_12582 ? phv_data_415 : _GEN_934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_936 = 9'h1a0 == _GEN_12582 ? phv_data_416 : _GEN_935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_937 = 9'h1a1 == _GEN_12582 ? phv_data_417 : _GEN_936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_938 = 9'h1a2 == _GEN_12582 ? phv_data_418 : _GEN_937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_939 = 9'h1a3 == _GEN_12582 ? phv_data_419 : _GEN_938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_940 = 9'h1a4 == _GEN_12582 ? phv_data_420 : _GEN_939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_941 = 9'h1a5 == _GEN_12582 ? phv_data_421 : _GEN_940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_942 = 9'h1a6 == _GEN_12582 ? phv_data_422 : _GEN_941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_943 = 9'h1a7 == _GEN_12582 ? phv_data_423 : _GEN_942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_944 = 9'h1a8 == _GEN_12582 ? phv_data_424 : _GEN_943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_945 = 9'h1a9 == _GEN_12582 ? phv_data_425 : _GEN_944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_946 = 9'h1aa == _GEN_12582 ? phv_data_426 : _GEN_945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_947 = 9'h1ab == _GEN_12582 ? phv_data_427 : _GEN_946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_948 = 9'h1ac == _GEN_12582 ? phv_data_428 : _GEN_947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_949 = 9'h1ad == _GEN_12582 ? phv_data_429 : _GEN_948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_950 = 9'h1ae == _GEN_12582 ? phv_data_430 : _GEN_949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_951 = 9'h1af == _GEN_12582 ? phv_data_431 : _GEN_950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_952 = 9'h1b0 == _GEN_12582 ? phv_data_432 : _GEN_951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_953 = 9'h1b1 == _GEN_12582 ? phv_data_433 : _GEN_952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_954 = 9'h1b2 == _GEN_12582 ? phv_data_434 : _GEN_953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_955 = 9'h1b3 == _GEN_12582 ? phv_data_435 : _GEN_954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_956 = 9'h1b4 == _GEN_12582 ? phv_data_436 : _GEN_955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_957 = 9'h1b5 == _GEN_12582 ? phv_data_437 : _GEN_956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_958 = 9'h1b6 == _GEN_12582 ? phv_data_438 : _GEN_957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_959 = 9'h1b7 == _GEN_12582 ? phv_data_439 : _GEN_958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_960 = 9'h1b8 == _GEN_12582 ? phv_data_440 : _GEN_959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_961 = 9'h1b9 == _GEN_12582 ? phv_data_441 : _GEN_960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_962 = 9'h1ba == _GEN_12582 ? phv_data_442 : _GEN_961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_963 = 9'h1bb == _GEN_12582 ? phv_data_443 : _GEN_962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_964 = 9'h1bc == _GEN_12582 ? phv_data_444 : _GEN_963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_965 = 9'h1bd == _GEN_12582 ? phv_data_445 : _GEN_964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_966 = 9'h1be == _GEN_12582 ? phv_data_446 : _GEN_965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_967 = 9'h1bf == _GEN_12582 ? phv_data_447 : _GEN_966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_968 = 9'h1c0 == _GEN_12582 ? phv_data_448 : _GEN_967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_969 = 9'h1c1 == _GEN_12582 ? phv_data_449 : _GEN_968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_970 = 9'h1c2 == _GEN_12582 ? phv_data_450 : _GEN_969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_971 = 9'h1c3 == _GEN_12582 ? phv_data_451 : _GEN_970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_972 = 9'h1c4 == _GEN_12582 ? phv_data_452 : _GEN_971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_973 = 9'h1c5 == _GEN_12582 ? phv_data_453 : _GEN_972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_974 = 9'h1c6 == _GEN_12582 ? phv_data_454 : _GEN_973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_975 = 9'h1c7 == _GEN_12582 ? phv_data_455 : _GEN_974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_976 = 9'h1c8 == _GEN_12582 ? phv_data_456 : _GEN_975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_977 = 9'h1c9 == _GEN_12582 ? phv_data_457 : _GEN_976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_978 = 9'h1ca == _GEN_12582 ? phv_data_458 : _GEN_977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_979 = 9'h1cb == _GEN_12582 ? phv_data_459 : _GEN_978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_980 = 9'h1cc == _GEN_12582 ? phv_data_460 : _GEN_979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_981 = 9'h1cd == _GEN_12582 ? phv_data_461 : _GEN_980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_982 = 9'h1ce == _GEN_12582 ? phv_data_462 : _GEN_981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_983 = 9'h1cf == _GEN_12582 ? phv_data_463 : _GEN_982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_984 = 9'h1d0 == _GEN_12582 ? phv_data_464 : _GEN_983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_985 = 9'h1d1 == _GEN_12582 ? phv_data_465 : _GEN_984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_986 = 9'h1d2 == _GEN_12582 ? phv_data_466 : _GEN_985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_987 = 9'h1d3 == _GEN_12582 ? phv_data_467 : _GEN_986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_988 = 9'h1d4 == _GEN_12582 ? phv_data_468 : _GEN_987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_989 = 9'h1d5 == _GEN_12582 ? phv_data_469 : _GEN_988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_990 = 9'h1d6 == _GEN_12582 ? phv_data_470 : _GEN_989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_991 = 9'h1d7 == _GEN_12582 ? phv_data_471 : _GEN_990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_992 = 9'h1d8 == _GEN_12582 ? phv_data_472 : _GEN_991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_993 = 9'h1d9 == _GEN_12582 ? phv_data_473 : _GEN_992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_994 = 9'h1da == _GEN_12582 ? phv_data_474 : _GEN_993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_995 = 9'h1db == _GEN_12582 ? phv_data_475 : _GEN_994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_996 = 9'h1dc == _GEN_12582 ? phv_data_476 : _GEN_995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_997 = 9'h1dd == _GEN_12582 ? phv_data_477 : _GEN_996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_998 = 9'h1de == _GEN_12582 ? phv_data_478 : _GEN_997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_999 = 9'h1df == _GEN_12582 ? phv_data_479 : _GEN_998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1000 = 9'h1e0 == _GEN_12582 ? phv_data_480 : _GEN_999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1001 = 9'h1e1 == _GEN_12582 ? phv_data_481 : _GEN_1000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1002 = 9'h1e2 == _GEN_12582 ? phv_data_482 : _GEN_1001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1003 = 9'h1e3 == _GEN_12582 ? phv_data_483 : _GEN_1002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1004 = 9'h1e4 == _GEN_12582 ? phv_data_484 : _GEN_1003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1005 = 9'h1e5 == _GEN_12582 ? phv_data_485 : _GEN_1004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1006 = 9'h1e6 == _GEN_12582 ? phv_data_486 : _GEN_1005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1007 = 9'h1e7 == _GEN_12582 ? phv_data_487 : _GEN_1006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1008 = 9'h1e8 == _GEN_12582 ? phv_data_488 : _GEN_1007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1009 = 9'h1e9 == _GEN_12582 ? phv_data_489 : _GEN_1008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1010 = 9'h1ea == _GEN_12582 ? phv_data_490 : _GEN_1009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1011 = 9'h1eb == _GEN_12582 ? phv_data_491 : _GEN_1010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1012 = 9'h1ec == _GEN_12582 ? phv_data_492 : _GEN_1011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1013 = 9'h1ed == _GEN_12582 ? phv_data_493 : _GEN_1012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1014 = 9'h1ee == _GEN_12582 ? phv_data_494 : _GEN_1013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1015 = 9'h1ef == _GEN_12582 ? phv_data_495 : _GEN_1014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1016 = 9'h1f0 == _GEN_12582 ? phv_data_496 : _GEN_1015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1017 = 9'h1f1 == _GEN_12582 ? phv_data_497 : _GEN_1016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1018 = 9'h1f2 == _GEN_12582 ? phv_data_498 : _GEN_1017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1019 = 9'h1f3 == _GEN_12582 ? phv_data_499 : _GEN_1018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1020 = 9'h1f4 == _GEN_12582 ? phv_data_500 : _GEN_1019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1021 = 9'h1f5 == _GEN_12582 ? phv_data_501 : _GEN_1020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1022 = 9'h1f6 == _GEN_12582 ? phv_data_502 : _GEN_1021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1023 = 9'h1f7 == _GEN_12582 ? phv_data_503 : _GEN_1022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1024 = 9'h1f8 == _GEN_12582 ? phv_data_504 : _GEN_1023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1025 = 9'h1f9 == _GEN_12582 ? phv_data_505 : _GEN_1024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1026 = 9'h1fa == _GEN_12582 ? phv_data_506 : _GEN_1025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1027 = 9'h1fb == _GEN_12582 ? phv_data_507 : _GEN_1026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1028 = 9'h1fc == _GEN_12582 ? phv_data_508 : _GEN_1027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1029 = 9'h1fd == _GEN_12582 ? phv_data_509 : _GEN_1028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1030 = 9'h1fe == _GEN_12582 ? phv_data_510 : _GEN_1029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1031 = 9'h1ff == _GEN_12582 ? phv_data_511 : _GEN_1030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1033 = 8'h1 == _match_key_qbytes_0_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1034 = 8'h2 == _match_key_qbytes_0_T ? phv_data_2 : _GEN_1033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1035 = 8'h3 == _match_key_qbytes_0_T ? phv_data_3 : _GEN_1034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1036 = 8'h4 == _match_key_qbytes_0_T ? phv_data_4 : _GEN_1035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1037 = 8'h5 == _match_key_qbytes_0_T ? phv_data_5 : _GEN_1036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1038 = 8'h6 == _match_key_qbytes_0_T ? phv_data_6 : _GEN_1037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1039 = 8'h7 == _match_key_qbytes_0_T ? phv_data_7 : _GEN_1038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1040 = 8'h8 == _match_key_qbytes_0_T ? phv_data_8 : _GEN_1039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1041 = 8'h9 == _match_key_qbytes_0_T ? phv_data_9 : _GEN_1040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1042 = 8'ha == _match_key_qbytes_0_T ? phv_data_10 : _GEN_1041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1043 = 8'hb == _match_key_qbytes_0_T ? phv_data_11 : _GEN_1042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1044 = 8'hc == _match_key_qbytes_0_T ? phv_data_12 : _GEN_1043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1045 = 8'hd == _match_key_qbytes_0_T ? phv_data_13 : _GEN_1044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1046 = 8'he == _match_key_qbytes_0_T ? phv_data_14 : _GEN_1045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1047 = 8'hf == _match_key_qbytes_0_T ? phv_data_15 : _GEN_1046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1048 = 8'h10 == _match_key_qbytes_0_T ? phv_data_16 : _GEN_1047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1049 = 8'h11 == _match_key_qbytes_0_T ? phv_data_17 : _GEN_1048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1050 = 8'h12 == _match_key_qbytes_0_T ? phv_data_18 : _GEN_1049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1051 = 8'h13 == _match_key_qbytes_0_T ? phv_data_19 : _GEN_1050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1052 = 8'h14 == _match_key_qbytes_0_T ? phv_data_20 : _GEN_1051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1053 = 8'h15 == _match_key_qbytes_0_T ? phv_data_21 : _GEN_1052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1054 = 8'h16 == _match_key_qbytes_0_T ? phv_data_22 : _GEN_1053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1055 = 8'h17 == _match_key_qbytes_0_T ? phv_data_23 : _GEN_1054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1056 = 8'h18 == _match_key_qbytes_0_T ? phv_data_24 : _GEN_1055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1057 = 8'h19 == _match_key_qbytes_0_T ? phv_data_25 : _GEN_1056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1058 = 8'h1a == _match_key_qbytes_0_T ? phv_data_26 : _GEN_1057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1059 = 8'h1b == _match_key_qbytes_0_T ? phv_data_27 : _GEN_1058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1060 = 8'h1c == _match_key_qbytes_0_T ? phv_data_28 : _GEN_1059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1061 = 8'h1d == _match_key_qbytes_0_T ? phv_data_29 : _GEN_1060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1062 = 8'h1e == _match_key_qbytes_0_T ? phv_data_30 : _GEN_1061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1063 = 8'h1f == _match_key_qbytes_0_T ? phv_data_31 : _GEN_1062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1064 = 8'h20 == _match_key_qbytes_0_T ? phv_data_32 : _GEN_1063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1065 = 8'h21 == _match_key_qbytes_0_T ? phv_data_33 : _GEN_1064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1066 = 8'h22 == _match_key_qbytes_0_T ? phv_data_34 : _GEN_1065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1067 = 8'h23 == _match_key_qbytes_0_T ? phv_data_35 : _GEN_1066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1068 = 8'h24 == _match_key_qbytes_0_T ? phv_data_36 : _GEN_1067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1069 = 8'h25 == _match_key_qbytes_0_T ? phv_data_37 : _GEN_1068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1070 = 8'h26 == _match_key_qbytes_0_T ? phv_data_38 : _GEN_1069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1071 = 8'h27 == _match_key_qbytes_0_T ? phv_data_39 : _GEN_1070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1072 = 8'h28 == _match_key_qbytes_0_T ? phv_data_40 : _GEN_1071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1073 = 8'h29 == _match_key_qbytes_0_T ? phv_data_41 : _GEN_1072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1074 = 8'h2a == _match_key_qbytes_0_T ? phv_data_42 : _GEN_1073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1075 = 8'h2b == _match_key_qbytes_0_T ? phv_data_43 : _GEN_1074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1076 = 8'h2c == _match_key_qbytes_0_T ? phv_data_44 : _GEN_1075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1077 = 8'h2d == _match_key_qbytes_0_T ? phv_data_45 : _GEN_1076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1078 = 8'h2e == _match_key_qbytes_0_T ? phv_data_46 : _GEN_1077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1079 = 8'h2f == _match_key_qbytes_0_T ? phv_data_47 : _GEN_1078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1080 = 8'h30 == _match_key_qbytes_0_T ? phv_data_48 : _GEN_1079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1081 = 8'h31 == _match_key_qbytes_0_T ? phv_data_49 : _GEN_1080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1082 = 8'h32 == _match_key_qbytes_0_T ? phv_data_50 : _GEN_1081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1083 = 8'h33 == _match_key_qbytes_0_T ? phv_data_51 : _GEN_1082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1084 = 8'h34 == _match_key_qbytes_0_T ? phv_data_52 : _GEN_1083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1085 = 8'h35 == _match_key_qbytes_0_T ? phv_data_53 : _GEN_1084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1086 = 8'h36 == _match_key_qbytes_0_T ? phv_data_54 : _GEN_1085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1087 = 8'h37 == _match_key_qbytes_0_T ? phv_data_55 : _GEN_1086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1088 = 8'h38 == _match_key_qbytes_0_T ? phv_data_56 : _GEN_1087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1089 = 8'h39 == _match_key_qbytes_0_T ? phv_data_57 : _GEN_1088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1090 = 8'h3a == _match_key_qbytes_0_T ? phv_data_58 : _GEN_1089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1091 = 8'h3b == _match_key_qbytes_0_T ? phv_data_59 : _GEN_1090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1092 = 8'h3c == _match_key_qbytes_0_T ? phv_data_60 : _GEN_1091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1093 = 8'h3d == _match_key_qbytes_0_T ? phv_data_61 : _GEN_1092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1094 = 8'h3e == _match_key_qbytes_0_T ? phv_data_62 : _GEN_1093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1095 = 8'h3f == _match_key_qbytes_0_T ? phv_data_63 : _GEN_1094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1096 = 8'h40 == _match_key_qbytes_0_T ? phv_data_64 : _GEN_1095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1097 = 8'h41 == _match_key_qbytes_0_T ? phv_data_65 : _GEN_1096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1098 = 8'h42 == _match_key_qbytes_0_T ? phv_data_66 : _GEN_1097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1099 = 8'h43 == _match_key_qbytes_0_T ? phv_data_67 : _GEN_1098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1100 = 8'h44 == _match_key_qbytes_0_T ? phv_data_68 : _GEN_1099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1101 = 8'h45 == _match_key_qbytes_0_T ? phv_data_69 : _GEN_1100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1102 = 8'h46 == _match_key_qbytes_0_T ? phv_data_70 : _GEN_1101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1103 = 8'h47 == _match_key_qbytes_0_T ? phv_data_71 : _GEN_1102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1104 = 8'h48 == _match_key_qbytes_0_T ? phv_data_72 : _GEN_1103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1105 = 8'h49 == _match_key_qbytes_0_T ? phv_data_73 : _GEN_1104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1106 = 8'h4a == _match_key_qbytes_0_T ? phv_data_74 : _GEN_1105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1107 = 8'h4b == _match_key_qbytes_0_T ? phv_data_75 : _GEN_1106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1108 = 8'h4c == _match_key_qbytes_0_T ? phv_data_76 : _GEN_1107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1109 = 8'h4d == _match_key_qbytes_0_T ? phv_data_77 : _GEN_1108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1110 = 8'h4e == _match_key_qbytes_0_T ? phv_data_78 : _GEN_1109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1111 = 8'h4f == _match_key_qbytes_0_T ? phv_data_79 : _GEN_1110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1112 = 8'h50 == _match_key_qbytes_0_T ? phv_data_80 : _GEN_1111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1113 = 8'h51 == _match_key_qbytes_0_T ? phv_data_81 : _GEN_1112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1114 = 8'h52 == _match_key_qbytes_0_T ? phv_data_82 : _GEN_1113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1115 = 8'h53 == _match_key_qbytes_0_T ? phv_data_83 : _GEN_1114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1116 = 8'h54 == _match_key_qbytes_0_T ? phv_data_84 : _GEN_1115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1117 = 8'h55 == _match_key_qbytes_0_T ? phv_data_85 : _GEN_1116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1118 = 8'h56 == _match_key_qbytes_0_T ? phv_data_86 : _GEN_1117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1119 = 8'h57 == _match_key_qbytes_0_T ? phv_data_87 : _GEN_1118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1120 = 8'h58 == _match_key_qbytes_0_T ? phv_data_88 : _GEN_1119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1121 = 8'h59 == _match_key_qbytes_0_T ? phv_data_89 : _GEN_1120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1122 = 8'h5a == _match_key_qbytes_0_T ? phv_data_90 : _GEN_1121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1123 = 8'h5b == _match_key_qbytes_0_T ? phv_data_91 : _GEN_1122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1124 = 8'h5c == _match_key_qbytes_0_T ? phv_data_92 : _GEN_1123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1125 = 8'h5d == _match_key_qbytes_0_T ? phv_data_93 : _GEN_1124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1126 = 8'h5e == _match_key_qbytes_0_T ? phv_data_94 : _GEN_1125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1127 = 8'h5f == _match_key_qbytes_0_T ? phv_data_95 : _GEN_1126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1128 = 8'h60 == _match_key_qbytes_0_T ? phv_data_96 : _GEN_1127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1129 = 8'h61 == _match_key_qbytes_0_T ? phv_data_97 : _GEN_1128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1130 = 8'h62 == _match_key_qbytes_0_T ? phv_data_98 : _GEN_1129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1131 = 8'h63 == _match_key_qbytes_0_T ? phv_data_99 : _GEN_1130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1132 = 8'h64 == _match_key_qbytes_0_T ? phv_data_100 : _GEN_1131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1133 = 8'h65 == _match_key_qbytes_0_T ? phv_data_101 : _GEN_1132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1134 = 8'h66 == _match_key_qbytes_0_T ? phv_data_102 : _GEN_1133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1135 = 8'h67 == _match_key_qbytes_0_T ? phv_data_103 : _GEN_1134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1136 = 8'h68 == _match_key_qbytes_0_T ? phv_data_104 : _GEN_1135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1137 = 8'h69 == _match_key_qbytes_0_T ? phv_data_105 : _GEN_1136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1138 = 8'h6a == _match_key_qbytes_0_T ? phv_data_106 : _GEN_1137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1139 = 8'h6b == _match_key_qbytes_0_T ? phv_data_107 : _GEN_1138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1140 = 8'h6c == _match_key_qbytes_0_T ? phv_data_108 : _GEN_1139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1141 = 8'h6d == _match_key_qbytes_0_T ? phv_data_109 : _GEN_1140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1142 = 8'h6e == _match_key_qbytes_0_T ? phv_data_110 : _GEN_1141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1143 = 8'h6f == _match_key_qbytes_0_T ? phv_data_111 : _GEN_1142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1144 = 8'h70 == _match_key_qbytes_0_T ? phv_data_112 : _GEN_1143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1145 = 8'h71 == _match_key_qbytes_0_T ? phv_data_113 : _GEN_1144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1146 = 8'h72 == _match_key_qbytes_0_T ? phv_data_114 : _GEN_1145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1147 = 8'h73 == _match_key_qbytes_0_T ? phv_data_115 : _GEN_1146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1148 = 8'h74 == _match_key_qbytes_0_T ? phv_data_116 : _GEN_1147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1149 = 8'h75 == _match_key_qbytes_0_T ? phv_data_117 : _GEN_1148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1150 = 8'h76 == _match_key_qbytes_0_T ? phv_data_118 : _GEN_1149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1151 = 8'h77 == _match_key_qbytes_0_T ? phv_data_119 : _GEN_1150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1152 = 8'h78 == _match_key_qbytes_0_T ? phv_data_120 : _GEN_1151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1153 = 8'h79 == _match_key_qbytes_0_T ? phv_data_121 : _GEN_1152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1154 = 8'h7a == _match_key_qbytes_0_T ? phv_data_122 : _GEN_1153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1155 = 8'h7b == _match_key_qbytes_0_T ? phv_data_123 : _GEN_1154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1156 = 8'h7c == _match_key_qbytes_0_T ? phv_data_124 : _GEN_1155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1157 = 8'h7d == _match_key_qbytes_0_T ? phv_data_125 : _GEN_1156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1158 = 8'h7e == _match_key_qbytes_0_T ? phv_data_126 : _GEN_1157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1159 = 8'h7f == _match_key_qbytes_0_T ? phv_data_127 : _GEN_1158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1160 = 8'h80 == _match_key_qbytes_0_T ? phv_data_128 : _GEN_1159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1161 = 8'h81 == _match_key_qbytes_0_T ? phv_data_129 : _GEN_1160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1162 = 8'h82 == _match_key_qbytes_0_T ? phv_data_130 : _GEN_1161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1163 = 8'h83 == _match_key_qbytes_0_T ? phv_data_131 : _GEN_1162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1164 = 8'h84 == _match_key_qbytes_0_T ? phv_data_132 : _GEN_1163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1165 = 8'h85 == _match_key_qbytes_0_T ? phv_data_133 : _GEN_1164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1166 = 8'h86 == _match_key_qbytes_0_T ? phv_data_134 : _GEN_1165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1167 = 8'h87 == _match_key_qbytes_0_T ? phv_data_135 : _GEN_1166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1168 = 8'h88 == _match_key_qbytes_0_T ? phv_data_136 : _GEN_1167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1169 = 8'h89 == _match_key_qbytes_0_T ? phv_data_137 : _GEN_1168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1170 = 8'h8a == _match_key_qbytes_0_T ? phv_data_138 : _GEN_1169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1171 = 8'h8b == _match_key_qbytes_0_T ? phv_data_139 : _GEN_1170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1172 = 8'h8c == _match_key_qbytes_0_T ? phv_data_140 : _GEN_1171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1173 = 8'h8d == _match_key_qbytes_0_T ? phv_data_141 : _GEN_1172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1174 = 8'h8e == _match_key_qbytes_0_T ? phv_data_142 : _GEN_1173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1175 = 8'h8f == _match_key_qbytes_0_T ? phv_data_143 : _GEN_1174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1176 = 8'h90 == _match_key_qbytes_0_T ? phv_data_144 : _GEN_1175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1177 = 8'h91 == _match_key_qbytes_0_T ? phv_data_145 : _GEN_1176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1178 = 8'h92 == _match_key_qbytes_0_T ? phv_data_146 : _GEN_1177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1179 = 8'h93 == _match_key_qbytes_0_T ? phv_data_147 : _GEN_1178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1180 = 8'h94 == _match_key_qbytes_0_T ? phv_data_148 : _GEN_1179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1181 = 8'h95 == _match_key_qbytes_0_T ? phv_data_149 : _GEN_1180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1182 = 8'h96 == _match_key_qbytes_0_T ? phv_data_150 : _GEN_1181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1183 = 8'h97 == _match_key_qbytes_0_T ? phv_data_151 : _GEN_1182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1184 = 8'h98 == _match_key_qbytes_0_T ? phv_data_152 : _GEN_1183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1185 = 8'h99 == _match_key_qbytes_0_T ? phv_data_153 : _GEN_1184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1186 = 8'h9a == _match_key_qbytes_0_T ? phv_data_154 : _GEN_1185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1187 = 8'h9b == _match_key_qbytes_0_T ? phv_data_155 : _GEN_1186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1188 = 8'h9c == _match_key_qbytes_0_T ? phv_data_156 : _GEN_1187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1189 = 8'h9d == _match_key_qbytes_0_T ? phv_data_157 : _GEN_1188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1190 = 8'h9e == _match_key_qbytes_0_T ? phv_data_158 : _GEN_1189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1191 = 8'h9f == _match_key_qbytes_0_T ? phv_data_159 : _GEN_1190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1192 = 8'ha0 == _match_key_qbytes_0_T ? phv_data_160 : _GEN_1191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1193 = 8'ha1 == _match_key_qbytes_0_T ? phv_data_161 : _GEN_1192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1194 = 8'ha2 == _match_key_qbytes_0_T ? phv_data_162 : _GEN_1193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1195 = 8'ha3 == _match_key_qbytes_0_T ? phv_data_163 : _GEN_1194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1196 = 8'ha4 == _match_key_qbytes_0_T ? phv_data_164 : _GEN_1195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1197 = 8'ha5 == _match_key_qbytes_0_T ? phv_data_165 : _GEN_1196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1198 = 8'ha6 == _match_key_qbytes_0_T ? phv_data_166 : _GEN_1197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1199 = 8'ha7 == _match_key_qbytes_0_T ? phv_data_167 : _GEN_1198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1200 = 8'ha8 == _match_key_qbytes_0_T ? phv_data_168 : _GEN_1199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1201 = 8'ha9 == _match_key_qbytes_0_T ? phv_data_169 : _GEN_1200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1202 = 8'haa == _match_key_qbytes_0_T ? phv_data_170 : _GEN_1201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1203 = 8'hab == _match_key_qbytes_0_T ? phv_data_171 : _GEN_1202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1204 = 8'hac == _match_key_qbytes_0_T ? phv_data_172 : _GEN_1203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1205 = 8'had == _match_key_qbytes_0_T ? phv_data_173 : _GEN_1204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1206 = 8'hae == _match_key_qbytes_0_T ? phv_data_174 : _GEN_1205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1207 = 8'haf == _match_key_qbytes_0_T ? phv_data_175 : _GEN_1206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1208 = 8'hb0 == _match_key_qbytes_0_T ? phv_data_176 : _GEN_1207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1209 = 8'hb1 == _match_key_qbytes_0_T ? phv_data_177 : _GEN_1208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1210 = 8'hb2 == _match_key_qbytes_0_T ? phv_data_178 : _GEN_1209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1211 = 8'hb3 == _match_key_qbytes_0_T ? phv_data_179 : _GEN_1210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1212 = 8'hb4 == _match_key_qbytes_0_T ? phv_data_180 : _GEN_1211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1213 = 8'hb5 == _match_key_qbytes_0_T ? phv_data_181 : _GEN_1212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1214 = 8'hb6 == _match_key_qbytes_0_T ? phv_data_182 : _GEN_1213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1215 = 8'hb7 == _match_key_qbytes_0_T ? phv_data_183 : _GEN_1214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1216 = 8'hb8 == _match_key_qbytes_0_T ? phv_data_184 : _GEN_1215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1217 = 8'hb9 == _match_key_qbytes_0_T ? phv_data_185 : _GEN_1216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1218 = 8'hba == _match_key_qbytes_0_T ? phv_data_186 : _GEN_1217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1219 = 8'hbb == _match_key_qbytes_0_T ? phv_data_187 : _GEN_1218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1220 = 8'hbc == _match_key_qbytes_0_T ? phv_data_188 : _GEN_1219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1221 = 8'hbd == _match_key_qbytes_0_T ? phv_data_189 : _GEN_1220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1222 = 8'hbe == _match_key_qbytes_0_T ? phv_data_190 : _GEN_1221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1223 = 8'hbf == _match_key_qbytes_0_T ? phv_data_191 : _GEN_1222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1224 = 8'hc0 == _match_key_qbytes_0_T ? phv_data_192 : _GEN_1223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1225 = 8'hc1 == _match_key_qbytes_0_T ? phv_data_193 : _GEN_1224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1226 = 8'hc2 == _match_key_qbytes_0_T ? phv_data_194 : _GEN_1225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1227 = 8'hc3 == _match_key_qbytes_0_T ? phv_data_195 : _GEN_1226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1228 = 8'hc4 == _match_key_qbytes_0_T ? phv_data_196 : _GEN_1227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1229 = 8'hc5 == _match_key_qbytes_0_T ? phv_data_197 : _GEN_1228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1230 = 8'hc6 == _match_key_qbytes_0_T ? phv_data_198 : _GEN_1229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1231 = 8'hc7 == _match_key_qbytes_0_T ? phv_data_199 : _GEN_1230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1232 = 8'hc8 == _match_key_qbytes_0_T ? phv_data_200 : _GEN_1231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1233 = 8'hc9 == _match_key_qbytes_0_T ? phv_data_201 : _GEN_1232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1234 = 8'hca == _match_key_qbytes_0_T ? phv_data_202 : _GEN_1233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1235 = 8'hcb == _match_key_qbytes_0_T ? phv_data_203 : _GEN_1234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1236 = 8'hcc == _match_key_qbytes_0_T ? phv_data_204 : _GEN_1235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1237 = 8'hcd == _match_key_qbytes_0_T ? phv_data_205 : _GEN_1236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1238 = 8'hce == _match_key_qbytes_0_T ? phv_data_206 : _GEN_1237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1239 = 8'hcf == _match_key_qbytes_0_T ? phv_data_207 : _GEN_1238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1240 = 8'hd0 == _match_key_qbytes_0_T ? phv_data_208 : _GEN_1239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1241 = 8'hd1 == _match_key_qbytes_0_T ? phv_data_209 : _GEN_1240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1242 = 8'hd2 == _match_key_qbytes_0_T ? phv_data_210 : _GEN_1241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1243 = 8'hd3 == _match_key_qbytes_0_T ? phv_data_211 : _GEN_1242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1244 = 8'hd4 == _match_key_qbytes_0_T ? phv_data_212 : _GEN_1243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1245 = 8'hd5 == _match_key_qbytes_0_T ? phv_data_213 : _GEN_1244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1246 = 8'hd6 == _match_key_qbytes_0_T ? phv_data_214 : _GEN_1245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1247 = 8'hd7 == _match_key_qbytes_0_T ? phv_data_215 : _GEN_1246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1248 = 8'hd8 == _match_key_qbytes_0_T ? phv_data_216 : _GEN_1247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1249 = 8'hd9 == _match_key_qbytes_0_T ? phv_data_217 : _GEN_1248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1250 = 8'hda == _match_key_qbytes_0_T ? phv_data_218 : _GEN_1249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1251 = 8'hdb == _match_key_qbytes_0_T ? phv_data_219 : _GEN_1250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1252 = 8'hdc == _match_key_qbytes_0_T ? phv_data_220 : _GEN_1251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1253 = 8'hdd == _match_key_qbytes_0_T ? phv_data_221 : _GEN_1252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1254 = 8'hde == _match_key_qbytes_0_T ? phv_data_222 : _GEN_1253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1255 = 8'hdf == _match_key_qbytes_0_T ? phv_data_223 : _GEN_1254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1256 = 8'he0 == _match_key_qbytes_0_T ? phv_data_224 : _GEN_1255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1257 = 8'he1 == _match_key_qbytes_0_T ? phv_data_225 : _GEN_1256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1258 = 8'he2 == _match_key_qbytes_0_T ? phv_data_226 : _GEN_1257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1259 = 8'he3 == _match_key_qbytes_0_T ? phv_data_227 : _GEN_1258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1260 = 8'he4 == _match_key_qbytes_0_T ? phv_data_228 : _GEN_1259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1261 = 8'he5 == _match_key_qbytes_0_T ? phv_data_229 : _GEN_1260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1262 = 8'he6 == _match_key_qbytes_0_T ? phv_data_230 : _GEN_1261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1263 = 8'he7 == _match_key_qbytes_0_T ? phv_data_231 : _GEN_1262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1264 = 8'he8 == _match_key_qbytes_0_T ? phv_data_232 : _GEN_1263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1265 = 8'he9 == _match_key_qbytes_0_T ? phv_data_233 : _GEN_1264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1266 = 8'hea == _match_key_qbytes_0_T ? phv_data_234 : _GEN_1265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1267 = 8'heb == _match_key_qbytes_0_T ? phv_data_235 : _GEN_1266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1268 = 8'hec == _match_key_qbytes_0_T ? phv_data_236 : _GEN_1267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1269 = 8'hed == _match_key_qbytes_0_T ? phv_data_237 : _GEN_1268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1270 = 8'hee == _match_key_qbytes_0_T ? phv_data_238 : _GEN_1269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1271 = 8'hef == _match_key_qbytes_0_T ? phv_data_239 : _GEN_1270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1272 = 8'hf0 == _match_key_qbytes_0_T ? phv_data_240 : _GEN_1271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1273 = 8'hf1 == _match_key_qbytes_0_T ? phv_data_241 : _GEN_1272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1274 = 8'hf2 == _match_key_qbytes_0_T ? phv_data_242 : _GEN_1273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1275 = 8'hf3 == _match_key_qbytes_0_T ? phv_data_243 : _GEN_1274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1276 = 8'hf4 == _match_key_qbytes_0_T ? phv_data_244 : _GEN_1275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1277 = 8'hf5 == _match_key_qbytes_0_T ? phv_data_245 : _GEN_1276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1278 = 8'hf6 == _match_key_qbytes_0_T ? phv_data_246 : _GEN_1277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1279 = 8'hf7 == _match_key_qbytes_0_T ? phv_data_247 : _GEN_1278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1280 = 8'hf8 == _match_key_qbytes_0_T ? phv_data_248 : _GEN_1279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1281 = 8'hf9 == _match_key_qbytes_0_T ? phv_data_249 : _GEN_1280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1282 = 8'hfa == _match_key_qbytes_0_T ? phv_data_250 : _GEN_1281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1283 = 8'hfb == _match_key_qbytes_0_T ? phv_data_251 : _GEN_1282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1284 = 8'hfc == _match_key_qbytes_0_T ? phv_data_252 : _GEN_1283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1285 = 8'hfd == _match_key_qbytes_0_T ? phv_data_253 : _GEN_1284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1286 = 8'hfe == _match_key_qbytes_0_T ? phv_data_254 : _GEN_1285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1287 = 8'hff == _match_key_qbytes_0_T ? phv_data_255 : _GEN_1286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_12838 = {{1'd0}, _match_key_qbytes_0_T}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1288 = 9'h100 == _GEN_12838 ? phv_data_256 : _GEN_1287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1289 = 9'h101 == _GEN_12838 ? phv_data_257 : _GEN_1288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1290 = 9'h102 == _GEN_12838 ? phv_data_258 : _GEN_1289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1291 = 9'h103 == _GEN_12838 ? phv_data_259 : _GEN_1290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1292 = 9'h104 == _GEN_12838 ? phv_data_260 : _GEN_1291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1293 = 9'h105 == _GEN_12838 ? phv_data_261 : _GEN_1292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1294 = 9'h106 == _GEN_12838 ? phv_data_262 : _GEN_1293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1295 = 9'h107 == _GEN_12838 ? phv_data_263 : _GEN_1294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1296 = 9'h108 == _GEN_12838 ? phv_data_264 : _GEN_1295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1297 = 9'h109 == _GEN_12838 ? phv_data_265 : _GEN_1296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1298 = 9'h10a == _GEN_12838 ? phv_data_266 : _GEN_1297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1299 = 9'h10b == _GEN_12838 ? phv_data_267 : _GEN_1298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1300 = 9'h10c == _GEN_12838 ? phv_data_268 : _GEN_1299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1301 = 9'h10d == _GEN_12838 ? phv_data_269 : _GEN_1300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1302 = 9'h10e == _GEN_12838 ? phv_data_270 : _GEN_1301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1303 = 9'h10f == _GEN_12838 ? phv_data_271 : _GEN_1302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1304 = 9'h110 == _GEN_12838 ? phv_data_272 : _GEN_1303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1305 = 9'h111 == _GEN_12838 ? phv_data_273 : _GEN_1304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1306 = 9'h112 == _GEN_12838 ? phv_data_274 : _GEN_1305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1307 = 9'h113 == _GEN_12838 ? phv_data_275 : _GEN_1306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1308 = 9'h114 == _GEN_12838 ? phv_data_276 : _GEN_1307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1309 = 9'h115 == _GEN_12838 ? phv_data_277 : _GEN_1308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1310 = 9'h116 == _GEN_12838 ? phv_data_278 : _GEN_1309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1311 = 9'h117 == _GEN_12838 ? phv_data_279 : _GEN_1310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1312 = 9'h118 == _GEN_12838 ? phv_data_280 : _GEN_1311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1313 = 9'h119 == _GEN_12838 ? phv_data_281 : _GEN_1312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1314 = 9'h11a == _GEN_12838 ? phv_data_282 : _GEN_1313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1315 = 9'h11b == _GEN_12838 ? phv_data_283 : _GEN_1314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1316 = 9'h11c == _GEN_12838 ? phv_data_284 : _GEN_1315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1317 = 9'h11d == _GEN_12838 ? phv_data_285 : _GEN_1316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1318 = 9'h11e == _GEN_12838 ? phv_data_286 : _GEN_1317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1319 = 9'h11f == _GEN_12838 ? phv_data_287 : _GEN_1318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1320 = 9'h120 == _GEN_12838 ? phv_data_288 : _GEN_1319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1321 = 9'h121 == _GEN_12838 ? phv_data_289 : _GEN_1320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1322 = 9'h122 == _GEN_12838 ? phv_data_290 : _GEN_1321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1323 = 9'h123 == _GEN_12838 ? phv_data_291 : _GEN_1322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1324 = 9'h124 == _GEN_12838 ? phv_data_292 : _GEN_1323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1325 = 9'h125 == _GEN_12838 ? phv_data_293 : _GEN_1324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1326 = 9'h126 == _GEN_12838 ? phv_data_294 : _GEN_1325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1327 = 9'h127 == _GEN_12838 ? phv_data_295 : _GEN_1326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1328 = 9'h128 == _GEN_12838 ? phv_data_296 : _GEN_1327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1329 = 9'h129 == _GEN_12838 ? phv_data_297 : _GEN_1328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1330 = 9'h12a == _GEN_12838 ? phv_data_298 : _GEN_1329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1331 = 9'h12b == _GEN_12838 ? phv_data_299 : _GEN_1330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1332 = 9'h12c == _GEN_12838 ? phv_data_300 : _GEN_1331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1333 = 9'h12d == _GEN_12838 ? phv_data_301 : _GEN_1332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1334 = 9'h12e == _GEN_12838 ? phv_data_302 : _GEN_1333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1335 = 9'h12f == _GEN_12838 ? phv_data_303 : _GEN_1334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1336 = 9'h130 == _GEN_12838 ? phv_data_304 : _GEN_1335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1337 = 9'h131 == _GEN_12838 ? phv_data_305 : _GEN_1336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1338 = 9'h132 == _GEN_12838 ? phv_data_306 : _GEN_1337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1339 = 9'h133 == _GEN_12838 ? phv_data_307 : _GEN_1338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1340 = 9'h134 == _GEN_12838 ? phv_data_308 : _GEN_1339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1341 = 9'h135 == _GEN_12838 ? phv_data_309 : _GEN_1340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1342 = 9'h136 == _GEN_12838 ? phv_data_310 : _GEN_1341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1343 = 9'h137 == _GEN_12838 ? phv_data_311 : _GEN_1342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1344 = 9'h138 == _GEN_12838 ? phv_data_312 : _GEN_1343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1345 = 9'h139 == _GEN_12838 ? phv_data_313 : _GEN_1344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1346 = 9'h13a == _GEN_12838 ? phv_data_314 : _GEN_1345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1347 = 9'h13b == _GEN_12838 ? phv_data_315 : _GEN_1346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1348 = 9'h13c == _GEN_12838 ? phv_data_316 : _GEN_1347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1349 = 9'h13d == _GEN_12838 ? phv_data_317 : _GEN_1348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1350 = 9'h13e == _GEN_12838 ? phv_data_318 : _GEN_1349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1351 = 9'h13f == _GEN_12838 ? phv_data_319 : _GEN_1350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1352 = 9'h140 == _GEN_12838 ? phv_data_320 : _GEN_1351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1353 = 9'h141 == _GEN_12838 ? phv_data_321 : _GEN_1352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1354 = 9'h142 == _GEN_12838 ? phv_data_322 : _GEN_1353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1355 = 9'h143 == _GEN_12838 ? phv_data_323 : _GEN_1354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1356 = 9'h144 == _GEN_12838 ? phv_data_324 : _GEN_1355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1357 = 9'h145 == _GEN_12838 ? phv_data_325 : _GEN_1356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1358 = 9'h146 == _GEN_12838 ? phv_data_326 : _GEN_1357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1359 = 9'h147 == _GEN_12838 ? phv_data_327 : _GEN_1358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1360 = 9'h148 == _GEN_12838 ? phv_data_328 : _GEN_1359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1361 = 9'h149 == _GEN_12838 ? phv_data_329 : _GEN_1360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1362 = 9'h14a == _GEN_12838 ? phv_data_330 : _GEN_1361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1363 = 9'h14b == _GEN_12838 ? phv_data_331 : _GEN_1362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1364 = 9'h14c == _GEN_12838 ? phv_data_332 : _GEN_1363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1365 = 9'h14d == _GEN_12838 ? phv_data_333 : _GEN_1364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1366 = 9'h14e == _GEN_12838 ? phv_data_334 : _GEN_1365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1367 = 9'h14f == _GEN_12838 ? phv_data_335 : _GEN_1366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1368 = 9'h150 == _GEN_12838 ? phv_data_336 : _GEN_1367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1369 = 9'h151 == _GEN_12838 ? phv_data_337 : _GEN_1368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1370 = 9'h152 == _GEN_12838 ? phv_data_338 : _GEN_1369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1371 = 9'h153 == _GEN_12838 ? phv_data_339 : _GEN_1370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1372 = 9'h154 == _GEN_12838 ? phv_data_340 : _GEN_1371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1373 = 9'h155 == _GEN_12838 ? phv_data_341 : _GEN_1372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1374 = 9'h156 == _GEN_12838 ? phv_data_342 : _GEN_1373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1375 = 9'h157 == _GEN_12838 ? phv_data_343 : _GEN_1374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1376 = 9'h158 == _GEN_12838 ? phv_data_344 : _GEN_1375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1377 = 9'h159 == _GEN_12838 ? phv_data_345 : _GEN_1376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1378 = 9'h15a == _GEN_12838 ? phv_data_346 : _GEN_1377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1379 = 9'h15b == _GEN_12838 ? phv_data_347 : _GEN_1378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1380 = 9'h15c == _GEN_12838 ? phv_data_348 : _GEN_1379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1381 = 9'h15d == _GEN_12838 ? phv_data_349 : _GEN_1380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1382 = 9'h15e == _GEN_12838 ? phv_data_350 : _GEN_1381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1383 = 9'h15f == _GEN_12838 ? phv_data_351 : _GEN_1382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1384 = 9'h160 == _GEN_12838 ? phv_data_352 : _GEN_1383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1385 = 9'h161 == _GEN_12838 ? phv_data_353 : _GEN_1384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1386 = 9'h162 == _GEN_12838 ? phv_data_354 : _GEN_1385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1387 = 9'h163 == _GEN_12838 ? phv_data_355 : _GEN_1386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1388 = 9'h164 == _GEN_12838 ? phv_data_356 : _GEN_1387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1389 = 9'h165 == _GEN_12838 ? phv_data_357 : _GEN_1388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1390 = 9'h166 == _GEN_12838 ? phv_data_358 : _GEN_1389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1391 = 9'h167 == _GEN_12838 ? phv_data_359 : _GEN_1390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1392 = 9'h168 == _GEN_12838 ? phv_data_360 : _GEN_1391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1393 = 9'h169 == _GEN_12838 ? phv_data_361 : _GEN_1392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1394 = 9'h16a == _GEN_12838 ? phv_data_362 : _GEN_1393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1395 = 9'h16b == _GEN_12838 ? phv_data_363 : _GEN_1394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1396 = 9'h16c == _GEN_12838 ? phv_data_364 : _GEN_1395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1397 = 9'h16d == _GEN_12838 ? phv_data_365 : _GEN_1396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1398 = 9'h16e == _GEN_12838 ? phv_data_366 : _GEN_1397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1399 = 9'h16f == _GEN_12838 ? phv_data_367 : _GEN_1398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1400 = 9'h170 == _GEN_12838 ? phv_data_368 : _GEN_1399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1401 = 9'h171 == _GEN_12838 ? phv_data_369 : _GEN_1400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1402 = 9'h172 == _GEN_12838 ? phv_data_370 : _GEN_1401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1403 = 9'h173 == _GEN_12838 ? phv_data_371 : _GEN_1402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1404 = 9'h174 == _GEN_12838 ? phv_data_372 : _GEN_1403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1405 = 9'h175 == _GEN_12838 ? phv_data_373 : _GEN_1404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1406 = 9'h176 == _GEN_12838 ? phv_data_374 : _GEN_1405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1407 = 9'h177 == _GEN_12838 ? phv_data_375 : _GEN_1406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1408 = 9'h178 == _GEN_12838 ? phv_data_376 : _GEN_1407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1409 = 9'h179 == _GEN_12838 ? phv_data_377 : _GEN_1408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1410 = 9'h17a == _GEN_12838 ? phv_data_378 : _GEN_1409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1411 = 9'h17b == _GEN_12838 ? phv_data_379 : _GEN_1410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1412 = 9'h17c == _GEN_12838 ? phv_data_380 : _GEN_1411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1413 = 9'h17d == _GEN_12838 ? phv_data_381 : _GEN_1412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1414 = 9'h17e == _GEN_12838 ? phv_data_382 : _GEN_1413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1415 = 9'h17f == _GEN_12838 ? phv_data_383 : _GEN_1414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1416 = 9'h180 == _GEN_12838 ? phv_data_384 : _GEN_1415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1417 = 9'h181 == _GEN_12838 ? phv_data_385 : _GEN_1416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1418 = 9'h182 == _GEN_12838 ? phv_data_386 : _GEN_1417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1419 = 9'h183 == _GEN_12838 ? phv_data_387 : _GEN_1418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1420 = 9'h184 == _GEN_12838 ? phv_data_388 : _GEN_1419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1421 = 9'h185 == _GEN_12838 ? phv_data_389 : _GEN_1420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1422 = 9'h186 == _GEN_12838 ? phv_data_390 : _GEN_1421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1423 = 9'h187 == _GEN_12838 ? phv_data_391 : _GEN_1422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1424 = 9'h188 == _GEN_12838 ? phv_data_392 : _GEN_1423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1425 = 9'h189 == _GEN_12838 ? phv_data_393 : _GEN_1424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1426 = 9'h18a == _GEN_12838 ? phv_data_394 : _GEN_1425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1427 = 9'h18b == _GEN_12838 ? phv_data_395 : _GEN_1426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1428 = 9'h18c == _GEN_12838 ? phv_data_396 : _GEN_1427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1429 = 9'h18d == _GEN_12838 ? phv_data_397 : _GEN_1428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1430 = 9'h18e == _GEN_12838 ? phv_data_398 : _GEN_1429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1431 = 9'h18f == _GEN_12838 ? phv_data_399 : _GEN_1430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1432 = 9'h190 == _GEN_12838 ? phv_data_400 : _GEN_1431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1433 = 9'h191 == _GEN_12838 ? phv_data_401 : _GEN_1432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1434 = 9'h192 == _GEN_12838 ? phv_data_402 : _GEN_1433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1435 = 9'h193 == _GEN_12838 ? phv_data_403 : _GEN_1434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1436 = 9'h194 == _GEN_12838 ? phv_data_404 : _GEN_1435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1437 = 9'h195 == _GEN_12838 ? phv_data_405 : _GEN_1436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1438 = 9'h196 == _GEN_12838 ? phv_data_406 : _GEN_1437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1439 = 9'h197 == _GEN_12838 ? phv_data_407 : _GEN_1438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1440 = 9'h198 == _GEN_12838 ? phv_data_408 : _GEN_1439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1441 = 9'h199 == _GEN_12838 ? phv_data_409 : _GEN_1440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1442 = 9'h19a == _GEN_12838 ? phv_data_410 : _GEN_1441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1443 = 9'h19b == _GEN_12838 ? phv_data_411 : _GEN_1442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1444 = 9'h19c == _GEN_12838 ? phv_data_412 : _GEN_1443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1445 = 9'h19d == _GEN_12838 ? phv_data_413 : _GEN_1444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1446 = 9'h19e == _GEN_12838 ? phv_data_414 : _GEN_1445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1447 = 9'h19f == _GEN_12838 ? phv_data_415 : _GEN_1446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1448 = 9'h1a0 == _GEN_12838 ? phv_data_416 : _GEN_1447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1449 = 9'h1a1 == _GEN_12838 ? phv_data_417 : _GEN_1448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1450 = 9'h1a2 == _GEN_12838 ? phv_data_418 : _GEN_1449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1451 = 9'h1a3 == _GEN_12838 ? phv_data_419 : _GEN_1450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1452 = 9'h1a4 == _GEN_12838 ? phv_data_420 : _GEN_1451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1453 = 9'h1a5 == _GEN_12838 ? phv_data_421 : _GEN_1452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1454 = 9'h1a6 == _GEN_12838 ? phv_data_422 : _GEN_1453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1455 = 9'h1a7 == _GEN_12838 ? phv_data_423 : _GEN_1454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1456 = 9'h1a8 == _GEN_12838 ? phv_data_424 : _GEN_1455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1457 = 9'h1a9 == _GEN_12838 ? phv_data_425 : _GEN_1456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1458 = 9'h1aa == _GEN_12838 ? phv_data_426 : _GEN_1457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1459 = 9'h1ab == _GEN_12838 ? phv_data_427 : _GEN_1458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1460 = 9'h1ac == _GEN_12838 ? phv_data_428 : _GEN_1459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1461 = 9'h1ad == _GEN_12838 ? phv_data_429 : _GEN_1460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1462 = 9'h1ae == _GEN_12838 ? phv_data_430 : _GEN_1461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1463 = 9'h1af == _GEN_12838 ? phv_data_431 : _GEN_1462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1464 = 9'h1b0 == _GEN_12838 ? phv_data_432 : _GEN_1463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1465 = 9'h1b1 == _GEN_12838 ? phv_data_433 : _GEN_1464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1466 = 9'h1b2 == _GEN_12838 ? phv_data_434 : _GEN_1465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1467 = 9'h1b3 == _GEN_12838 ? phv_data_435 : _GEN_1466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1468 = 9'h1b4 == _GEN_12838 ? phv_data_436 : _GEN_1467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1469 = 9'h1b5 == _GEN_12838 ? phv_data_437 : _GEN_1468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1470 = 9'h1b6 == _GEN_12838 ? phv_data_438 : _GEN_1469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1471 = 9'h1b7 == _GEN_12838 ? phv_data_439 : _GEN_1470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1472 = 9'h1b8 == _GEN_12838 ? phv_data_440 : _GEN_1471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1473 = 9'h1b9 == _GEN_12838 ? phv_data_441 : _GEN_1472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1474 = 9'h1ba == _GEN_12838 ? phv_data_442 : _GEN_1473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1475 = 9'h1bb == _GEN_12838 ? phv_data_443 : _GEN_1474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1476 = 9'h1bc == _GEN_12838 ? phv_data_444 : _GEN_1475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1477 = 9'h1bd == _GEN_12838 ? phv_data_445 : _GEN_1476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1478 = 9'h1be == _GEN_12838 ? phv_data_446 : _GEN_1477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1479 = 9'h1bf == _GEN_12838 ? phv_data_447 : _GEN_1478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1480 = 9'h1c0 == _GEN_12838 ? phv_data_448 : _GEN_1479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1481 = 9'h1c1 == _GEN_12838 ? phv_data_449 : _GEN_1480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1482 = 9'h1c2 == _GEN_12838 ? phv_data_450 : _GEN_1481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1483 = 9'h1c3 == _GEN_12838 ? phv_data_451 : _GEN_1482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1484 = 9'h1c4 == _GEN_12838 ? phv_data_452 : _GEN_1483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1485 = 9'h1c5 == _GEN_12838 ? phv_data_453 : _GEN_1484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1486 = 9'h1c6 == _GEN_12838 ? phv_data_454 : _GEN_1485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1487 = 9'h1c7 == _GEN_12838 ? phv_data_455 : _GEN_1486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1488 = 9'h1c8 == _GEN_12838 ? phv_data_456 : _GEN_1487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1489 = 9'h1c9 == _GEN_12838 ? phv_data_457 : _GEN_1488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1490 = 9'h1ca == _GEN_12838 ? phv_data_458 : _GEN_1489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1491 = 9'h1cb == _GEN_12838 ? phv_data_459 : _GEN_1490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1492 = 9'h1cc == _GEN_12838 ? phv_data_460 : _GEN_1491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1493 = 9'h1cd == _GEN_12838 ? phv_data_461 : _GEN_1492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1494 = 9'h1ce == _GEN_12838 ? phv_data_462 : _GEN_1493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1495 = 9'h1cf == _GEN_12838 ? phv_data_463 : _GEN_1494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1496 = 9'h1d0 == _GEN_12838 ? phv_data_464 : _GEN_1495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1497 = 9'h1d1 == _GEN_12838 ? phv_data_465 : _GEN_1496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1498 = 9'h1d2 == _GEN_12838 ? phv_data_466 : _GEN_1497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1499 = 9'h1d3 == _GEN_12838 ? phv_data_467 : _GEN_1498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1500 = 9'h1d4 == _GEN_12838 ? phv_data_468 : _GEN_1499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1501 = 9'h1d5 == _GEN_12838 ? phv_data_469 : _GEN_1500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1502 = 9'h1d6 == _GEN_12838 ? phv_data_470 : _GEN_1501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1503 = 9'h1d7 == _GEN_12838 ? phv_data_471 : _GEN_1502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1504 = 9'h1d8 == _GEN_12838 ? phv_data_472 : _GEN_1503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1505 = 9'h1d9 == _GEN_12838 ? phv_data_473 : _GEN_1504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1506 = 9'h1da == _GEN_12838 ? phv_data_474 : _GEN_1505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1507 = 9'h1db == _GEN_12838 ? phv_data_475 : _GEN_1506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1508 = 9'h1dc == _GEN_12838 ? phv_data_476 : _GEN_1507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1509 = 9'h1dd == _GEN_12838 ? phv_data_477 : _GEN_1508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1510 = 9'h1de == _GEN_12838 ? phv_data_478 : _GEN_1509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1511 = 9'h1df == _GEN_12838 ? phv_data_479 : _GEN_1510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1512 = 9'h1e0 == _GEN_12838 ? phv_data_480 : _GEN_1511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1513 = 9'h1e1 == _GEN_12838 ? phv_data_481 : _GEN_1512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1514 = 9'h1e2 == _GEN_12838 ? phv_data_482 : _GEN_1513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1515 = 9'h1e3 == _GEN_12838 ? phv_data_483 : _GEN_1514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1516 = 9'h1e4 == _GEN_12838 ? phv_data_484 : _GEN_1515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1517 = 9'h1e5 == _GEN_12838 ? phv_data_485 : _GEN_1516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1518 = 9'h1e6 == _GEN_12838 ? phv_data_486 : _GEN_1517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1519 = 9'h1e7 == _GEN_12838 ? phv_data_487 : _GEN_1518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1520 = 9'h1e8 == _GEN_12838 ? phv_data_488 : _GEN_1519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1521 = 9'h1e9 == _GEN_12838 ? phv_data_489 : _GEN_1520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1522 = 9'h1ea == _GEN_12838 ? phv_data_490 : _GEN_1521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1523 = 9'h1eb == _GEN_12838 ? phv_data_491 : _GEN_1522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1524 = 9'h1ec == _GEN_12838 ? phv_data_492 : _GEN_1523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1525 = 9'h1ed == _GEN_12838 ? phv_data_493 : _GEN_1524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1526 = 9'h1ee == _GEN_12838 ? phv_data_494 : _GEN_1525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1527 = 9'h1ef == _GEN_12838 ? phv_data_495 : _GEN_1526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1528 = 9'h1f0 == _GEN_12838 ? phv_data_496 : _GEN_1527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1529 = 9'h1f1 == _GEN_12838 ? phv_data_497 : _GEN_1528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1530 = 9'h1f2 == _GEN_12838 ? phv_data_498 : _GEN_1529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1531 = 9'h1f3 == _GEN_12838 ? phv_data_499 : _GEN_1530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1532 = 9'h1f4 == _GEN_12838 ? phv_data_500 : _GEN_1531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1533 = 9'h1f5 == _GEN_12838 ? phv_data_501 : _GEN_1532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1534 = 9'h1f6 == _GEN_12838 ? phv_data_502 : _GEN_1533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1535 = 9'h1f7 == _GEN_12838 ? phv_data_503 : _GEN_1534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1536 = 9'h1f8 == _GEN_12838 ? phv_data_504 : _GEN_1535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1537 = 9'h1f9 == _GEN_12838 ? phv_data_505 : _GEN_1536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1538 = 9'h1fa == _GEN_12838 ? phv_data_506 : _GEN_1537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1539 = 9'h1fb == _GEN_12838 ? phv_data_507 : _GEN_1538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1540 = 9'h1fc == _GEN_12838 ? phv_data_508 : _GEN_1539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1541 = 9'h1fd == _GEN_12838 ? phv_data_509 : _GEN_1540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1542 = 9'h1fe == _GEN_12838 ? phv_data_510 : _GEN_1541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1543 = 9'h1ff == _GEN_12838 ? phv_data_511 : _GEN_1542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1545 = 8'h1 == _match_key_qbytes_0_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1546 = 8'h2 == _match_key_qbytes_0_T_1 ? phv_data_2 : _GEN_1545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1547 = 8'h3 == _match_key_qbytes_0_T_1 ? phv_data_3 : _GEN_1546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1548 = 8'h4 == _match_key_qbytes_0_T_1 ? phv_data_4 : _GEN_1547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1549 = 8'h5 == _match_key_qbytes_0_T_1 ? phv_data_5 : _GEN_1548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1550 = 8'h6 == _match_key_qbytes_0_T_1 ? phv_data_6 : _GEN_1549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1551 = 8'h7 == _match_key_qbytes_0_T_1 ? phv_data_7 : _GEN_1550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1552 = 8'h8 == _match_key_qbytes_0_T_1 ? phv_data_8 : _GEN_1551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1553 = 8'h9 == _match_key_qbytes_0_T_1 ? phv_data_9 : _GEN_1552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1554 = 8'ha == _match_key_qbytes_0_T_1 ? phv_data_10 : _GEN_1553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1555 = 8'hb == _match_key_qbytes_0_T_1 ? phv_data_11 : _GEN_1554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1556 = 8'hc == _match_key_qbytes_0_T_1 ? phv_data_12 : _GEN_1555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1557 = 8'hd == _match_key_qbytes_0_T_1 ? phv_data_13 : _GEN_1556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1558 = 8'he == _match_key_qbytes_0_T_1 ? phv_data_14 : _GEN_1557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1559 = 8'hf == _match_key_qbytes_0_T_1 ? phv_data_15 : _GEN_1558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1560 = 8'h10 == _match_key_qbytes_0_T_1 ? phv_data_16 : _GEN_1559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1561 = 8'h11 == _match_key_qbytes_0_T_1 ? phv_data_17 : _GEN_1560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1562 = 8'h12 == _match_key_qbytes_0_T_1 ? phv_data_18 : _GEN_1561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1563 = 8'h13 == _match_key_qbytes_0_T_1 ? phv_data_19 : _GEN_1562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1564 = 8'h14 == _match_key_qbytes_0_T_1 ? phv_data_20 : _GEN_1563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1565 = 8'h15 == _match_key_qbytes_0_T_1 ? phv_data_21 : _GEN_1564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1566 = 8'h16 == _match_key_qbytes_0_T_1 ? phv_data_22 : _GEN_1565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1567 = 8'h17 == _match_key_qbytes_0_T_1 ? phv_data_23 : _GEN_1566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1568 = 8'h18 == _match_key_qbytes_0_T_1 ? phv_data_24 : _GEN_1567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1569 = 8'h19 == _match_key_qbytes_0_T_1 ? phv_data_25 : _GEN_1568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1570 = 8'h1a == _match_key_qbytes_0_T_1 ? phv_data_26 : _GEN_1569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1571 = 8'h1b == _match_key_qbytes_0_T_1 ? phv_data_27 : _GEN_1570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1572 = 8'h1c == _match_key_qbytes_0_T_1 ? phv_data_28 : _GEN_1571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1573 = 8'h1d == _match_key_qbytes_0_T_1 ? phv_data_29 : _GEN_1572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1574 = 8'h1e == _match_key_qbytes_0_T_1 ? phv_data_30 : _GEN_1573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1575 = 8'h1f == _match_key_qbytes_0_T_1 ? phv_data_31 : _GEN_1574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1576 = 8'h20 == _match_key_qbytes_0_T_1 ? phv_data_32 : _GEN_1575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1577 = 8'h21 == _match_key_qbytes_0_T_1 ? phv_data_33 : _GEN_1576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1578 = 8'h22 == _match_key_qbytes_0_T_1 ? phv_data_34 : _GEN_1577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1579 = 8'h23 == _match_key_qbytes_0_T_1 ? phv_data_35 : _GEN_1578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1580 = 8'h24 == _match_key_qbytes_0_T_1 ? phv_data_36 : _GEN_1579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1581 = 8'h25 == _match_key_qbytes_0_T_1 ? phv_data_37 : _GEN_1580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1582 = 8'h26 == _match_key_qbytes_0_T_1 ? phv_data_38 : _GEN_1581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1583 = 8'h27 == _match_key_qbytes_0_T_1 ? phv_data_39 : _GEN_1582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1584 = 8'h28 == _match_key_qbytes_0_T_1 ? phv_data_40 : _GEN_1583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1585 = 8'h29 == _match_key_qbytes_0_T_1 ? phv_data_41 : _GEN_1584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1586 = 8'h2a == _match_key_qbytes_0_T_1 ? phv_data_42 : _GEN_1585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1587 = 8'h2b == _match_key_qbytes_0_T_1 ? phv_data_43 : _GEN_1586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1588 = 8'h2c == _match_key_qbytes_0_T_1 ? phv_data_44 : _GEN_1587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1589 = 8'h2d == _match_key_qbytes_0_T_1 ? phv_data_45 : _GEN_1588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1590 = 8'h2e == _match_key_qbytes_0_T_1 ? phv_data_46 : _GEN_1589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1591 = 8'h2f == _match_key_qbytes_0_T_1 ? phv_data_47 : _GEN_1590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1592 = 8'h30 == _match_key_qbytes_0_T_1 ? phv_data_48 : _GEN_1591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1593 = 8'h31 == _match_key_qbytes_0_T_1 ? phv_data_49 : _GEN_1592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1594 = 8'h32 == _match_key_qbytes_0_T_1 ? phv_data_50 : _GEN_1593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1595 = 8'h33 == _match_key_qbytes_0_T_1 ? phv_data_51 : _GEN_1594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1596 = 8'h34 == _match_key_qbytes_0_T_1 ? phv_data_52 : _GEN_1595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1597 = 8'h35 == _match_key_qbytes_0_T_1 ? phv_data_53 : _GEN_1596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1598 = 8'h36 == _match_key_qbytes_0_T_1 ? phv_data_54 : _GEN_1597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1599 = 8'h37 == _match_key_qbytes_0_T_1 ? phv_data_55 : _GEN_1598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1600 = 8'h38 == _match_key_qbytes_0_T_1 ? phv_data_56 : _GEN_1599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1601 = 8'h39 == _match_key_qbytes_0_T_1 ? phv_data_57 : _GEN_1600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1602 = 8'h3a == _match_key_qbytes_0_T_1 ? phv_data_58 : _GEN_1601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1603 = 8'h3b == _match_key_qbytes_0_T_1 ? phv_data_59 : _GEN_1602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1604 = 8'h3c == _match_key_qbytes_0_T_1 ? phv_data_60 : _GEN_1603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1605 = 8'h3d == _match_key_qbytes_0_T_1 ? phv_data_61 : _GEN_1604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1606 = 8'h3e == _match_key_qbytes_0_T_1 ? phv_data_62 : _GEN_1605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1607 = 8'h3f == _match_key_qbytes_0_T_1 ? phv_data_63 : _GEN_1606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1608 = 8'h40 == _match_key_qbytes_0_T_1 ? phv_data_64 : _GEN_1607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1609 = 8'h41 == _match_key_qbytes_0_T_1 ? phv_data_65 : _GEN_1608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1610 = 8'h42 == _match_key_qbytes_0_T_1 ? phv_data_66 : _GEN_1609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1611 = 8'h43 == _match_key_qbytes_0_T_1 ? phv_data_67 : _GEN_1610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1612 = 8'h44 == _match_key_qbytes_0_T_1 ? phv_data_68 : _GEN_1611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1613 = 8'h45 == _match_key_qbytes_0_T_1 ? phv_data_69 : _GEN_1612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1614 = 8'h46 == _match_key_qbytes_0_T_1 ? phv_data_70 : _GEN_1613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1615 = 8'h47 == _match_key_qbytes_0_T_1 ? phv_data_71 : _GEN_1614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1616 = 8'h48 == _match_key_qbytes_0_T_1 ? phv_data_72 : _GEN_1615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1617 = 8'h49 == _match_key_qbytes_0_T_1 ? phv_data_73 : _GEN_1616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1618 = 8'h4a == _match_key_qbytes_0_T_1 ? phv_data_74 : _GEN_1617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1619 = 8'h4b == _match_key_qbytes_0_T_1 ? phv_data_75 : _GEN_1618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1620 = 8'h4c == _match_key_qbytes_0_T_1 ? phv_data_76 : _GEN_1619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1621 = 8'h4d == _match_key_qbytes_0_T_1 ? phv_data_77 : _GEN_1620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1622 = 8'h4e == _match_key_qbytes_0_T_1 ? phv_data_78 : _GEN_1621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1623 = 8'h4f == _match_key_qbytes_0_T_1 ? phv_data_79 : _GEN_1622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1624 = 8'h50 == _match_key_qbytes_0_T_1 ? phv_data_80 : _GEN_1623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1625 = 8'h51 == _match_key_qbytes_0_T_1 ? phv_data_81 : _GEN_1624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1626 = 8'h52 == _match_key_qbytes_0_T_1 ? phv_data_82 : _GEN_1625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1627 = 8'h53 == _match_key_qbytes_0_T_1 ? phv_data_83 : _GEN_1626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1628 = 8'h54 == _match_key_qbytes_0_T_1 ? phv_data_84 : _GEN_1627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1629 = 8'h55 == _match_key_qbytes_0_T_1 ? phv_data_85 : _GEN_1628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1630 = 8'h56 == _match_key_qbytes_0_T_1 ? phv_data_86 : _GEN_1629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1631 = 8'h57 == _match_key_qbytes_0_T_1 ? phv_data_87 : _GEN_1630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1632 = 8'h58 == _match_key_qbytes_0_T_1 ? phv_data_88 : _GEN_1631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1633 = 8'h59 == _match_key_qbytes_0_T_1 ? phv_data_89 : _GEN_1632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1634 = 8'h5a == _match_key_qbytes_0_T_1 ? phv_data_90 : _GEN_1633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1635 = 8'h5b == _match_key_qbytes_0_T_1 ? phv_data_91 : _GEN_1634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1636 = 8'h5c == _match_key_qbytes_0_T_1 ? phv_data_92 : _GEN_1635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1637 = 8'h5d == _match_key_qbytes_0_T_1 ? phv_data_93 : _GEN_1636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1638 = 8'h5e == _match_key_qbytes_0_T_1 ? phv_data_94 : _GEN_1637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1639 = 8'h5f == _match_key_qbytes_0_T_1 ? phv_data_95 : _GEN_1638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1640 = 8'h60 == _match_key_qbytes_0_T_1 ? phv_data_96 : _GEN_1639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1641 = 8'h61 == _match_key_qbytes_0_T_1 ? phv_data_97 : _GEN_1640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1642 = 8'h62 == _match_key_qbytes_0_T_1 ? phv_data_98 : _GEN_1641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1643 = 8'h63 == _match_key_qbytes_0_T_1 ? phv_data_99 : _GEN_1642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1644 = 8'h64 == _match_key_qbytes_0_T_1 ? phv_data_100 : _GEN_1643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1645 = 8'h65 == _match_key_qbytes_0_T_1 ? phv_data_101 : _GEN_1644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1646 = 8'h66 == _match_key_qbytes_0_T_1 ? phv_data_102 : _GEN_1645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1647 = 8'h67 == _match_key_qbytes_0_T_1 ? phv_data_103 : _GEN_1646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1648 = 8'h68 == _match_key_qbytes_0_T_1 ? phv_data_104 : _GEN_1647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1649 = 8'h69 == _match_key_qbytes_0_T_1 ? phv_data_105 : _GEN_1648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1650 = 8'h6a == _match_key_qbytes_0_T_1 ? phv_data_106 : _GEN_1649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1651 = 8'h6b == _match_key_qbytes_0_T_1 ? phv_data_107 : _GEN_1650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1652 = 8'h6c == _match_key_qbytes_0_T_1 ? phv_data_108 : _GEN_1651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1653 = 8'h6d == _match_key_qbytes_0_T_1 ? phv_data_109 : _GEN_1652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1654 = 8'h6e == _match_key_qbytes_0_T_1 ? phv_data_110 : _GEN_1653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1655 = 8'h6f == _match_key_qbytes_0_T_1 ? phv_data_111 : _GEN_1654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1656 = 8'h70 == _match_key_qbytes_0_T_1 ? phv_data_112 : _GEN_1655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1657 = 8'h71 == _match_key_qbytes_0_T_1 ? phv_data_113 : _GEN_1656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1658 = 8'h72 == _match_key_qbytes_0_T_1 ? phv_data_114 : _GEN_1657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1659 = 8'h73 == _match_key_qbytes_0_T_1 ? phv_data_115 : _GEN_1658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1660 = 8'h74 == _match_key_qbytes_0_T_1 ? phv_data_116 : _GEN_1659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1661 = 8'h75 == _match_key_qbytes_0_T_1 ? phv_data_117 : _GEN_1660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1662 = 8'h76 == _match_key_qbytes_0_T_1 ? phv_data_118 : _GEN_1661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1663 = 8'h77 == _match_key_qbytes_0_T_1 ? phv_data_119 : _GEN_1662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1664 = 8'h78 == _match_key_qbytes_0_T_1 ? phv_data_120 : _GEN_1663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1665 = 8'h79 == _match_key_qbytes_0_T_1 ? phv_data_121 : _GEN_1664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1666 = 8'h7a == _match_key_qbytes_0_T_1 ? phv_data_122 : _GEN_1665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1667 = 8'h7b == _match_key_qbytes_0_T_1 ? phv_data_123 : _GEN_1666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1668 = 8'h7c == _match_key_qbytes_0_T_1 ? phv_data_124 : _GEN_1667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1669 = 8'h7d == _match_key_qbytes_0_T_1 ? phv_data_125 : _GEN_1668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1670 = 8'h7e == _match_key_qbytes_0_T_1 ? phv_data_126 : _GEN_1669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1671 = 8'h7f == _match_key_qbytes_0_T_1 ? phv_data_127 : _GEN_1670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1672 = 8'h80 == _match_key_qbytes_0_T_1 ? phv_data_128 : _GEN_1671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1673 = 8'h81 == _match_key_qbytes_0_T_1 ? phv_data_129 : _GEN_1672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1674 = 8'h82 == _match_key_qbytes_0_T_1 ? phv_data_130 : _GEN_1673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1675 = 8'h83 == _match_key_qbytes_0_T_1 ? phv_data_131 : _GEN_1674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1676 = 8'h84 == _match_key_qbytes_0_T_1 ? phv_data_132 : _GEN_1675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1677 = 8'h85 == _match_key_qbytes_0_T_1 ? phv_data_133 : _GEN_1676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1678 = 8'h86 == _match_key_qbytes_0_T_1 ? phv_data_134 : _GEN_1677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1679 = 8'h87 == _match_key_qbytes_0_T_1 ? phv_data_135 : _GEN_1678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1680 = 8'h88 == _match_key_qbytes_0_T_1 ? phv_data_136 : _GEN_1679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1681 = 8'h89 == _match_key_qbytes_0_T_1 ? phv_data_137 : _GEN_1680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1682 = 8'h8a == _match_key_qbytes_0_T_1 ? phv_data_138 : _GEN_1681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1683 = 8'h8b == _match_key_qbytes_0_T_1 ? phv_data_139 : _GEN_1682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1684 = 8'h8c == _match_key_qbytes_0_T_1 ? phv_data_140 : _GEN_1683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1685 = 8'h8d == _match_key_qbytes_0_T_1 ? phv_data_141 : _GEN_1684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1686 = 8'h8e == _match_key_qbytes_0_T_1 ? phv_data_142 : _GEN_1685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1687 = 8'h8f == _match_key_qbytes_0_T_1 ? phv_data_143 : _GEN_1686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1688 = 8'h90 == _match_key_qbytes_0_T_1 ? phv_data_144 : _GEN_1687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1689 = 8'h91 == _match_key_qbytes_0_T_1 ? phv_data_145 : _GEN_1688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1690 = 8'h92 == _match_key_qbytes_0_T_1 ? phv_data_146 : _GEN_1689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1691 = 8'h93 == _match_key_qbytes_0_T_1 ? phv_data_147 : _GEN_1690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1692 = 8'h94 == _match_key_qbytes_0_T_1 ? phv_data_148 : _GEN_1691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1693 = 8'h95 == _match_key_qbytes_0_T_1 ? phv_data_149 : _GEN_1692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1694 = 8'h96 == _match_key_qbytes_0_T_1 ? phv_data_150 : _GEN_1693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1695 = 8'h97 == _match_key_qbytes_0_T_1 ? phv_data_151 : _GEN_1694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1696 = 8'h98 == _match_key_qbytes_0_T_1 ? phv_data_152 : _GEN_1695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1697 = 8'h99 == _match_key_qbytes_0_T_1 ? phv_data_153 : _GEN_1696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1698 = 8'h9a == _match_key_qbytes_0_T_1 ? phv_data_154 : _GEN_1697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1699 = 8'h9b == _match_key_qbytes_0_T_1 ? phv_data_155 : _GEN_1698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1700 = 8'h9c == _match_key_qbytes_0_T_1 ? phv_data_156 : _GEN_1699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1701 = 8'h9d == _match_key_qbytes_0_T_1 ? phv_data_157 : _GEN_1700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1702 = 8'h9e == _match_key_qbytes_0_T_1 ? phv_data_158 : _GEN_1701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1703 = 8'h9f == _match_key_qbytes_0_T_1 ? phv_data_159 : _GEN_1702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1704 = 8'ha0 == _match_key_qbytes_0_T_1 ? phv_data_160 : _GEN_1703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1705 = 8'ha1 == _match_key_qbytes_0_T_1 ? phv_data_161 : _GEN_1704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1706 = 8'ha2 == _match_key_qbytes_0_T_1 ? phv_data_162 : _GEN_1705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1707 = 8'ha3 == _match_key_qbytes_0_T_1 ? phv_data_163 : _GEN_1706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1708 = 8'ha4 == _match_key_qbytes_0_T_1 ? phv_data_164 : _GEN_1707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1709 = 8'ha5 == _match_key_qbytes_0_T_1 ? phv_data_165 : _GEN_1708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1710 = 8'ha6 == _match_key_qbytes_0_T_1 ? phv_data_166 : _GEN_1709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1711 = 8'ha7 == _match_key_qbytes_0_T_1 ? phv_data_167 : _GEN_1710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1712 = 8'ha8 == _match_key_qbytes_0_T_1 ? phv_data_168 : _GEN_1711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1713 = 8'ha9 == _match_key_qbytes_0_T_1 ? phv_data_169 : _GEN_1712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1714 = 8'haa == _match_key_qbytes_0_T_1 ? phv_data_170 : _GEN_1713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1715 = 8'hab == _match_key_qbytes_0_T_1 ? phv_data_171 : _GEN_1714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1716 = 8'hac == _match_key_qbytes_0_T_1 ? phv_data_172 : _GEN_1715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1717 = 8'had == _match_key_qbytes_0_T_1 ? phv_data_173 : _GEN_1716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1718 = 8'hae == _match_key_qbytes_0_T_1 ? phv_data_174 : _GEN_1717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1719 = 8'haf == _match_key_qbytes_0_T_1 ? phv_data_175 : _GEN_1718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1720 = 8'hb0 == _match_key_qbytes_0_T_1 ? phv_data_176 : _GEN_1719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1721 = 8'hb1 == _match_key_qbytes_0_T_1 ? phv_data_177 : _GEN_1720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1722 = 8'hb2 == _match_key_qbytes_0_T_1 ? phv_data_178 : _GEN_1721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1723 = 8'hb3 == _match_key_qbytes_0_T_1 ? phv_data_179 : _GEN_1722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1724 = 8'hb4 == _match_key_qbytes_0_T_1 ? phv_data_180 : _GEN_1723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1725 = 8'hb5 == _match_key_qbytes_0_T_1 ? phv_data_181 : _GEN_1724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1726 = 8'hb6 == _match_key_qbytes_0_T_1 ? phv_data_182 : _GEN_1725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1727 = 8'hb7 == _match_key_qbytes_0_T_1 ? phv_data_183 : _GEN_1726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1728 = 8'hb8 == _match_key_qbytes_0_T_1 ? phv_data_184 : _GEN_1727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1729 = 8'hb9 == _match_key_qbytes_0_T_1 ? phv_data_185 : _GEN_1728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1730 = 8'hba == _match_key_qbytes_0_T_1 ? phv_data_186 : _GEN_1729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1731 = 8'hbb == _match_key_qbytes_0_T_1 ? phv_data_187 : _GEN_1730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1732 = 8'hbc == _match_key_qbytes_0_T_1 ? phv_data_188 : _GEN_1731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1733 = 8'hbd == _match_key_qbytes_0_T_1 ? phv_data_189 : _GEN_1732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1734 = 8'hbe == _match_key_qbytes_0_T_1 ? phv_data_190 : _GEN_1733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1735 = 8'hbf == _match_key_qbytes_0_T_1 ? phv_data_191 : _GEN_1734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1736 = 8'hc0 == _match_key_qbytes_0_T_1 ? phv_data_192 : _GEN_1735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1737 = 8'hc1 == _match_key_qbytes_0_T_1 ? phv_data_193 : _GEN_1736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1738 = 8'hc2 == _match_key_qbytes_0_T_1 ? phv_data_194 : _GEN_1737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1739 = 8'hc3 == _match_key_qbytes_0_T_1 ? phv_data_195 : _GEN_1738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1740 = 8'hc4 == _match_key_qbytes_0_T_1 ? phv_data_196 : _GEN_1739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1741 = 8'hc5 == _match_key_qbytes_0_T_1 ? phv_data_197 : _GEN_1740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1742 = 8'hc6 == _match_key_qbytes_0_T_1 ? phv_data_198 : _GEN_1741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1743 = 8'hc7 == _match_key_qbytes_0_T_1 ? phv_data_199 : _GEN_1742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1744 = 8'hc8 == _match_key_qbytes_0_T_1 ? phv_data_200 : _GEN_1743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1745 = 8'hc9 == _match_key_qbytes_0_T_1 ? phv_data_201 : _GEN_1744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1746 = 8'hca == _match_key_qbytes_0_T_1 ? phv_data_202 : _GEN_1745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1747 = 8'hcb == _match_key_qbytes_0_T_1 ? phv_data_203 : _GEN_1746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1748 = 8'hcc == _match_key_qbytes_0_T_1 ? phv_data_204 : _GEN_1747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1749 = 8'hcd == _match_key_qbytes_0_T_1 ? phv_data_205 : _GEN_1748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1750 = 8'hce == _match_key_qbytes_0_T_1 ? phv_data_206 : _GEN_1749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1751 = 8'hcf == _match_key_qbytes_0_T_1 ? phv_data_207 : _GEN_1750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1752 = 8'hd0 == _match_key_qbytes_0_T_1 ? phv_data_208 : _GEN_1751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1753 = 8'hd1 == _match_key_qbytes_0_T_1 ? phv_data_209 : _GEN_1752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1754 = 8'hd2 == _match_key_qbytes_0_T_1 ? phv_data_210 : _GEN_1753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1755 = 8'hd3 == _match_key_qbytes_0_T_1 ? phv_data_211 : _GEN_1754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1756 = 8'hd4 == _match_key_qbytes_0_T_1 ? phv_data_212 : _GEN_1755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1757 = 8'hd5 == _match_key_qbytes_0_T_1 ? phv_data_213 : _GEN_1756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1758 = 8'hd6 == _match_key_qbytes_0_T_1 ? phv_data_214 : _GEN_1757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1759 = 8'hd7 == _match_key_qbytes_0_T_1 ? phv_data_215 : _GEN_1758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1760 = 8'hd8 == _match_key_qbytes_0_T_1 ? phv_data_216 : _GEN_1759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1761 = 8'hd9 == _match_key_qbytes_0_T_1 ? phv_data_217 : _GEN_1760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1762 = 8'hda == _match_key_qbytes_0_T_1 ? phv_data_218 : _GEN_1761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1763 = 8'hdb == _match_key_qbytes_0_T_1 ? phv_data_219 : _GEN_1762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1764 = 8'hdc == _match_key_qbytes_0_T_1 ? phv_data_220 : _GEN_1763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1765 = 8'hdd == _match_key_qbytes_0_T_1 ? phv_data_221 : _GEN_1764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1766 = 8'hde == _match_key_qbytes_0_T_1 ? phv_data_222 : _GEN_1765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1767 = 8'hdf == _match_key_qbytes_0_T_1 ? phv_data_223 : _GEN_1766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1768 = 8'he0 == _match_key_qbytes_0_T_1 ? phv_data_224 : _GEN_1767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1769 = 8'he1 == _match_key_qbytes_0_T_1 ? phv_data_225 : _GEN_1768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1770 = 8'he2 == _match_key_qbytes_0_T_1 ? phv_data_226 : _GEN_1769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1771 = 8'he3 == _match_key_qbytes_0_T_1 ? phv_data_227 : _GEN_1770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1772 = 8'he4 == _match_key_qbytes_0_T_1 ? phv_data_228 : _GEN_1771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1773 = 8'he5 == _match_key_qbytes_0_T_1 ? phv_data_229 : _GEN_1772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1774 = 8'he6 == _match_key_qbytes_0_T_1 ? phv_data_230 : _GEN_1773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1775 = 8'he7 == _match_key_qbytes_0_T_1 ? phv_data_231 : _GEN_1774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1776 = 8'he8 == _match_key_qbytes_0_T_1 ? phv_data_232 : _GEN_1775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1777 = 8'he9 == _match_key_qbytes_0_T_1 ? phv_data_233 : _GEN_1776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1778 = 8'hea == _match_key_qbytes_0_T_1 ? phv_data_234 : _GEN_1777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1779 = 8'heb == _match_key_qbytes_0_T_1 ? phv_data_235 : _GEN_1778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1780 = 8'hec == _match_key_qbytes_0_T_1 ? phv_data_236 : _GEN_1779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1781 = 8'hed == _match_key_qbytes_0_T_1 ? phv_data_237 : _GEN_1780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1782 = 8'hee == _match_key_qbytes_0_T_1 ? phv_data_238 : _GEN_1781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1783 = 8'hef == _match_key_qbytes_0_T_1 ? phv_data_239 : _GEN_1782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1784 = 8'hf0 == _match_key_qbytes_0_T_1 ? phv_data_240 : _GEN_1783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1785 = 8'hf1 == _match_key_qbytes_0_T_1 ? phv_data_241 : _GEN_1784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1786 = 8'hf2 == _match_key_qbytes_0_T_1 ? phv_data_242 : _GEN_1785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1787 = 8'hf3 == _match_key_qbytes_0_T_1 ? phv_data_243 : _GEN_1786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1788 = 8'hf4 == _match_key_qbytes_0_T_1 ? phv_data_244 : _GEN_1787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1789 = 8'hf5 == _match_key_qbytes_0_T_1 ? phv_data_245 : _GEN_1788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1790 = 8'hf6 == _match_key_qbytes_0_T_1 ? phv_data_246 : _GEN_1789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1791 = 8'hf7 == _match_key_qbytes_0_T_1 ? phv_data_247 : _GEN_1790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1792 = 8'hf8 == _match_key_qbytes_0_T_1 ? phv_data_248 : _GEN_1791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1793 = 8'hf9 == _match_key_qbytes_0_T_1 ? phv_data_249 : _GEN_1792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1794 = 8'hfa == _match_key_qbytes_0_T_1 ? phv_data_250 : _GEN_1793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1795 = 8'hfb == _match_key_qbytes_0_T_1 ? phv_data_251 : _GEN_1794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1796 = 8'hfc == _match_key_qbytes_0_T_1 ? phv_data_252 : _GEN_1795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1797 = 8'hfd == _match_key_qbytes_0_T_1 ? phv_data_253 : _GEN_1796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1798 = 8'hfe == _match_key_qbytes_0_T_1 ? phv_data_254 : _GEN_1797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1799 = 8'hff == _match_key_qbytes_0_T_1 ? phv_data_255 : _GEN_1798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_13094 = {{1'd0}, _match_key_qbytes_0_T_1}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1800 = 9'h100 == _GEN_13094 ? phv_data_256 : _GEN_1799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1801 = 9'h101 == _GEN_13094 ? phv_data_257 : _GEN_1800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1802 = 9'h102 == _GEN_13094 ? phv_data_258 : _GEN_1801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1803 = 9'h103 == _GEN_13094 ? phv_data_259 : _GEN_1802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1804 = 9'h104 == _GEN_13094 ? phv_data_260 : _GEN_1803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1805 = 9'h105 == _GEN_13094 ? phv_data_261 : _GEN_1804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1806 = 9'h106 == _GEN_13094 ? phv_data_262 : _GEN_1805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1807 = 9'h107 == _GEN_13094 ? phv_data_263 : _GEN_1806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1808 = 9'h108 == _GEN_13094 ? phv_data_264 : _GEN_1807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1809 = 9'h109 == _GEN_13094 ? phv_data_265 : _GEN_1808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1810 = 9'h10a == _GEN_13094 ? phv_data_266 : _GEN_1809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1811 = 9'h10b == _GEN_13094 ? phv_data_267 : _GEN_1810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1812 = 9'h10c == _GEN_13094 ? phv_data_268 : _GEN_1811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1813 = 9'h10d == _GEN_13094 ? phv_data_269 : _GEN_1812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1814 = 9'h10e == _GEN_13094 ? phv_data_270 : _GEN_1813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1815 = 9'h10f == _GEN_13094 ? phv_data_271 : _GEN_1814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1816 = 9'h110 == _GEN_13094 ? phv_data_272 : _GEN_1815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1817 = 9'h111 == _GEN_13094 ? phv_data_273 : _GEN_1816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1818 = 9'h112 == _GEN_13094 ? phv_data_274 : _GEN_1817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1819 = 9'h113 == _GEN_13094 ? phv_data_275 : _GEN_1818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1820 = 9'h114 == _GEN_13094 ? phv_data_276 : _GEN_1819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1821 = 9'h115 == _GEN_13094 ? phv_data_277 : _GEN_1820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1822 = 9'h116 == _GEN_13094 ? phv_data_278 : _GEN_1821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1823 = 9'h117 == _GEN_13094 ? phv_data_279 : _GEN_1822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1824 = 9'h118 == _GEN_13094 ? phv_data_280 : _GEN_1823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1825 = 9'h119 == _GEN_13094 ? phv_data_281 : _GEN_1824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1826 = 9'h11a == _GEN_13094 ? phv_data_282 : _GEN_1825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1827 = 9'h11b == _GEN_13094 ? phv_data_283 : _GEN_1826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1828 = 9'h11c == _GEN_13094 ? phv_data_284 : _GEN_1827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1829 = 9'h11d == _GEN_13094 ? phv_data_285 : _GEN_1828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1830 = 9'h11e == _GEN_13094 ? phv_data_286 : _GEN_1829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1831 = 9'h11f == _GEN_13094 ? phv_data_287 : _GEN_1830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1832 = 9'h120 == _GEN_13094 ? phv_data_288 : _GEN_1831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1833 = 9'h121 == _GEN_13094 ? phv_data_289 : _GEN_1832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1834 = 9'h122 == _GEN_13094 ? phv_data_290 : _GEN_1833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1835 = 9'h123 == _GEN_13094 ? phv_data_291 : _GEN_1834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1836 = 9'h124 == _GEN_13094 ? phv_data_292 : _GEN_1835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1837 = 9'h125 == _GEN_13094 ? phv_data_293 : _GEN_1836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1838 = 9'h126 == _GEN_13094 ? phv_data_294 : _GEN_1837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1839 = 9'h127 == _GEN_13094 ? phv_data_295 : _GEN_1838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1840 = 9'h128 == _GEN_13094 ? phv_data_296 : _GEN_1839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1841 = 9'h129 == _GEN_13094 ? phv_data_297 : _GEN_1840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1842 = 9'h12a == _GEN_13094 ? phv_data_298 : _GEN_1841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1843 = 9'h12b == _GEN_13094 ? phv_data_299 : _GEN_1842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1844 = 9'h12c == _GEN_13094 ? phv_data_300 : _GEN_1843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1845 = 9'h12d == _GEN_13094 ? phv_data_301 : _GEN_1844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1846 = 9'h12e == _GEN_13094 ? phv_data_302 : _GEN_1845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1847 = 9'h12f == _GEN_13094 ? phv_data_303 : _GEN_1846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1848 = 9'h130 == _GEN_13094 ? phv_data_304 : _GEN_1847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1849 = 9'h131 == _GEN_13094 ? phv_data_305 : _GEN_1848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1850 = 9'h132 == _GEN_13094 ? phv_data_306 : _GEN_1849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1851 = 9'h133 == _GEN_13094 ? phv_data_307 : _GEN_1850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1852 = 9'h134 == _GEN_13094 ? phv_data_308 : _GEN_1851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1853 = 9'h135 == _GEN_13094 ? phv_data_309 : _GEN_1852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1854 = 9'h136 == _GEN_13094 ? phv_data_310 : _GEN_1853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1855 = 9'h137 == _GEN_13094 ? phv_data_311 : _GEN_1854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1856 = 9'h138 == _GEN_13094 ? phv_data_312 : _GEN_1855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1857 = 9'h139 == _GEN_13094 ? phv_data_313 : _GEN_1856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1858 = 9'h13a == _GEN_13094 ? phv_data_314 : _GEN_1857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1859 = 9'h13b == _GEN_13094 ? phv_data_315 : _GEN_1858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1860 = 9'h13c == _GEN_13094 ? phv_data_316 : _GEN_1859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1861 = 9'h13d == _GEN_13094 ? phv_data_317 : _GEN_1860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1862 = 9'h13e == _GEN_13094 ? phv_data_318 : _GEN_1861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1863 = 9'h13f == _GEN_13094 ? phv_data_319 : _GEN_1862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1864 = 9'h140 == _GEN_13094 ? phv_data_320 : _GEN_1863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1865 = 9'h141 == _GEN_13094 ? phv_data_321 : _GEN_1864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1866 = 9'h142 == _GEN_13094 ? phv_data_322 : _GEN_1865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1867 = 9'h143 == _GEN_13094 ? phv_data_323 : _GEN_1866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1868 = 9'h144 == _GEN_13094 ? phv_data_324 : _GEN_1867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1869 = 9'h145 == _GEN_13094 ? phv_data_325 : _GEN_1868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1870 = 9'h146 == _GEN_13094 ? phv_data_326 : _GEN_1869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1871 = 9'h147 == _GEN_13094 ? phv_data_327 : _GEN_1870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1872 = 9'h148 == _GEN_13094 ? phv_data_328 : _GEN_1871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1873 = 9'h149 == _GEN_13094 ? phv_data_329 : _GEN_1872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1874 = 9'h14a == _GEN_13094 ? phv_data_330 : _GEN_1873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1875 = 9'h14b == _GEN_13094 ? phv_data_331 : _GEN_1874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1876 = 9'h14c == _GEN_13094 ? phv_data_332 : _GEN_1875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1877 = 9'h14d == _GEN_13094 ? phv_data_333 : _GEN_1876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1878 = 9'h14e == _GEN_13094 ? phv_data_334 : _GEN_1877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1879 = 9'h14f == _GEN_13094 ? phv_data_335 : _GEN_1878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1880 = 9'h150 == _GEN_13094 ? phv_data_336 : _GEN_1879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1881 = 9'h151 == _GEN_13094 ? phv_data_337 : _GEN_1880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1882 = 9'h152 == _GEN_13094 ? phv_data_338 : _GEN_1881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1883 = 9'h153 == _GEN_13094 ? phv_data_339 : _GEN_1882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1884 = 9'h154 == _GEN_13094 ? phv_data_340 : _GEN_1883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1885 = 9'h155 == _GEN_13094 ? phv_data_341 : _GEN_1884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1886 = 9'h156 == _GEN_13094 ? phv_data_342 : _GEN_1885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1887 = 9'h157 == _GEN_13094 ? phv_data_343 : _GEN_1886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1888 = 9'h158 == _GEN_13094 ? phv_data_344 : _GEN_1887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1889 = 9'h159 == _GEN_13094 ? phv_data_345 : _GEN_1888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1890 = 9'h15a == _GEN_13094 ? phv_data_346 : _GEN_1889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1891 = 9'h15b == _GEN_13094 ? phv_data_347 : _GEN_1890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1892 = 9'h15c == _GEN_13094 ? phv_data_348 : _GEN_1891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1893 = 9'h15d == _GEN_13094 ? phv_data_349 : _GEN_1892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1894 = 9'h15e == _GEN_13094 ? phv_data_350 : _GEN_1893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1895 = 9'h15f == _GEN_13094 ? phv_data_351 : _GEN_1894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1896 = 9'h160 == _GEN_13094 ? phv_data_352 : _GEN_1895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1897 = 9'h161 == _GEN_13094 ? phv_data_353 : _GEN_1896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1898 = 9'h162 == _GEN_13094 ? phv_data_354 : _GEN_1897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1899 = 9'h163 == _GEN_13094 ? phv_data_355 : _GEN_1898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1900 = 9'h164 == _GEN_13094 ? phv_data_356 : _GEN_1899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1901 = 9'h165 == _GEN_13094 ? phv_data_357 : _GEN_1900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1902 = 9'h166 == _GEN_13094 ? phv_data_358 : _GEN_1901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1903 = 9'h167 == _GEN_13094 ? phv_data_359 : _GEN_1902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1904 = 9'h168 == _GEN_13094 ? phv_data_360 : _GEN_1903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1905 = 9'h169 == _GEN_13094 ? phv_data_361 : _GEN_1904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1906 = 9'h16a == _GEN_13094 ? phv_data_362 : _GEN_1905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1907 = 9'h16b == _GEN_13094 ? phv_data_363 : _GEN_1906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1908 = 9'h16c == _GEN_13094 ? phv_data_364 : _GEN_1907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1909 = 9'h16d == _GEN_13094 ? phv_data_365 : _GEN_1908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1910 = 9'h16e == _GEN_13094 ? phv_data_366 : _GEN_1909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1911 = 9'h16f == _GEN_13094 ? phv_data_367 : _GEN_1910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1912 = 9'h170 == _GEN_13094 ? phv_data_368 : _GEN_1911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1913 = 9'h171 == _GEN_13094 ? phv_data_369 : _GEN_1912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1914 = 9'h172 == _GEN_13094 ? phv_data_370 : _GEN_1913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1915 = 9'h173 == _GEN_13094 ? phv_data_371 : _GEN_1914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1916 = 9'h174 == _GEN_13094 ? phv_data_372 : _GEN_1915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1917 = 9'h175 == _GEN_13094 ? phv_data_373 : _GEN_1916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1918 = 9'h176 == _GEN_13094 ? phv_data_374 : _GEN_1917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1919 = 9'h177 == _GEN_13094 ? phv_data_375 : _GEN_1918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1920 = 9'h178 == _GEN_13094 ? phv_data_376 : _GEN_1919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1921 = 9'h179 == _GEN_13094 ? phv_data_377 : _GEN_1920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1922 = 9'h17a == _GEN_13094 ? phv_data_378 : _GEN_1921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1923 = 9'h17b == _GEN_13094 ? phv_data_379 : _GEN_1922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1924 = 9'h17c == _GEN_13094 ? phv_data_380 : _GEN_1923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1925 = 9'h17d == _GEN_13094 ? phv_data_381 : _GEN_1924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1926 = 9'h17e == _GEN_13094 ? phv_data_382 : _GEN_1925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1927 = 9'h17f == _GEN_13094 ? phv_data_383 : _GEN_1926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1928 = 9'h180 == _GEN_13094 ? phv_data_384 : _GEN_1927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1929 = 9'h181 == _GEN_13094 ? phv_data_385 : _GEN_1928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1930 = 9'h182 == _GEN_13094 ? phv_data_386 : _GEN_1929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1931 = 9'h183 == _GEN_13094 ? phv_data_387 : _GEN_1930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1932 = 9'h184 == _GEN_13094 ? phv_data_388 : _GEN_1931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1933 = 9'h185 == _GEN_13094 ? phv_data_389 : _GEN_1932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1934 = 9'h186 == _GEN_13094 ? phv_data_390 : _GEN_1933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1935 = 9'h187 == _GEN_13094 ? phv_data_391 : _GEN_1934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1936 = 9'h188 == _GEN_13094 ? phv_data_392 : _GEN_1935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1937 = 9'h189 == _GEN_13094 ? phv_data_393 : _GEN_1936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1938 = 9'h18a == _GEN_13094 ? phv_data_394 : _GEN_1937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1939 = 9'h18b == _GEN_13094 ? phv_data_395 : _GEN_1938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1940 = 9'h18c == _GEN_13094 ? phv_data_396 : _GEN_1939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1941 = 9'h18d == _GEN_13094 ? phv_data_397 : _GEN_1940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1942 = 9'h18e == _GEN_13094 ? phv_data_398 : _GEN_1941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1943 = 9'h18f == _GEN_13094 ? phv_data_399 : _GEN_1942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1944 = 9'h190 == _GEN_13094 ? phv_data_400 : _GEN_1943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1945 = 9'h191 == _GEN_13094 ? phv_data_401 : _GEN_1944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1946 = 9'h192 == _GEN_13094 ? phv_data_402 : _GEN_1945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1947 = 9'h193 == _GEN_13094 ? phv_data_403 : _GEN_1946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1948 = 9'h194 == _GEN_13094 ? phv_data_404 : _GEN_1947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1949 = 9'h195 == _GEN_13094 ? phv_data_405 : _GEN_1948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1950 = 9'h196 == _GEN_13094 ? phv_data_406 : _GEN_1949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1951 = 9'h197 == _GEN_13094 ? phv_data_407 : _GEN_1950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1952 = 9'h198 == _GEN_13094 ? phv_data_408 : _GEN_1951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1953 = 9'h199 == _GEN_13094 ? phv_data_409 : _GEN_1952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1954 = 9'h19a == _GEN_13094 ? phv_data_410 : _GEN_1953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1955 = 9'h19b == _GEN_13094 ? phv_data_411 : _GEN_1954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1956 = 9'h19c == _GEN_13094 ? phv_data_412 : _GEN_1955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1957 = 9'h19d == _GEN_13094 ? phv_data_413 : _GEN_1956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1958 = 9'h19e == _GEN_13094 ? phv_data_414 : _GEN_1957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1959 = 9'h19f == _GEN_13094 ? phv_data_415 : _GEN_1958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1960 = 9'h1a0 == _GEN_13094 ? phv_data_416 : _GEN_1959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1961 = 9'h1a1 == _GEN_13094 ? phv_data_417 : _GEN_1960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1962 = 9'h1a2 == _GEN_13094 ? phv_data_418 : _GEN_1961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1963 = 9'h1a3 == _GEN_13094 ? phv_data_419 : _GEN_1962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1964 = 9'h1a4 == _GEN_13094 ? phv_data_420 : _GEN_1963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1965 = 9'h1a5 == _GEN_13094 ? phv_data_421 : _GEN_1964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1966 = 9'h1a6 == _GEN_13094 ? phv_data_422 : _GEN_1965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1967 = 9'h1a7 == _GEN_13094 ? phv_data_423 : _GEN_1966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1968 = 9'h1a8 == _GEN_13094 ? phv_data_424 : _GEN_1967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1969 = 9'h1a9 == _GEN_13094 ? phv_data_425 : _GEN_1968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1970 = 9'h1aa == _GEN_13094 ? phv_data_426 : _GEN_1969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1971 = 9'h1ab == _GEN_13094 ? phv_data_427 : _GEN_1970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1972 = 9'h1ac == _GEN_13094 ? phv_data_428 : _GEN_1971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1973 = 9'h1ad == _GEN_13094 ? phv_data_429 : _GEN_1972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1974 = 9'h1ae == _GEN_13094 ? phv_data_430 : _GEN_1973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1975 = 9'h1af == _GEN_13094 ? phv_data_431 : _GEN_1974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1976 = 9'h1b0 == _GEN_13094 ? phv_data_432 : _GEN_1975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1977 = 9'h1b1 == _GEN_13094 ? phv_data_433 : _GEN_1976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1978 = 9'h1b2 == _GEN_13094 ? phv_data_434 : _GEN_1977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1979 = 9'h1b3 == _GEN_13094 ? phv_data_435 : _GEN_1978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1980 = 9'h1b4 == _GEN_13094 ? phv_data_436 : _GEN_1979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1981 = 9'h1b5 == _GEN_13094 ? phv_data_437 : _GEN_1980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1982 = 9'h1b6 == _GEN_13094 ? phv_data_438 : _GEN_1981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1983 = 9'h1b7 == _GEN_13094 ? phv_data_439 : _GEN_1982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1984 = 9'h1b8 == _GEN_13094 ? phv_data_440 : _GEN_1983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1985 = 9'h1b9 == _GEN_13094 ? phv_data_441 : _GEN_1984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1986 = 9'h1ba == _GEN_13094 ? phv_data_442 : _GEN_1985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1987 = 9'h1bb == _GEN_13094 ? phv_data_443 : _GEN_1986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1988 = 9'h1bc == _GEN_13094 ? phv_data_444 : _GEN_1987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1989 = 9'h1bd == _GEN_13094 ? phv_data_445 : _GEN_1988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1990 = 9'h1be == _GEN_13094 ? phv_data_446 : _GEN_1989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1991 = 9'h1bf == _GEN_13094 ? phv_data_447 : _GEN_1990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1992 = 9'h1c0 == _GEN_13094 ? phv_data_448 : _GEN_1991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1993 = 9'h1c1 == _GEN_13094 ? phv_data_449 : _GEN_1992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1994 = 9'h1c2 == _GEN_13094 ? phv_data_450 : _GEN_1993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1995 = 9'h1c3 == _GEN_13094 ? phv_data_451 : _GEN_1994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1996 = 9'h1c4 == _GEN_13094 ? phv_data_452 : _GEN_1995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1997 = 9'h1c5 == _GEN_13094 ? phv_data_453 : _GEN_1996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1998 = 9'h1c6 == _GEN_13094 ? phv_data_454 : _GEN_1997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_1999 = 9'h1c7 == _GEN_13094 ? phv_data_455 : _GEN_1998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2000 = 9'h1c8 == _GEN_13094 ? phv_data_456 : _GEN_1999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2001 = 9'h1c9 == _GEN_13094 ? phv_data_457 : _GEN_2000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2002 = 9'h1ca == _GEN_13094 ? phv_data_458 : _GEN_2001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2003 = 9'h1cb == _GEN_13094 ? phv_data_459 : _GEN_2002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2004 = 9'h1cc == _GEN_13094 ? phv_data_460 : _GEN_2003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2005 = 9'h1cd == _GEN_13094 ? phv_data_461 : _GEN_2004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2006 = 9'h1ce == _GEN_13094 ? phv_data_462 : _GEN_2005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2007 = 9'h1cf == _GEN_13094 ? phv_data_463 : _GEN_2006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2008 = 9'h1d0 == _GEN_13094 ? phv_data_464 : _GEN_2007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2009 = 9'h1d1 == _GEN_13094 ? phv_data_465 : _GEN_2008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2010 = 9'h1d2 == _GEN_13094 ? phv_data_466 : _GEN_2009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2011 = 9'h1d3 == _GEN_13094 ? phv_data_467 : _GEN_2010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2012 = 9'h1d4 == _GEN_13094 ? phv_data_468 : _GEN_2011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2013 = 9'h1d5 == _GEN_13094 ? phv_data_469 : _GEN_2012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2014 = 9'h1d6 == _GEN_13094 ? phv_data_470 : _GEN_2013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2015 = 9'h1d7 == _GEN_13094 ? phv_data_471 : _GEN_2014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2016 = 9'h1d8 == _GEN_13094 ? phv_data_472 : _GEN_2015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2017 = 9'h1d9 == _GEN_13094 ? phv_data_473 : _GEN_2016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2018 = 9'h1da == _GEN_13094 ? phv_data_474 : _GEN_2017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2019 = 9'h1db == _GEN_13094 ? phv_data_475 : _GEN_2018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2020 = 9'h1dc == _GEN_13094 ? phv_data_476 : _GEN_2019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2021 = 9'h1dd == _GEN_13094 ? phv_data_477 : _GEN_2020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2022 = 9'h1de == _GEN_13094 ? phv_data_478 : _GEN_2021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2023 = 9'h1df == _GEN_13094 ? phv_data_479 : _GEN_2022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2024 = 9'h1e0 == _GEN_13094 ? phv_data_480 : _GEN_2023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2025 = 9'h1e1 == _GEN_13094 ? phv_data_481 : _GEN_2024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2026 = 9'h1e2 == _GEN_13094 ? phv_data_482 : _GEN_2025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2027 = 9'h1e3 == _GEN_13094 ? phv_data_483 : _GEN_2026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2028 = 9'h1e4 == _GEN_13094 ? phv_data_484 : _GEN_2027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2029 = 9'h1e5 == _GEN_13094 ? phv_data_485 : _GEN_2028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2030 = 9'h1e6 == _GEN_13094 ? phv_data_486 : _GEN_2029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2031 = 9'h1e7 == _GEN_13094 ? phv_data_487 : _GEN_2030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2032 = 9'h1e8 == _GEN_13094 ? phv_data_488 : _GEN_2031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2033 = 9'h1e9 == _GEN_13094 ? phv_data_489 : _GEN_2032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2034 = 9'h1ea == _GEN_13094 ? phv_data_490 : _GEN_2033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2035 = 9'h1eb == _GEN_13094 ? phv_data_491 : _GEN_2034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2036 = 9'h1ec == _GEN_13094 ? phv_data_492 : _GEN_2035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2037 = 9'h1ed == _GEN_13094 ? phv_data_493 : _GEN_2036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2038 = 9'h1ee == _GEN_13094 ? phv_data_494 : _GEN_2037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2039 = 9'h1ef == _GEN_13094 ? phv_data_495 : _GEN_2038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2040 = 9'h1f0 == _GEN_13094 ? phv_data_496 : _GEN_2039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2041 = 9'h1f1 == _GEN_13094 ? phv_data_497 : _GEN_2040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2042 = 9'h1f2 == _GEN_13094 ? phv_data_498 : _GEN_2041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2043 = 9'h1f3 == _GEN_13094 ? phv_data_499 : _GEN_2042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2044 = 9'h1f4 == _GEN_13094 ? phv_data_500 : _GEN_2043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2045 = 9'h1f5 == _GEN_13094 ? phv_data_501 : _GEN_2044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2046 = 9'h1f6 == _GEN_13094 ? phv_data_502 : _GEN_2045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2047 = 9'h1f7 == _GEN_13094 ? phv_data_503 : _GEN_2046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2048 = 9'h1f8 == _GEN_13094 ? phv_data_504 : _GEN_2047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2049 = 9'h1f9 == _GEN_13094 ? phv_data_505 : _GEN_2048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2050 = 9'h1fa == _GEN_13094 ? phv_data_506 : _GEN_2049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2051 = 9'h1fb == _GEN_13094 ? phv_data_507 : _GEN_2050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2052 = 9'h1fc == _GEN_13094 ? phv_data_508 : _GEN_2051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2053 = 9'h1fd == _GEN_13094 ? phv_data_509 : _GEN_2052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2054 = 9'h1fe == _GEN_13094 ? phv_data_510 : _GEN_2053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2055 = 9'h1ff == _GEN_13094 ? phv_data_511 : _GEN_2054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_0_T_3 = {_GEN_1543,_GEN_2055,_GEN_519,_GEN_1031}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_0 = local_offset < end_offset ? _match_key_qbytes_0_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_1 = 8'h4 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_1_hi = local_offset_1[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_1_T = {match_key_qbytes_1_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_1_T_1 = {match_key_qbytes_1_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_1_T_2 = {match_key_qbytes_1_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2058 = 8'h1 == _match_key_qbytes_1_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2059 = 8'h2 == _match_key_qbytes_1_T_2 ? phv_data_2 : _GEN_2058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2060 = 8'h3 == _match_key_qbytes_1_T_2 ? phv_data_3 : _GEN_2059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2061 = 8'h4 == _match_key_qbytes_1_T_2 ? phv_data_4 : _GEN_2060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2062 = 8'h5 == _match_key_qbytes_1_T_2 ? phv_data_5 : _GEN_2061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2063 = 8'h6 == _match_key_qbytes_1_T_2 ? phv_data_6 : _GEN_2062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2064 = 8'h7 == _match_key_qbytes_1_T_2 ? phv_data_7 : _GEN_2063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2065 = 8'h8 == _match_key_qbytes_1_T_2 ? phv_data_8 : _GEN_2064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2066 = 8'h9 == _match_key_qbytes_1_T_2 ? phv_data_9 : _GEN_2065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2067 = 8'ha == _match_key_qbytes_1_T_2 ? phv_data_10 : _GEN_2066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2068 = 8'hb == _match_key_qbytes_1_T_2 ? phv_data_11 : _GEN_2067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2069 = 8'hc == _match_key_qbytes_1_T_2 ? phv_data_12 : _GEN_2068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2070 = 8'hd == _match_key_qbytes_1_T_2 ? phv_data_13 : _GEN_2069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2071 = 8'he == _match_key_qbytes_1_T_2 ? phv_data_14 : _GEN_2070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2072 = 8'hf == _match_key_qbytes_1_T_2 ? phv_data_15 : _GEN_2071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2073 = 8'h10 == _match_key_qbytes_1_T_2 ? phv_data_16 : _GEN_2072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2074 = 8'h11 == _match_key_qbytes_1_T_2 ? phv_data_17 : _GEN_2073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2075 = 8'h12 == _match_key_qbytes_1_T_2 ? phv_data_18 : _GEN_2074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2076 = 8'h13 == _match_key_qbytes_1_T_2 ? phv_data_19 : _GEN_2075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2077 = 8'h14 == _match_key_qbytes_1_T_2 ? phv_data_20 : _GEN_2076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2078 = 8'h15 == _match_key_qbytes_1_T_2 ? phv_data_21 : _GEN_2077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2079 = 8'h16 == _match_key_qbytes_1_T_2 ? phv_data_22 : _GEN_2078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2080 = 8'h17 == _match_key_qbytes_1_T_2 ? phv_data_23 : _GEN_2079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2081 = 8'h18 == _match_key_qbytes_1_T_2 ? phv_data_24 : _GEN_2080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2082 = 8'h19 == _match_key_qbytes_1_T_2 ? phv_data_25 : _GEN_2081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2083 = 8'h1a == _match_key_qbytes_1_T_2 ? phv_data_26 : _GEN_2082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2084 = 8'h1b == _match_key_qbytes_1_T_2 ? phv_data_27 : _GEN_2083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2085 = 8'h1c == _match_key_qbytes_1_T_2 ? phv_data_28 : _GEN_2084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2086 = 8'h1d == _match_key_qbytes_1_T_2 ? phv_data_29 : _GEN_2085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2087 = 8'h1e == _match_key_qbytes_1_T_2 ? phv_data_30 : _GEN_2086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2088 = 8'h1f == _match_key_qbytes_1_T_2 ? phv_data_31 : _GEN_2087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2089 = 8'h20 == _match_key_qbytes_1_T_2 ? phv_data_32 : _GEN_2088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2090 = 8'h21 == _match_key_qbytes_1_T_2 ? phv_data_33 : _GEN_2089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2091 = 8'h22 == _match_key_qbytes_1_T_2 ? phv_data_34 : _GEN_2090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2092 = 8'h23 == _match_key_qbytes_1_T_2 ? phv_data_35 : _GEN_2091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2093 = 8'h24 == _match_key_qbytes_1_T_2 ? phv_data_36 : _GEN_2092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2094 = 8'h25 == _match_key_qbytes_1_T_2 ? phv_data_37 : _GEN_2093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2095 = 8'h26 == _match_key_qbytes_1_T_2 ? phv_data_38 : _GEN_2094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2096 = 8'h27 == _match_key_qbytes_1_T_2 ? phv_data_39 : _GEN_2095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2097 = 8'h28 == _match_key_qbytes_1_T_2 ? phv_data_40 : _GEN_2096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2098 = 8'h29 == _match_key_qbytes_1_T_2 ? phv_data_41 : _GEN_2097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2099 = 8'h2a == _match_key_qbytes_1_T_2 ? phv_data_42 : _GEN_2098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2100 = 8'h2b == _match_key_qbytes_1_T_2 ? phv_data_43 : _GEN_2099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2101 = 8'h2c == _match_key_qbytes_1_T_2 ? phv_data_44 : _GEN_2100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2102 = 8'h2d == _match_key_qbytes_1_T_2 ? phv_data_45 : _GEN_2101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2103 = 8'h2e == _match_key_qbytes_1_T_2 ? phv_data_46 : _GEN_2102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2104 = 8'h2f == _match_key_qbytes_1_T_2 ? phv_data_47 : _GEN_2103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2105 = 8'h30 == _match_key_qbytes_1_T_2 ? phv_data_48 : _GEN_2104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2106 = 8'h31 == _match_key_qbytes_1_T_2 ? phv_data_49 : _GEN_2105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2107 = 8'h32 == _match_key_qbytes_1_T_2 ? phv_data_50 : _GEN_2106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2108 = 8'h33 == _match_key_qbytes_1_T_2 ? phv_data_51 : _GEN_2107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2109 = 8'h34 == _match_key_qbytes_1_T_2 ? phv_data_52 : _GEN_2108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2110 = 8'h35 == _match_key_qbytes_1_T_2 ? phv_data_53 : _GEN_2109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2111 = 8'h36 == _match_key_qbytes_1_T_2 ? phv_data_54 : _GEN_2110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2112 = 8'h37 == _match_key_qbytes_1_T_2 ? phv_data_55 : _GEN_2111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2113 = 8'h38 == _match_key_qbytes_1_T_2 ? phv_data_56 : _GEN_2112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2114 = 8'h39 == _match_key_qbytes_1_T_2 ? phv_data_57 : _GEN_2113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2115 = 8'h3a == _match_key_qbytes_1_T_2 ? phv_data_58 : _GEN_2114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2116 = 8'h3b == _match_key_qbytes_1_T_2 ? phv_data_59 : _GEN_2115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2117 = 8'h3c == _match_key_qbytes_1_T_2 ? phv_data_60 : _GEN_2116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2118 = 8'h3d == _match_key_qbytes_1_T_2 ? phv_data_61 : _GEN_2117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2119 = 8'h3e == _match_key_qbytes_1_T_2 ? phv_data_62 : _GEN_2118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2120 = 8'h3f == _match_key_qbytes_1_T_2 ? phv_data_63 : _GEN_2119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2121 = 8'h40 == _match_key_qbytes_1_T_2 ? phv_data_64 : _GEN_2120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2122 = 8'h41 == _match_key_qbytes_1_T_2 ? phv_data_65 : _GEN_2121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2123 = 8'h42 == _match_key_qbytes_1_T_2 ? phv_data_66 : _GEN_2122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2124 = 8'h43 == _match_key_qbytes_1_T_2 ? phv_data_67 : _GEN_2123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2125 = 8'h44 == _match_key_qbytes_1_T_2 ? phv_data_68 : _GEN_2124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2126 = 8'h45 == _match_key_qbytes_1_T_2 ? phv_data_69 : _GEN_2125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2127 = 8'h46 == _match_key_qbytes_1_T_2 ? phv_data_70 : _GEN_2126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2128 = 8'h47 == _match_key_qbytes_1_T_2 ? phv_data_71 : _GEN_2127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2129 = 8'h48 == _match_key_qbytes_1_T_2 ? phv_data_72 : _GEN_2128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2130 = 8'h49 == _match_key_qbytes_1_T_2 ? phv_data_73 : _GEN_2129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2131 = 8'h4a == _match_key_qbytes_1_T_2 ? phv_data_74 : _GEN_2130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2132 = 8'h4b == _match_key_qbytes_1_T_2 ? phv_data_75 : _GEN_2131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2133 = 8'h4c == _match_key_qbytes_1_T_2 ? phv_data_76 : _GEN_2132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2134 = 8'h4d == _match_key_qbytes_1_T_2 ? phv_data_77 : _GEN_2133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2135 = 8'h4e == _match_key_qbytes_1_T_2 ? phv_data_78 : _GEN_2134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2136 = 8'h4f == _match_key_qbytes_1_T_2 ? phv_data_79 : _GEN_2135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2137 = 8'h50 == _match_key_qbytes_1_T_2 ? phv_data_80 : _GEN_2136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2138 = 8'h51 == _match_key_qbytes_1_T_2 ? phv_data_81 : _GEN_2137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2139 = 8'h52 == _match_key_qbytes_1_T_2 ? phv_data_82 : _GEN_2138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2140 = 8'h53 == _match_key_qbytes_1_T_2 ? phv_data_83 : _GEN_2139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2141 = 8'h54 == _match_key_qbytes_1_T_2 ? phv_data_84 : _GEN_2140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2142 = 8'h55 == _match_key_qbytes_1_T_2 ? phv_data_85 : _GEN_2141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2143 = 8'h56 == _match_key_qbytes_1_T_2 ? phv_data_86 : _GEN_2142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2144 = 8'h57 == _match_key_qbytes_1_T_2 ? phv_data_87 : _GEN_2143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2145 = 8'h58 == _match_key_qbytes_1_T_2 ? phv_data_88 : _GEN_2144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2146 = 8'h59 == _match_key_qbytes_1_T_2 ? phv_data_89 : _GEN_2145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2147 = 8'h5a == _match_key_qbytes_1_T_2 ? phv_data_90 : _GEN_2146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2148 = 8'h5b == _match_key_qbytes_1_T_2 ? phv_data_91 : _GEN_2147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2149 = 8'h5c == _match_key_qbytes_1_T_2 ? phv_data_92 : _GEN_2148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2150 = 8'h5d == _match_key_qbytes_1_T_2 ? phv_data_93 : _GEN_2149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2151 = 8'h5e == _match_key_qbytes_1_T_2 ? phv_data_94 : _GEN_2150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2152 = 8'h5f == _match_key_qbytes_1_T_2 ? phv_data_95 : _GEN_2151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2153 = 8'h60 == _match_key_qbytes_1_T_2 ? phv_data_96 : _GEN_2152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2154 = 8'h61 == _match_key_qbytes_1_T_2 ? phv_data_97 : _GEN_2153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2155 = 8'h62 == _match_key_qbytes_1_T_2 ? phv_data_98 : _GEN_2154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2156 = 8'h63 == _match_key_qbytes_1_T_2 ? phv_data_99 : _GEN_2155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2157 = 8'h64 == _match_key_qbytes_1_T_2 ? phv_data_100 : _GEN_2156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2158 = 8'h65 == _match_key_qbytes_1_T_2 ? phv_data_101 : _GEN_2157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2159 = 8'h66 == _match_key_qbytes_1_T_2 ? phv_data_102 : _GEN_2158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2160 = 8'h67 == _match_key_qbytes_1_T_2 ? phv_data_103 : _GEN_2159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2161 = 8'h68 == _match_key_qbytes_1_T_2 ? phv_data_104 : _GEN_2160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2162 = 8'h69 == _match_key_qbytes_1_T_2 ? phv_data_105 : _GEN_2161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2163 = 8'h6a == _match_key_qbytes_1_T_2 ? phv_data_106 : _GEN_2162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2164 = 8'h6b == _match_key_qbytes_1_T_2 ? phv_data_107 : _GEN_2163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2165 = 8'h6c == _match_key_qbytes_1_T_2 ? phv_data_108 : _GEN_2164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2166 = 8'h6d == _match_key_qbytes_1_T_2 ? phv_data_109 : _GEN_2165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2167 = 8'h6e == _match_key_qbytes_1_T_2 ? phv_data_110 : _GEN_2166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2168 = 8'h6f == _match_key_qbytes_1_T_2 ? phv_data_111 : _GEN_2167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2169 = 8'h70 == _match_key_qbytes_1_T_2 ? phv_data_112 : _GEN_2168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2170 = 8'h71 == _match_key_qbytes_1_T_2 ? phv_data_113 : _GEN_2169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2171 = 8'h72 == _match_key_qbytes_1_T_2 ? phv_data_114 : _GEN_2170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2172 = 8'h73 == _match_key_qbytes_1_T_2 ? phv_data_115 : _GEN_2171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2173 = 8'h74 == _match_key_qbytes_1_T_2 ? phv_data_116 : _GEN_2172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2174 = 8'h75 == _match_key_qbytes_1_T_2 ? phv_data_117 : _GEN_2173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2175 = 8'h76 == _match_key_qbytes_1_T_2 ? phv_data_118 : _GEN_2174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2176 = 8'h77 == _match_key_qbytes_1_T_2 ? phv_data_119 : _GEN_2175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2177 = 8'h78 == _match_key_qbytes_1_T_2 ? phv_data_120 : _GEN_2176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2178 = 8'h79 == _match_key_qbytes_1_T_2 ? phv_data_121 : _GEN_2177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2179 = 8'h7a == _match_key_qbytes_1_T_2 ? phv_data_122 : _GEN_2178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2180 = 8'h7b == _match_key_qbytes_1_T_2 ? phv_data_123 : _GEN_2179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2181 = 8'h7c == _match_key_qbytes_1_T_2 ? phv_data_124 : _GEN_2180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2182 = 8'h7d == _match_key_qbytes_1_T_2 ? phv_data_125 : _GEN_2181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2183 = 8'h7e == _match_key_qbytes_1_T_2 ? phv_data_126 : _GEN_2182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2184 = 8'h7f == _match_key_qbytes_1_T_2 ? phv_data_127 : _GEN_2183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2185 = 8'h80 == _match_key_qbytes_1_T_2 ? phv_data_128 : _GEN_2184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2186 = 8'h81 == _match_key_qbytes_1_T_2 ? phv_data_129 : _GEN_2185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2187 = 8'h82 == _match_key_qbytes_1_T_2 ? phv_data_130 : _GEN_2186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2188 = 8'h83 == _match_key_qbytes_1_T_2 ? phv_data_131 : _GEN_2187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2189 = 8'h84 == _match_key_qbytes_1_T_2 ? phv_data_132 : _GEN_2188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2190 = 8'h85 == _match_key_qbytes_1_T_2 ? phv_data_133 : _GEN_2189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2191 = 8'h86 == _match_key_qbytes_1_T_2 ? phv_data_134 : _GEN_2190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2192 = 8'h87 == _match_key_qbytes_1_T_2 ? phv_data_135 : _GEN_2191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2193 = 8'h88 == _match_key_qbytes_1_T_2 ? phv_data_136 : _GEN_2192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2194 = 8'h89 == _match_key_qbytes_1_T_2 ? phv_data_137 : _GEN_2193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2195 = 8'h8a == _match_key_qbytes_1_T_2 ? phv_data_138 : _GEN_2194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2196 = 8'h8b == _match_key_qbytes_1_T_2 ? phv_data_139 : _GEN_2195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2197 = 8'h8c == _match_key_qbytes_1_T_2 ? phv_data_140 : _GEN_2196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2198 = 8'h8d == _match_key_qbytes_1_T_2 ? phv_data_141 : _GEN_2197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2199 = 8'h8e == _match_key_qbytes_1_T_2 ? phv_data_142 : _GEN_2198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2200 = 8'h8f == _match_key_qbytes_1_T_2 ? phv_data_143 : _GEN_2199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2201 = 8'h90 == _match_key_qbytes_1_T_2 ? phv_data_144 : _GEN_2200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2202 = 8'h91 == _match_key_qbytes_1_T_2 ? phv_data_145 : _GEN_2201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2203 = 8'h92 == _match_key_qbytes_1_T_2 ? phv_data_146 : _GEN_2202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2204 = 8'h93 == _match_key_qbytes_1_T_2 ? phv_data_147 : _GEN_2203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2205 = 8'h94 == _match_key_qbytes_1_T_2 ? phv_data_148 : _GEN_2204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2206 = 8'h95 == _match_key_qbytes_1_T_2 ? phv_data_149 : _GEN_2205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2207 = 8'h96 == _match_key_qbytes_1_T_2 ? phv_data_150 : _GEN_2206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2208 = 8'h97 == _match_key_qbytes_1_T_2 ? phv_data_151 : _GEN_2207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2209 = 8'h98 == _match_key_qbytes_1_T_2 ? phv_data_152 : _GEN_2208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2210 = 8'h99 == _match_key_qbytes_1_T_2 ? phv_data_153 : _GEN_2209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2211 = 8'h9a == _match_key_qbytes_1_T_2 ? phv_data_154 : _GEN_2210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2212 = 8'h9b == _match_key_qbytes_1_T_2 ? phv_data_155 : _GEN_2211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2213 = 8'h9c == _match_key_qbytes_1_T_2 ? phv_data_156 : _GEN_2212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2214 = 8'h9d == _match_key_qbytes_1_T_2 ? phv_data_157 : _GEN_2213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2215 = 8'h9e == _match_key_qbytes_1_T_2 ? phv_data_158 : _GEN_2214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2216 = 8'h9f == _match_key_qbytes_1_T_2 ? phv_data_159 : _GEN_2215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2217 = 8'ha0 == _match_key_qbytes_1_T_2 ? phv_data_160 : _GEN_2216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2218 = 8'ha1 == _match_key_qbytes_1_T_2 ? phv_data_161 : _GEN_2217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2219 = 8'ha2 == _match_key_qbytes_1_T_2 ? phv_data_162 : _GEN_2218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2220 = 8'ha3 == _match_key_qbytes_1_T_2 ? phv_data_163 : _GEN_2219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2221 = 8'ha4 == _match_key_qbytes_1_T_2 ? phv_data_164 : _GEN_2220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2222 = 8'ha5 == _match_key_qbytes_1_T_2 ? phv_data_165 : _GEN_2221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2223 = 8'ha6 == _match_key_qbytes_1_T_2 ? phv_data_166 : _GEN_2222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2224 = 8'ha7 == _match_key_qbytes_1_T_2 ? phv_data_167 : _GEN_2223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2225 = 8'ha8 == _match_key_qbytes_1_T_2 ? phv_data_168 : _GEN_2224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2226 = 8'ha9 == _match_key_qbytes_1_T_2 ? phv_data_169 : _GEN_2225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2227 = 8'haa == _match_key_qbytes_1_T_2 ? phv_data_170 : _GEN_2226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2228 = 8'hab == _match_key_qbytes_1_T_2 ? phv_data_171 : _GEN_2227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2229 = 8'hac == _match_key_qbytes_1_T_2 ? phv_data_172 : _GEN_2228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2230 = 8'had == _match_key_qbytes_1_T_2 ? phv_data_173 : _GEN_2229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2231 = 8'hae == _match_key_qbytes_1_T_2 ? phv_data_174 : _GEN_2230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2232 = 8'haf == _match_key_qbytes_1_T_2 ? phv_data_175 : _GEN_2231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2233 = 8'hb0 == _match_key_qbytes_1_T_2 ? phv_data_176 : _GEN_2232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2234 = 8'hb1 == _match_key_qbytes_1_T_2 ? phv_data_177 : _GEN_2233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2235 = 8'hb2 == _match_key_qbytes_1_T_2 ? phv_data_178 : _GEN_2234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2236 = 8'hb3 == _match_key_qbytes_1_T_2 ? phv_data_179 : _GEN_2235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2237 = 8'hb4 == _match_key_qbytes_1_T_2 ? phv_data_180 : _GEN_2236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2238 = 8'hb5 == _match_key_qbytes_1_T_2 ? phv_data_181 : _GEN_2237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2239 = 8'hb6 == _match_key_qbytes_1_T_2 ? phv_data_182 : _GEN_2238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2240 = 8'hb7 == _match_key_qbytes_1_T_2 ? phv_data_183 : _GEN_2239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2241 = 8'hb8 == _match_key_qbytes_1_T_2 ? phv_data_184 : _GEN_2240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2242 = 8'hb9 == _match_key_qbytes_1_T_2 ? phv_data_185 : _GEN_2241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2243 = 8'hba == _match_key_qbytes_1_T_2 ? phv_data_186 : _GEN_2242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2244 = 8'hbb == _match_key_qbytes_1_T_2 ? phv_data_187 : _GEN_2243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2245 = 8'hbc == _match_key_qbytes_1_T_2 ? phv_data_188 : _GEN_2244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2246 = 8'hbd == _match_key_qbytes_1_T_2 ? phv_data_189 : _GEN_2245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2247 = 8'hbe == _match_key_qbytes_1_T_2 ? phv_data_190 : _GEN_2246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2248 = 8'hbf == _match_key_qbytes_1_T_2 ? phv_data_191 : _GEN_2247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2249 = 8'hc0 == _match_key_qbytes_1_T_2 ? phv_data_192 : _GEN_2248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2250 = 8'hc1 == _match_key_qbytes_1_T_2 ? phv_data_193 : _GEN_2249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2251 = 8'hc2 == _match_key_qbytes_1_T_2 ? phv_data_194 : _GEN_2250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2252 = 8'hc3 == _match_key_qbytes_1_T_2 ? phv_data_195 : _GEN_2251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2253 = 8'hc4 == _match_key_qbytes_1_T_2 ? phv_data_196 : _GEN_2252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2254 = 8'hc5 == _match_key_qbytes_1_T_2 ? phv_data_197 : _GEN_2253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2255 = 8'hc6 == _match_key_qbytes_1_T_2 ? phv_data_198 : _GEN_2254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2256 = 8'hc7 == _match_key_qbytes_1_T_2 ? phv_data_199 : _GEN_2255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2257 = 8'hc8 == _match_key_qbytes_1_T_2 ? phv_data_200 : _GEN_2256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2258 = 8'hc9 == _match_key_qbytes_1_T_2 ? phv_data_201 : _GEN_2257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2259 = 8'hca == _match_key_qbytes_1_T_2 ? phv_data_202 : _GEN_2258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2260 = 8'hcb == _match_key_qbytes_1_T_2 ? phv_data_203 : _GEN_2259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2261 = 8'hcc == _match_key_qbytes_1_T_2 ? phv_data_204 : _GEN_2260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2262 = 8'hcd == _match_key_qbytes_1_T_2 ? phv_data_205 : _GEN_2261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2263 = 8'hce == _match_key_qbytes_1_T_2 ? phv_data_206 : _GEN_2262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2264 = 8'hcf == _match_key_qbytes_1_T_2 ? phv_data_207 : _GEN_2263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2265 = 8'hd0 == _match_key_qbytes_1_T_2 ? phv_data_208 : _GEN_2264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2266 = 8'hd1 == _match_key_qbytes_1_T_2 ? phv_data_209 : _GEN_2265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2267 = 8'hd2 == _match_key_qbytes_1_T_2 ? phv_data_210 : _GEN_2266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2268 = 8'hd3 == _match_key_qbytes_1_T_2 ? phv_data_211 : _GEN_2267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2269 = 8'hd4 == _match_key_qbytes_1_T_2 ? phv_data_212 : _GEN_2268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2270 = 8'hd5 == _match_key_qbytes_1_T_2 ? phv_data_213 : _GEN_2269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2271 = 8'hd6 == _match_key_qbytes_1_T_2 ? phv_data_214 : _GEN_2270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2272 = 8'hd7 == _match_key_qbytes_1_T_2 ? phv_data_215 : _GEN_2271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2273 = 8'hd8 == _match_key_qbytes_1_T_2 ? phv_data_216 : _GEN_2272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2274 = 8'hd9 == _match_key_qbytes_1_T_2 ? phv_data_217 : _GEN_2273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2275 = 8'hda == _match_key_qbytes_1_T_2 ? phv_data_218 : _GEN_2274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2276 = 8'hdb == _match_key_qbytes_1_T_2 ? phv_data_219 : _GEN_2275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2277 = 8'hdc == _match_key_qbytes_1_T_2 ? phv_data_220 : _GEN_2276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2278 = 8'hdd == _match_key_qbytes_1_T_2 ? phv_data_221 : _GEN_2277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2279 = 8'hde == _match_key_qbytes_1_T_2 ? phv_data_222 : _GEN_2278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2280 = 8'hdf == _match_key_qbytes_1_T_2 ? phv_data_223 : _GEN_2279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2281 = 8'he0 == _match_key_qbytes_1_T_2 ? phv_data_224 : _GEN_2280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2282 = 8'he1 == _match_key_qbytes_1_T_2 ? phv_data_225 : _GEN_2281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2283 = 8'he2 == _match_key_qbytes_1_T_2 ? phv_data_226 : _GEN_2282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2284 = 8'he3 == _match_key_qbytes_1_T_2 ? phv_data_227 : _GEN_2283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2285 = 8'he4 == _match_key_qbytes_1_T_2 ? phv_data_228 : _GEN_2284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2286 = 8'he5 == _match_key_qbytes_1_T_2 ? phv_data_229 : _GEN_2285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2287 = 8'he6 == _match_key_qbytes_1_T_2 ? phv_data_230 : _GEN_2286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2288 = 8'he7 == _match_key_qbytes_1_T_2 ? phv_data_231 : _GEN_2287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2289 = 8'he8 == _match_key_qbytes_1_T_2 ? phv_data_232 : _GEN_2288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2290 = 8'he9 == _match_key_qbytes_1_T_2 ? phv_data_233 : _GEN_2289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2291 = 8'hea == _match_key_qbytes_1_T_2 ? phv_data_234 : _GEN_2290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2292 = 8'heb == _match_key_qbytes_1_T_2 ? phv_data_235 : _GEN_2291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2293 = 8'hec == _match_key_qbytes_1_T_2 ? phv_data_236 : _GEN_2292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2294 = 8'hed == _match_key_qbytes_1_T_2 ? phv_data_237 : _GEN_2293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2295 = 8'hee == _match_key_qbytes_1_T_2 ? phv_data_238 : _GEN_2294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2296 = 8'hef == _match_key_qbytes_1_T_2 ? phv_data_239 : _GEN_2295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2297 = 8'hf0 == _match_key_qbytes_1_T_2 ? phv_data_240 : _GEN_2296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2298 = 8'hf1 == _match_key_qbytes_1_T_2 ? phv_data_241 : _GEN_2297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2299 = 8'hf2 == _match_key_qbytes_1_T_2 ? phv_data_242 : _GEN_2298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2300 = 8'hf3 == _match_key_qbytes_1_T_2 ? phv_data_243 : _GEN_2299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2301 = 8'hf4 == _match_key_qbytes_1_T_2 ? phv_data_244 : _GEN_2300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2302 = 8'hf5 == _match_key_qbytes_1_T_2 ? phv_data_245 : _GEN_2301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2303 = 8'hf6 == _match_key_qbytes_1_T_2 ? phv_data_246 : _GEN_2302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2304 = 8'hf7 == _match_key_qbytes_1_T_2 ? phv_data_247 : _GEN_2303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2305 = 8'hf8 == _match_key_qbytes_1_T_2 ? phv_data_248 : _GEN_2304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2306 = 8'hf9 == _match_key_qbytes_1_T_2 ? phv_data_249 : _GEN_2305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2307 = 8'hfa == _match_key_qbytes_1_T_2 ? phv_data_250 : _GEN_2306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2308 = 8'hfb == _match_key_qbytes_1_T_2 ? phv_data_251 : _GEN_2307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2309 = 8'hfc == _match_key_qbytes_1_T_2 ? phv_data_252 : _GEN_2308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2310 = 8'hfd == _match_key_qbytes_1_T_2 ? phv_data_253 : _GEN_2309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2311 = 8'hfe == _match_key_qbytes_1_T_2 ? phv_data_254 : _GEN_2310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2312 = 8'hff == _match_key_qbytes_1_T_2 ? phv_data_255 : _GEN_2311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_13350 = {{1'd0}, _match_key_qbytes_1_T_2}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2313 = 9'h100 == _GEN_13350 ? phv_data_256 : _GEN_2312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2314 = 9'h101 == _GEN_13350 ? phv_data_257 : _GEN_2313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2315 = 9'h102 == _GEN_13350 ? phv_data_258 : _GEN_2314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2316 = 9'h103 == _GEN_13350 ? phv_data_259 : _GEN_2315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2317 = 9'h104 == _GEN_13350 ? phv_data_260 : _GEN_2316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2318 = 9'h105 == _GEN_13350 ? phv_data_261 : _GEN_2317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2319 = 9'h106 == _GEN_13350 ? phv_data_262 : _GEN_2318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2320 = 9'h107 == _GEN_13350 ? phv_data_263 : _GEN_2319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2321 = 9'h108 == _GEN_13350 ? phv_data_264 : _GEN_2320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2322 = 9'h109 == _GEN_13350 ? phv_data_265 : _GEN_2321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2323 = 9'h10a == _GEN_13350 ? phv_data_266 : _GEN_2322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2324 = 9'h10b == _GEN_13350 ? phv_data_267 : _GEN_2323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2325 = 9'h10c == _GEN_13350 ? phv_data_268 : _GEN_2324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2326 = 9'h10d == _GEN_13350 ? phv_data_269 : _GEN_2325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2327 = 9'h10e == _GEN_13350 ? phv_data_270 : _GEN_2326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2328 = 9'h10f == _GEN_13350 ? phv_data_271 : _GEN_2327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2329 = 9'h110 == _GEN_13350 ? phv_data_272 : _GEN_2328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2330 = 9'h111 == _GEN_13350 ? phv_data_273 : _GEN_2329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2331 = 9'h112 == _GEN_13350 ? phv_data_274 : _GEN_2330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2332 = 9'h113 == _GEN_13350 ? phv_data_275 : _GEN_2331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2333 = 9'h114 == _GEN_13350 ? phv_data_276 : _GEN_2332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2334 = 9'h115 == _GEN_13350 ? phv_data_277 : _GEN_2333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2335 = 9'h116 == _GEN_13350 ? phv_data_278 : _GEN_2334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2336 = 9'h117 == _GEN_13350 ? phv_data_279 : _GEN_2335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2337 = 9'h118 == _GEN_13350 ? phv_data_280 : _GEN_2336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2338 = 9'h119 == _GEN_13350 ? phv_data_281 : _GEN_2337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2339 = 9'h11a == _GEN_13350 ? phv_data_282 : _GEN_2338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2340 = 9'h11b == _GEN_13350 ? phv_data_283 : _GEN_2339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2341 = 9'h11c == _GEN_13350 ? phv_data_284 : _GEN_2340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2342 = 9'h11d == _GEN_13350 ? phv_data_285 : _GEN_2341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2343 = 9'h11e == _GEN_13350 ? phv_data_286 : _GEN_2342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2344 = 9'h11f == _GEN_13350 ? phv_data_287 : _GEN_2343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2345 = 9'h120 == _GEN_13350 ? phv_data_288 : _GEN_2344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2346 = 9'h121 == _GEN_13350 ? phv_data_289 : _GEN_2345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2347 = 9'h122 == _GEN_13350 ? phv_data_290 : _GEN_2346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2348 = 9'h123 == _GEN_13350 ? phv_data_291 : _GEN_2347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2349 = 9'h124 == _GEN_13350 ? phv_data_292 : _GEN_2348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2350 = 9'h125 == _GEN_13350 ? phv_data_293 : _GEN_2349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2351 = 9'h126 == _GEN_13350 ? phv_data_294 : _GEN_2350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2352 = 9'h127 == _GEN_13350 ? phv_data_295 : _GEN_2351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2353 = 9'h128 == _GEN_13350 ? phv_data_296 : _GEN_2352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2354 = 9'h129 == _GEN_13350 ? phv_data_297 : _GEN_2353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2355 = 9'h12a == _GEN_13350 ? phv_data_298 : _GEN_2354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2356 = 9'h12b == _GEN_13350 ? phv_data_299 : _GEN_2355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2357 = 9'h12c == _GEN_13350 ? phv_data_300 : _GEN_2356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2358 = 9'h12d == _GEN_13350 ? phv_data_301 : _GEN_2357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2359 = 9'h12e == _GEN_13350 ? phv_data_302 : _GEN_2358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2360 = 9'h12f == _GEN_13350 ? phv_data_303 : _GEN_2359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2361 = 9'h130 == _GEN_13350 ? phv_data_304 : _GEN_2360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2362 = 9'h131 == _GEN_13350 ? phv_data_305 : _GEN_2361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2363 = 9'h132 == _GEN_13350 ? phv_data_306 : _GEN_2362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2364 = 9'h133 == _GEN_13350 ? phv_data_307 : _GEN_2363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2365 = 9'h134 == _GEN_13350 ? phv_data_308 : _GEN_2364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2366 = 9'h135 == _GEN_13350 ? phv_data_309 : _GEN_2365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2367 = 9'h136 == _GEN_13350 ? phv_data_310 : _GEN_2366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2368 = 9'h137 == _GEN_13350 ? phv_data_311 : _GEN_2367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2369 = 9'h138 == _GEN_13350 ? phv_data_312 : _GEN_2368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2370 = 9'h139 == _GEN_13350 ? phv_data_313 : _GEN_2369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2371 = 9'h13a == _GEN_13350 ? phv_data_314 : _GEN_2370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2372 = 9'h13b == _GEN_13350 ? phv_data_315 : _GEN_2371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2373 = 9'h13c == _GEN_13350 ? phv_data_316 : _GEN_2372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2374 = 9'h13d == _GEN_13350 ? phv_data_317 : _GEN_2373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2375 = 9'h13e == _GEN_13350 ? phv_data_318 : _GEN_2374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2376 = 9'h13f == _GEN_13350 ? phv_data_319 : _GEN_2375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2377 = 9'h140 == _GEN_13350 ? phv_data_320 : _GEN_2376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2378 = 9'h141 == _GEN_13350 ? phv_data_321 : _GEN_2377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2379 = 9'h142 == _GEN_13350 ? phv_data_322 : _GEN_2378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2380 = 9'h143 == _GEN_13350 ? phv_data_323 : _GEN_2379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2381 = 9'h144 == _GEN_13350 ? phv_data_324 : _GEN_2380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2382 = 9'h145 == _GEN_13350 ? phv_data_325 : _GEN_2381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2383 = 9'h146 == _GEN_13350 ? phv_data_326 : _GEN_2382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2384 = 9'h147 == _GEN_13350 ? phv_data_327 : _GEN_2383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2385 = 9'h148 == _GEN_13350 ? phv_data_328 : _GEN_2384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2386 = 9'h149 == _GEN_13350 ? phv_data_329 : _GEN_2385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2387 = 9'h14a == _GEN_13350 ? phv_data_330 : _GEN_2386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2388 = 9'h14b == _GEN_13350 ? phv_data_331 : _GEN_2387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2389 = 9'h14c == _GEN_13350 ? phv_data_332 : _GEN_2388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2390 = 9'h14d == _GEN_13350 ? phv_data_333 : _GEN_2389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2391 = 9'h14e == _GEN_13350 ? phv_data_334 : _GEN_2390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2392 = 9'h14f == _GEN_13350 ? phv_data_335 : _GEN_2391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2393 = 9'h150 == _GEN_13350 ? phv_data_336 : _GEN_2392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2394 = 9'h151 == _GEN_13350 ? phv_data_337 : _GEN_2393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2395 = 9'h152 == _GEN_13350 ? phv_data_338 : _GEN_2394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2396 = 9'h153 == _GEN_13350 ? phv_data_339 : _GEN_2395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2397 = 9'h154 == _GEN_13350 ? phv_data_340 : _GEN_2396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2398 = 9'h155 == _GEN_13350 ? phv_data_341 : _GEN_2397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2399 = 9'h156 == _GEN_13350 ? phv_data_342 : _GEN_2398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2400 = 9'h157 == _GEN_13350 ? phv_data_343 : _GEN_2399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2401 = 9'h158 == _GEN_13350 ? phv_data_344 : _GEN_2400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2402 = 9'h159 == _GEN_13350 ? phv_data_345 : _GEN_2401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2403 = 9'h15a == _GEN_13350 ? phv_data_346 : _GEN_2402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2404 = 9'h15b == _GEN_13350 ? phv_data_347 : _GEN_2403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2405 = 9'h15c == _GEN_13350 ? phv_data_348 : _GEN_2404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2406 = 9'h15d == _GEN_13350 ? phv_data_349 : _GEN_2405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2407 = 9'h15e == _GEN_13350 ? phv_data_350 : _GEN_2406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2408 = 9'h15f == _GEN_13350 ? phv_data_351 : _GEN_2407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2409 = 9'h160 == _GEN_13350 ? phv_data_352 : _GEN_2408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2410 = 9'h161 == _GEN_13350 ? phv_data_353 : _GEN_2409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2411 = 9'h162 == _GEN_13350 ? phv_data_354 : _GEN_2410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2412 = 9'h163 == _GEN_13350 ? phv_data_355 : _GEN_2411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2413 = 9'h164 == _GEN_13350 ? phv_data_356 : _GEN_2412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2414 = 9'h165 == _GEN_13350 ? phv_data_357 : _GEN_2413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2415 = 9'h166 == _GEN_13350 ? phv_data_358 : _GEN_2414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2416 = 9'h167 == _GEN_13350 ? phv_data_359 : _GEN_2415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2417 = 9'h168 == _GEN_13350 ? phv_data_360 : _GEN_2416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2418 = 9'h169 == _GEN_13350 ? phv_data_361 : _GEN_2417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2419 = 9'h16a == _GEN_13350 ? phv_data_362 : _GEN_2418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2420 = 9'h16b == _GEN_13350 ? phv_data_363 : _GEN_2419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2421 = 9'h16c == _GEN_13350 ? phv_data_364 : _GEN_2420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2422 = 9'h16d == _GEN_13350 ? phv_data_365 : _GEN_2421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2423 = 9'h16e == _GEN_13350 ? phv_data_366 : _GEN_2422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2424 = 9'h16f == _GEN_13350 ? phv_data_367 : _GEN_2423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2425 = 9'h170 == _GEN_13350 ? phv_data_368 : _GEN_2424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2426 = 9'h171 == _GEN_13350 ? phv_data_369 : _GEN_2425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2427 = 9'h172 == _GEN_13350 ? phv_data_370 : _GEN_2426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2428 = 9'h173 == _GEN_13350 ? phv_data_371 : _GEN_2427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2429 = 9'h174 == _GEN_13350 ? phv_data_372 : _GEN_2428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2430 = 9'h175 == _GEN_13350 ? phv_data_373 : _GEN_2429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2431 = 9'h176 == _GEN_13350 ? phv_data_374 : _GEN_2430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2432 = 9'h177 == _GEN_13350 ? phv_data_375 : _GEN_2431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2433 = 9'h178 == _GEN_13350 ? phv_data_376 : _GEN_2432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2434 = 9'h179 == _GEN_13350 ? phv_data_377 : _GEN_2433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2435 = 9'h17a == _GEN_13350 ? phv_data_378 : _GEN_2434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2436 = 9'h17b == _GEN_13350 ? phv_data_379 : _GEN_2435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2437 = 9'h17c == _GEN_13350 ? phv_data_380 : _GEN_2436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2438 = 9'h17d == _GEN_13350 ? phv_data_381 : _GEN_2437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2439 = 9'h17e == _GEN_13350 ? phv_data_382 : _GEN_2438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2440 = 9'h17f == _GEN_13350 ? phv_data_383 : _GEN_2439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2441 = 9'h180 == _GEN_13350 ? phv_data_384 : _GEN_2440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2442 = 9'h181 == _GEN_13350 ? phv_data_385 : _GEN_2441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2443 = 9'h182 == _GEN_13350 ? phv_data_386 : _GEN_2442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2444 = 9'h183 == _GEN_13350 ? phv_data_387 : _GEN_2443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2445 = 9'h184 == _GEN_13350 ? phv_data_388 : _GEN_2444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2446 = 9'h185 == _GEN_13350 ? phv_data_389 : _GEN_2445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2447 = 9'h186 == _GEN_13350 ? phv_data_390 : _GEN_2446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2448 = 9'h187 == _GEN_13350 ? phv_data_391 : _GEN_2447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2449 = 9'h188 == _GEN_13350 ? phv_data_392 : _GEN_2448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2450 = 9'h189 == _GEN_13350 ? phv_data_393 : _GEN_2449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2451 = 9'h18a == _GEN_13350 ? phv_data_394 : _GEN_2450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2452 = 9'h18b == _GEN_13350 ? phv_data_395 : _GEN_2451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2453 = 9'h18c == _GEN_13350 ? phv_data_396 : _GEN_2452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2454 = 9'h18d == _GEN_13350 ? phv_data_397 : _GEN_2453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2455 = 9'h18e == _GEN_13350 ? phv_data_398 : _GEN_2454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2456 = 9'h18f == _GEN_13350 ? phv_data_399 : _GEN_2455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2457 = 9'h190 == _GEN_13350 ? phv_data_400 : _GEN_2456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2458 = 9'h191 == _GEN_13350 ? phv_data_401 : _GEN_2457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2459 = 9'h192 == _GEN_13350 ? phv_data_402 : _GEN_2458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2460 = 9'h193 == _GEN_13350 ? phv_data_403 : _GEN_2459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2461 = 9'h194 == _GEN_13350 ? phv_data_404 : _GEN_2460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2462 = 9'h195 == _GEN_13350 ? phv_data_405 : _GEN_2461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2463 = 9'h196 == _GEN_13350 ? phv_data_406 : _GEN_2462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2464 = 9'h197 == _GEN_13350 ? phv_data_407 : _GEN_2463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2465 = 9'h198 == _GEN_13350 ? phv_data_408 : _GEN_2464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2466 = 9'h199 == _GEN_13350 ? phv_data_409 : _GEN_2465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2467 = 9'h19a == _GEN_13350 ? phv_data_410 : _GEN_2466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2468 = 9'h19b == _GEN_13350 ? phv_data_411 : _GEN_2467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2469 = 9'h19c == _GEN_13350 ? phv_data_412 : _GEN_2468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2470 = 9'h19d == _GEN_13350 ? phv_data_413 : _GEN_2469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2471 = 9'h19e == _GEN_13350 ? phv_data_414 : _GEN_2470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2472 = 9'h19f == _GEN_13350 ? phv_data_415 : _GEN_2471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2473 = 9'h1a0 == _GEN_13350 ? phv_data_416 : _GEN_2472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2474 = 9'h1a1 == _GEN_13350 ? phv_data_417 : _GEN_2473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2475 = 9'h1a2 == _GEN_13350 ? phv_data_418 : _GEN_2474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2476 = 9'h1a3 == _GEN_13350 ? phv_data_419 : _GEN_2475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2477 = 9'h1a4 == _GEN_13350 ? phv_data_420 : _GEN_2476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2478 = 9'h1a5 == _GEN_13350 ? phv_data_421 : _GEN_2477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2479 = 9'h1a6 == _GEN_13350 ? phv_data_422 : _GEN_2478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2480 = 9'h1a7 == _GEN_13350 ? phv_data_423 : _GEN_2479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2481 = 9'h1a8 == _GEN_13350 ? phv_data_424 : _GEN_2480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2482 = 9'h1a9 == _GEN_13350 ? phv_data_425 : _GEN_2481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2483 = 9'h1aa == _GEN_13350 ? phv_data_426 : _GEN_2482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2484 = 9'h1ab == _GEN_13350 ? phv_data_427 : _GEN_2483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2485 = 9'h1ac == _GEN_13350 ? phv_data_428 : _GEN_2484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2486 = 9'h1ad == _GEN_13350 ? phv_data_429 : _GEN_2485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2487 = 9'h1ae == _GEN_13350 ? phv_data_430 : _GEN_2486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2488 = 9'h1af == _GEN_13350 ? phv_data_431 : _GEN_2487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2489 = 9'h1b0 == _GEN_13350 ? phv_data_432 : _GEN_2488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2490 = 9'h1b1 == _GEN_13350 ? phv_data_433 : _GEN_2489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2491 = 9'h1b2 == _GEN_13350 ? phv_data_434 : _GEN_2490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2492 = 9'h1b3 == _GEN_13350 ? phv_data_435 : _GEN_2491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2493 = 9'h1b4 == _GEN_13350 ? phv_data_436 : _GEN_2492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2494 = 9'h1b5 == _GEN_13350 ? phv_data_437 : _GEN_2493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2495 = 9'h1b6 == _GEN_13350 ? phv_data_438 : _GEN_2494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2496 = 9'h1b7 == _GEN_13350 ? phv_data_439 : _GEN_2495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2497 = 9'h1b8 == _GEN_13350 ? phv_data_440 : _GEN_2496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2498 = 9'h1b9 == _GEN_13350 ? phv_data_441 : _GEN_2497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2499 = 9'h1ba == _GEN_13350 ? phv_data_442 : _GEN_2498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2500 = 9'h1bb == _GEN_13350 ? phv_data_443 : _GEN_2499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2501 = 9'h1bc == _GEN_13350 ? phv_data_444 : _GEN_2500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2502 = 9'h1bd == _GEN_13350 ? phv_data_445 : _GEN_2501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2503 = 9'h1be == _GEN_13350 ? phv_data_446 : _GEN_2502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2504 = 9'h1bf == _GEN_13350 ? phv_data_447 : _GEN_2503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2505 = 9'h1c0 == _GEN_13350 ? phv_data_448 : _GEN_2504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2506 = 9'h1c1 == _GEN_13350 ? phv_data_449 : _GEN_2505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2507 = 9'h1c2 == _GEN_13350 ? phv_data_450 : _GEN_2506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2508 = 9'h1c3 == _GEN_13350 ? phv_data_451 : _GEN_2507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2509 = 9'h1c4 == _GEN_13350 ? phv_data_452 : _GEN_2508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2510 = 9'h1c5 == _GEN_13350 ? phv_data_453 : _GEN_2509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2511 = 9'h1c6 == _GEN_13350 ? phv_data_454 : _GEN_2510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2512 = 9'h1c7 == _GEN_13350 ? phv_data_455 : _GEN_2511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2513 = 9'h1c8 == _GEN_13350 ? phv_data_456 : _GEN_2512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2514 = 9'h1c9 == _GEN_13350 ? phv_data_457 : _GEN_2513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2515 = 9'h1ca == _GEN_13350 ? phv_data_458 : _GEN_2514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2516 = 9'h1cb == _GEN_13350 ? phv_data_459 : _GEN_2515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2517 = 9'h1cc == _GEN_13350 ? phv_data_460 : _GEN_2516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2518 = 9'h1cd == _GEN_13350 ? phv_data_461 : _GEN_2517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2519 = 9'h1ce == _GEN_13350 ? phv_data_462 : _GEN_2518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2520 = 9'h1cf == _GEN_13350 ? phv_data_463 : _GEN_2519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2521 = 9'h1d0 == _GEN_13350 ? phv_data_464 : _GEN_2520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2522 = 9'h1d1 == _GEN_13350 ? phv_data_465 : _GEN_2521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2523 = 9'h1d2 == _GEN_13350 ? phv_data_466 : _GEN_2522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2524 = 9'h1d3 == _GEN_13350 ? phv_data_467 : _GEN_2523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2525 = 9'h1d4 == _GEN_13350 ? phv_data_468 : _GEN_2524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2526 = 9'h1d5 == _GEN_13350 ? phv_data_469 : _GEN_2525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2527 = 9'h1d6 == _GEN_13350 ? phv_data_470 : _GEN_2526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2528 = 9'h1d7 == _GEN_13350 ? phv_data_471 : _GEN_2527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2529 = 9'h1d8 == _GEN_13350 ? phv_data_472 : _GEN_2528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2530 = 9'h1d9 == _GEN_13350 ? phv_data_473 : _GEN_2529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2531 = 9'h1da == _GEN_13350 ? phv_data_474 : _GEN_2530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2532 = 9'h1db == _GEN_13350 ? phv_data_475 : _GEN_2531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2533 = 9'h1dc == _GEN_13350 ? phv_data_476 : _GEN_2532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2534 = 9'h1dd == _GEN_13350 ? phv_data_477 : _GEN_2533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2535 = 9'h1de == _GEN_13350 ? phv_data_478 : _GEN_2534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2536 = 9'h1df == _GEN_13350 ? phv_data_479 : _GEN_2535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2537 = 9'h1e0 == _GEN_13350 ? phv_data_480 : _GEN_2536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2538 = 9'h1e1 == _GEN_13350 ? phv_data_481 : _GEN_2537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2539 = 9'h1e2 == _GEN_13350 ? phv_data_482 : _GEN_2538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2540 = 9'h1e3 == _GEN_13350 ? phv_data_483 : _GEN_2539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2541 = 9'h1e4 == _GEN_13350 ? phv_data_484 : _GEN_2540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2542 = 9'h1e5 == _GEN_13350 ? phv_data_485 : _GEN_2541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2543 = 9'h1e6 == _GEN_13350 ? phv_data_486 : _GEN_2542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2544 = 9'h1e7 == _GEN_13350 ? phv_data_487 : _GEN_2543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2545 = 9'h1e8 == _GEN_13350 ? phv_data_488 : _GEN_2544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2546 = 9'h1e9 == _GEN_13350 ? phv_data_489 : _GEN_2545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2547 = 9'h1ea == _GEN_13350 ? phv_data_490 : _GEN_2546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2548 = 9'h1eb == _GEN_13350 ? phv_data_491 : _GEN_2547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2549 = 9'h1ec == _GEN_13350 ? phv_data_492 : _GEN_2548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2550 = 9'h1ed == _GEN_13350 ? phv_data_493 : _GEN_2549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2551 = 9'h1ee == _GEN_13350 ? phv_data_494 : _GEN_2550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2552 = 9'h1ef == _GEN_13350 ? phv_data_495 : _GEN_2551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2553 = 9'h1f0 == _GEN_13350 ? phv_data_496 : _GEN_2552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2554 = 9'h1f1 == _GEN_13350 ? phv_data_497 : _GEN_2553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2555 = 9'h1f2 == _GEN_13350 ? phv_data_498 : _GEN_2554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2556 = 9'h1f3 == _GEN_13350 ? phv_data_499 : _GEN_2555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2557 = 9'h1f4 == _GEN_13350 ? phv_data_500 : _GEN_2556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2558 = 9'h1f5 == _GEN_13350 ? phv_data_501 : _GEN_2557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2559 = 9'h1f6 == _GEN_13350 ? phv_data_502 : _GEN_2558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2560 = 9'h1f7 == _GEN_13350 ? phv_data_503 : _GEN_2559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2561 = 9'h1f8 == _GEN_13350 ? phv_data_504 : _GEN_2560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2562 = 9'h1f9 == _GEN_13350 ? phv_data_505 : _GEN_2561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2563 = 9'h1fa == _GEN_13350 ? phv_data_506 : _GEN_2562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2564 = 9'h1fb == _GEN_13350 ? phv_data_507 : _GEN_2563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2565 = 9'h1fc == _GEN_13350 ? phv_data_508 : _GEN_2564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2566 = 9'h1fd == _GEN_13350 ? phv_data_509 : _GEN_2565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2567 = 9'h1fe == _GEN_13350 ? phv_data_510 : _GEN_2566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2568 = 9'h1ff == _GEN_13350 ? phv_data_511 : _GEN_2567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2570 = 8'h1 == local_offset_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2571 = 8'h2 == local_offset_1 ? phv_data_2 : _GEN_2570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2572 = 8'h3 == local_offset_1 ? phv_data_3 : _GEN_2571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2573 = 8'h4 == local_offset_1 ? phv_data_4 : _GEN_2572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2574 = 8'h5 == local_offset_1 ? phv_data_5 : _GEN_2573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2575 = 8'h6 == local_offset_1 ? phv_data_6 : _GEN_2574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2576 = 8'h7 == local_offset_1 ? phv_data_7 : _GEN_2575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2577 = 8'h8 == local_offset_1 ? phv_data_8 : _GEN_2576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2578 = 8'h9 == local_offset_1 ? phv_data_9 : _GEN_2577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2579 = 8'ha == local_offset_1 ? phv_data_10 : _GEN_2578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2580 = 8'hb == local_offset_1 ? phv_data_11 : _GEN_2579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2581 = 8'hc == local_offset_1 ? phv_data_12 : _GEN_2580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2582 = 8'hd == local_offset_1 ? phv_data_13 : _GEN_2581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2583 = 8'he == local_offset_1 ? phv_data_14 : _GEN_2582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2584 = 8'hf == local_offset_1 ? phv_data_15 : _GEN_2583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2585 = 8'h10 == local_offset_1 ? phv_data_16 : _GEN_2584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2586 = 8'h11 == local_offset_1 ? phv_data_17 : _GEN_2585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2587 = 8'h12 == local_offset_1 ? phv_data_18 : _GEN_2586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2588 = 8'h13 == local_offset_1 ? phv_data_19 : _GEN_2587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2589 = 8'h14 == local_offset_1 ? phv_data_20 : _GEN_2588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2590 = 8'h15 == local_offset_1 ? phv_data_21 : _GEN_2589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2591 = 8'h16 == local_offset_1 ? phv_data_22 : _GEN_2590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2592 = 8'h17 == local_offset_1 ? phv_data_23 : _GEN_2591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2593 = 8'h18 == local_offset_1 ? phv_data_24 : _GEN_2592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2594 = 8'h19 == local_offset_1 ? phv_data_25 : _GEN_2593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2595 = 8'h1a == local_offset_1 ? phv_data_26 : _GEN_2594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2596 = 8'h1b == local_offset_1 ? phv_data_27 : _GEN_2595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2597 = 8'h1c == local_offset_1 ? phv_data_28 : _GEN_2596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2598 = 8'h1d == local_offset_1 ? phv_data_29 : _GEN_2597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2599 = 8'h1e == local_offset_1 ? phv_data_30 : _GEN_2598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2600 = 8'h1f == local_offset_1 ? phv_data_31 : _GEN_2599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2601 = 8'h20 == local_offset_1 ? phv_data_32 : _GEN_2600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2602 = 8'h21 == local_offset_1 ? phv_data_33 : _GEN_2601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2603 = 8'h22 == local_offset_1 ? phv_data_34 : _GEN_2602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2604 = 8'h23 == local_offset_1 ? phv_data_35 : _GEN_2603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2605 = 8'h24 == local_offset_1 ? phv_data_36 : _GEN_2604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2606 = 8'h25 == local_offset_1 ? phv_data_37 : _GEN_2605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2607 = 8'h26 == local_offset_1 ? phv_data_38 : _GEN_2606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2608 = 8'h27 == local_offset_1 ? phv_data_39 : _GEN_2607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2609 = 8'h28 == local_offset_1 ? phv_data_40 : _GEN_2608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2610 = 8'h29 == local_offset_1 ? phv_data_41 : _GEN_2609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2611 = 8'h2a == local_offset_1 ? phv_data_42 : _GEN_2610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2612 = 8'h2b == local_offset_1 ? phv_data_43 : _GEN_2611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2613 = 8'h2c == local_offset_1 ? phv_data_44 : _GEN_2612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2614 = 8'h2d == local_offset_1 ? phv_data_45 : _GEN_2613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2615 = 8'h2e == local_offset_1 ? phv_data_46 : _GEN_2614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2616 = 8'h2f == local_offset_1 ? phv_data_47 : _GEN_2615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2617 = 8'h30 == local_offset_1 ? phv_data_48 : _GEN_2616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2618 = 8'h31 == local_offset_1 ? phv_data_49 : _GEN_2617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2619 = 8'h32 == local_offset_1 ? phv_data_50 : _GEN_2618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2620 = 8'h33 == local_offset_1 ? phv_data_51 : _GEN_2619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2621 = 8'h34 == local_offset_1 ? phv_data_52 : _GEN_2620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2622 = 8'h35 == local_offset_1 ? phv_data_53 : _GEN_2621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2623 = 8'h36 == local_offset_1 ? phv_data_54 : _GEN_2622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2624 = 8'h37 == local_offset_1 ? phv_data_55 : _GEN_2623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2625 = 8'h38 == local_offset_1 ? phv_data_56 : _GEN_2624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2626 = 8'h39 == local_offset_1 ? phv_data_57 : _GEN_2625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2627 = 8'h3a == local_offset_1 ? phv_data_58 : _GEN_2626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2628 = 8'h3b == local_offset_1 ? phv_data_59 : _GEN_2627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2629 = 8'h3c == local_offset_1 ? phv_data_60 : _GEN_2628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2630 = 8'h3d == local_offset_1 ? phv_data_61 : _GEN_2629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2631 = 8'h3e == local_offset_1 ? phv_data_62 : _GEN_2630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2632 = 8'h3f == local_offset_1 ? phv_data_63 : _GEN_2631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2633 = 8'h40 == local_offset_1 ? phv_data_64 : _GEN_2632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2634 = 8'h41 == local_offset_1 ? phv_data_65 : _GEN_2633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2635 = 8'h42 == local_offset_1 ? phv_data_66 : _GEN_2634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2636 = 8'h43 == local_offset_1 ? phv_data_67 : _GEN_2635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2637 = 8'h44 == local_offset_1 ? phv_data_68 : _GEN_2636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2638 = 8'h45 == local_offset_1 ? phv_data_69 : _GEN_2637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2639 = 8'h46 == local_offset_1 ? phv_data_70 : _GEN_2638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2640 = 8'h47 == local_offset_1 ? phv_data_71 : _GEN_2639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2641 = 8'h48 == local_offset_1 ? phv_data_72 : _GEN_2640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2642 = 8'h49 == local_offset_1 ? phv_data_73 : _GEN_2641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2643 = 8'h4a == local_offset_1 ? phv_data_74 : _GEN_2642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2644 = 8'h4b == local_offset_1 ? phv_data_75 : _GEN_2643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2645 = 8'h4c == local_offset_1 ? phv_data_76 : _GEN_2644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2646 = 8'h4d == local_offset_1 ? phv_data_77 : _GEN_2645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2647 = 8'h4e == local_offset_1 ? phv_data_78 : _GEN_2646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2648 = 8'h4f == local_offset_1 ? phv_data_79 : _GEN_2647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2649 = 8'h50 == local_offset_1 ? phv_data_80 : _GEN_2648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2650 = 8'h51 == local_offset_1 ? phv_data_81 : _GEN_2649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2651 = 8'h52 == local_offset_1 ? phv_data_82 : _GEN_2650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2652 = 8'h53 == local_offset_1 ? phv_data_83 : _GEN_2651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2653 = 8'h54 == local_offset_1 ? phv_data_84 : _GEN_2652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2654 = 8'h55 == local_offset_1 ? phv_data_85 : _GEN_2653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2655 = 8'h56 == local_offset_1 ? phv_data_86 : _GEN_2654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2656 = 8'h57 == local_offset_1 ? phv_data_87 : _GEN_2655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2657 = 8'h58 == local_offset_1 ? phv_data_88 : _GEN_2656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2658 = 8'h59 == local_offset_1 ? phv_data_89 : _GEN_2657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2659 = 8'h5a == local_offset_1 ? phv_data_90 : _GEN_2658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2660 = 8'h5b == local_offset_1 ? phv_data_91 : _GEN_2659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2661 = 8'h5c == local_offset_1 ? phv_data_92 : _GEN_2660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2662 = 8'h5d == local_offset_1 ? phv_data_93 : _GEN_2661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2663 = 8'h5e == local_offset_1 ? phv_data_94 : _GEN_2662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2664 = 8'h5f == local_offset_1 ? phv_data_95 : _GEN_2663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2665 = 8'h60 == local_offset_1 ? phv_data_96 : _GEN_2664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2666 = 8'h61 == local_offset_1 ? phv_data_97 : _GEN_2665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2667 = 8'h62 == local_offset_1 ? phv_data_98 : _GEN_2666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2668 = 8'h63 == local_offset_1 ? phv_data_99 : _GEN_2667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2669 = 8'h64 == local_offset_1 ? phv_data_100 : _GEN_2668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2670 = 8'h65 == local_offset_1 ? phv_data_101 : _GEN_2669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2671 = 8'h66 == local_offset_1 ? phv_data_102 : _GEN_2670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2672 = 8'h67 == local_offset_1 ? phv_data_103 : _GEN_2671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2673 = 8'h68 == local_offset_1 ? phv_data_104 : _GEN_2672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2674 = 8'h69 == local_offset_1 ? phv_data_105 : _GEN_2673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2675 = 8'h6a == local_offset_1 ? phv_data_106 : _GEN_2674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2676 = 8'h6b == local_offset_1 ? phv_data_107 : _GEN_2675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2677 = 8'h6c == local_offset_1 ? phv_data_108 : _GEN_2676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2678 = 8'h6d == local_offset_1 ? phv_data_109 : _GEN_2677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2679 = 8'h6e == local_offset_1 ? phv_data_110 : _GEN_2678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2680 = 8'h6f == local_offset_1 ? phv_data_111 : _GEN_2679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2681 = 8'h70 == local_offset_1 ? phv_data_112 : _GEN_2680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2682 = 8'h71 == local_offset_1 ? phv_data_113 : _GEN_2681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2683 = 8'h72 == local_offset_1 ? phv_data_114 : _GEN_2682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2684 = 8'h73 == local_offset_1 ? phv_data_115 : _GEN_2683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2685 = 8'h74 == local_offset_1 ? phv_data_116 : _GEN_2684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2686 = 8'h75 == local_offset_1 ? phv_data_117 : _GEN_2685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2687 = 8'h76 == local_offset_1 ? phv_data_118 : _GEN_2686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2688 = 8'h77 == local_offset_1 ? phv_data_119 : _GEN_2687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2689 = 8'h78 == local_offset_1 ? phv_data_120 : _GEN_2688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2690 = 8'h79 == local_offset_1 ? phv_data_121 : _GEN_2689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2691 = 8'h7a == local_offset_1 ? phv_data_122 : _GEN_2690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2692 = 8'h7b == local_offset_1 ? phv_data_123 : _GEN_2691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2693 = 8'h7c == local_offset_1 ? phv_data_124 : _GEN_2692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2694 = 8'h7d == local_offset_1 ? phv_data_125 : _GEN_2693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2695 = 8'h7e == local_offset_1 ? phv_data_126 : _GEN_2694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2696 = 8'h7f == local_offset_1 ? phv_data_127 : _GEN_2695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2697 = 8'h80 == local_offset_1 ? phv_data_128 : _GEN_2696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2698 = 8'h81 == local_offset_1 ? phv_data_129 : _GEN_2697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2699 = 8'h82 == local_offset_1 ? phv_data_130 : _GEN_2698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2700 = 8'h83 == local_offset_1 ? phv_data_131 : _GEN_2699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2701 = 8'h84 == local_offset_1 ? phv_data_132 : _GEN_2700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2702 = 8'h85 == local_offset_1 ? phv_data_133 : _GEN_2701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2703 = 8'h86 == local_offset_1 ? phv_data_134 : _GEN_2702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2704 = 8'h87 == local_offset_1 ? phv_data_135 : _GEN_2703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2705 = 8'h88 == local_offset_1 ? phv_data_136 : _GEN_2704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2706 = 8'h89 == local_offset_1 ? phv_data_137 : _GEN_2705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2707 = 8'h8a == local_offset_1 ? phv_data_138 : _GEN_2706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2708 = 8'h8b == local_offset_1 ? phv_data_139 : _GEN_2707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2709 = 8'h8c == local_offset_1 ? phv_data_140 : _GEN_2708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2710 = 8'h8d == local_offset_1 ? phv_data_141 : _GEN_2709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2711 = 8'h8e == local_offset_1 ? phv_data_142 : _GEN_2710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2712 = 8'h8f == local_offset_1 ? phv_data_143 : _GEN_2711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2713 = 8'h90 == local_offset_1 ? phv_data_144 : _GEN_2712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2714 = 8'h91 == local_offset_1 ? phv_data_145 : _GEN_2713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2715 = 8'h92 == local_offset_1 ? phv_data_146 : _GEN_2714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2716 = 8'h93 == local_offset_1 ? phv_data_147 : _GEN_2715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2717 = 8'h94 == local_offset_1 ? phv_data_148 : _GEN_2716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2718 = 8'h95 == local_offset_1 ? phv_data_149 : _GEN_2717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2719 = 8'h96 == local_offset_1 ? phv_data_150 : _GEN_2718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2720 = 8'h97 == local_offset_1 ? phv_data_151 : _GEN_2719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2721 = 8'h98 == local_offset_1 ? phv_data_152 : _GEN_2720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2722 = 8'h99 == local_offset_1 ? phv_data_153 : _GEN_2721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2723 = 8'h9a == local_offset_1 ? phv_data_154 : _GEN_2722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2724 = 8'h9b == local_offset_1 ? phv_data_155 : _GEN_2723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2725 = 8'h9c == local_offset_1 ? phv_data_156 : _GEN_2724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2726 = 8'h9d == local_offset_1 ? phv_data_157 : _GEN_2725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2727 = 8'h9e == local_offset_1 ? phv_data_158 : _GEN_2726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2728 = 8'h9f == local_offset_1 ? phv_data_159 : _GEN_2727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2729 = 8'ha0 == local_offset_1 ? phv_data_160 : _GEN_2728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2730 = 8'ha1 == local_offset_1 ? phv_data_161 : _GEN_2729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2731 = 8'ha2 == local_offset_1 ? phv_data_162 : _GEN_2730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2732 = 8'ha3 == local_offset_1 ? phv_data_163 : _GEN_2731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2733 = 8'ha4 == local_offset_1 ? phv_data_164 : _GEN_2732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2734 = 8'ha5 == local_offset_1 ? phv_data_165 : _GEN_2733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2735 = 8'ha6 == local_offset_1 ? phv_data_166 : _GEN_2734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2736 = 8'ha7 == local_offset_1 ? phv_data_167 : _GEN_2735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2737 = 8'ha8 == local_offset_1 ? phv_data_168 : _GEN_2736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2738 = 8'ha9 == local_offset_1 ? phv_data_169 : _GEN_2737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2739 = 8'haa == local_offset_1 ? phv_data_170 : _GEN_2738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2740 = 8'hab == local_offset_1 ? phv_data_171 : _GEN_2739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2741 = 8'hac == local_offset_1 ? phv_data_172 : _GEN_2740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2742 = 8'had == local_offset_1 ? phv_data_173 : _GEN_2741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2743 = 8'hae == local_offset_1 ? phv_data_174 : _GEN_2742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2744 = 8'haf == local_offset_1 ? phv_data_175 : _GEN_2743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2745 = 8'hb0 == local_offset_1 ? phv_data_176 : _GEN_2744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2746 = 8'hb1 == local_offset_1 ? phv_data_177 : _GEN_2745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2747 = 8'hb2 == local_offset_1 ? phv_data_178 : _GEN_2746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2748 = 8'hb3 == local_offset_1 ? phv_data_179 : _GEN_2747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2749 = 8'hb4 == local_offset_1 ? phv_data_180 : _GEN_2748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2750 = 8'hb5 == local_offset_1 ? phv_data_181 : _GEN_2749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2751 = 8'hb6 == local_offset_1 ? phv_data_182 : _GEN_2750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2752 = 8'hb7 == local_offset_1 ? phv_data_183 : _GEN_2751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2753 = 8'hb8 == local_offset_1 ? phv_data_184 : _GEN_2752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2754 = 8'hb9 == local_offset_1 ? phv_data_185 : _GEN_2753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2755 = 8'hba == local_offset_1 ? phv_data_186 : _GEN_2754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2756 = 8'hbb == local_offset_1 ? phv_data_187 : _GEN_2755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2757 = 8'hbc == local_offset_1 ? phv_data_188 : _GEN_2756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2758 = 8'hbd == local_offset_1 ? phv_data_189 : _GEN_2757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2759 = 8'hbe == local_offset_1 ? phv_data_190 : _GEN_2758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2760 = 8'hbf == local_offset_1 ? phv_data_191 : _GEN_2759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2761 = 8'hc0 == local_offset_1 ? phv_data_192 : _GEN_2760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2762 = 8'hc1 == local_offset_1 ? phv_data_193 : _GEN_2761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2763 = 8'hc2 == local_offset_1 ? phv_data_194 : _GEN_2762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2764 = 8'hc3 == local_offset_1 ? phv_data_195 : _GEN_2763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2765 = 8'hc4 == local_offset_1 ? phv_data_196 : _GEN_2764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2766 = 8'hc5 == local_offset_1 ? phv_data_197 : _GEN_2765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2767 = 8'hc6 == local_offset_1 ? phv_data_198 : _GEN_2766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2768 = 8'hc7 == local_offset_1 ? phv_data_199 : _GEN_2767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2769 = 8'hc8 == local_offset_1 ? phv_data_200 : _GEN_2768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2770 = 8'hc9 == local_offset_1 ? phv_data_201 : _GEN_2769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2771 = 8'hca == local_offset_1 ? phv_data_202 : _GEN_2770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2772 = 8'hcb == local_offset_1 ? phv_data_203 : _GEN_2771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2773 = 8'hcc == local_offset_1 ? phv_data_204 : _GEN_2772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2774 = 8'hcd == local_offset_1 ? phv_data_205 : _GEN_2773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2775 = 8'hce == local_offset_1 ? phv_data_206 : _GEN_2774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2776 = 8'hcf == local_offset_1 ? phv_data_207 : _GEN_2775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2777 = 8'hd0 == local_offset_1 ? phv_data_208 : _GEN_2776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2778 = 8'hd1 == local_offset_1 ? phv_data_209 : _GEN_2777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2779 = 8'hd2 == local_offset_1 ? phv_data_210 : _GEN_2778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2780 = 8'hd3 == local_offset_1 ? phv_data_211 : _GEN_2779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2781 = 8'hd4 == local_offset_1 ? phv_data_212 : _GEN_2780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2782 = 8'hd5 == local_offset_1 ? phv_data_213 : _GEN_2781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2783 = 8'hd6 == local_offset_1 ? phv_data_214 : _GEN_2782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2784 = 8'hd7 == local_offset_1 ? phv_data_215 : _GEN_2783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2785 = 8'hd8 == local_offset_1 ? phv_data_216 : _GEN_2784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2786 = 8'hd9 == local_offset_1 ? phv_data_217 : _GEN_2785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2787 = 8'hda == local_offset_1 ? phv_data_218 : _GEN_2786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2788 = 8'hdb == local_offset_1 ? phv_data_219 : _GEN_2787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2789 = 8'hdc == local_offset_1 ? phv_data_220 : _GEN_2788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2790 = 8'hdd == local_offset_1 ? phv_data_221 : _GEN_2789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2791 = 8'hde == local_offset_1 ? phv_data_222 : _GEN_2790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2792 = 8'hdf == local_offset_1 ? phv_data_223 : _GEN_2791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2793 = 8'he0 == local_offset_1 ? phv_data_224 : _GEN_2792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2794 = 8'he1 == local_offset_1 ? phv_data_225 : _GEN_2793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2795 = 8'he2 == local_offset_1 ? phv_data_226 : _GEN_2794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2796 = 8'he3 == local_offset_1 ? phv_data_227 : _GEN_2795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2797 = 8'he4 == local_offset_1 ? phv_data_228 : _GEN_2796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2798 = 8'he5 == local_offset_1 ? phv_data_229 : _GEN_2797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2799 = 8'he6 == local_offset_1 ? phv_data_230 : _GEN_2798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2800 = 8'he7 == local_offset_1 ? phv_data_231 : _GEN_2799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2801 = 8'he8 == local_offset_1 ? phv_data_232 : _GEN_2800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2802 = 8'he9 == local_offset_1 ? phv_data_233 : _GEN_2801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2803 = 8'hea == local_offset_1 ? phv_data_234 : _GEN_2802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2804 = 8'heb == local_offset_1 ? phv_data_235 : _GEN_2803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2805 = 8'hec == local_offset_1 ? phv_data_236 : _GEN_2804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2806 = 8'hed == local_offset_1 ? phv_data_237 : _GEN_2805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2807 = 8'hee == local_offset_1 ? phv_data_238 : _GEN_2806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2808 = 8'hef == local_offset_1 ? phv_data_239 : _GEN_2807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2809 = 8'hf0 == local_offset_1 ? phv_data_240 : _GEN_2808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2810 = 8'hf1 == local_offset_1 ? phv_data_241 : _GEN_2809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2811 = 8'hf2 == local_offset_1 ? phv_data_242 : _GEN_2810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2812 = 8'hf3 == local_offset_1 ? phv_data_243 : _GEN_2811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2813 = 8'hf4 == local_offset_1 ? phv_data_244 : _GEN_2812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2814 = 8'hf5 == local_offset_1 ? phv_data_245 : _GEN_2813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2815 = 8'hf6 == local_offset_1 ? phv_data_246 : _GEN_2814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2816 = 8'hf7 == local_offset_1 ? phv_data_247 : _GEN_2815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2817 = 8'hf8 == local_offset_1 ? phv_data_248 : _GEN_2816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2818 = 8'hf9 == local_offset_1 ? phv_data_249 : _GEN_2817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2819 = 8'hfa == local_offset_1 ? phv_data_250 : _GEN_2818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2820 = 8'hfb == local_offset_1 ? phv_data_251 : _GEN_2819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2821 = 8'hfc == local_offset_1 ? phv_data_252 : _GEN_2820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2822 = 8'hfd == local_offset_1 ? phv_data_253 : _GEN_2821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2823 = 8'hfe == local_offset_1 ? phv_data_254 : _GEN_2822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2824 = 8'hff == local_offset_1 ? phv_data_255 : _GEN_2823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_13606 = {{1'd0}, local_offset_1}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2825 = 9'h100 == _GEN_13606 ? phv_data_256 : _GEN_2824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2826 = 9'h101 == _GEN_13606 ? phv_data_257 : _GEN_2825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2827 = 9'h102 == _GEN_13606 ? phv_data_258 : _GEN_2826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2828 = 9'h103 == _GEN_13606 ? phv_data_259 : _GEN_2827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2829 = 9'h104 == _GEN_13606 ? phv_data_260 : _GEN_2828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2830 = 9'h105 == _GEN_13606 ? phv_data_261 : _GEN_2829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2831 = 9'h106 == _GEN_13606 ? phv_data_262 : _GEN_2830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2832 = 9'h107 == _GEN_13606 ? phv_data_263 : _GEN_2831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2833 = 9'h108 == _GEN_13606 ? phv_data_264 : _GEN_2832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2834 = 9'h109 == _GEN_13606 ? phv_data_265 : _GEN_2833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2835 = 9'h10a == _GEN_13606 ? phv_data_266 : _GEN_2834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2836 = 9'h10b == _GEN_13606 ? phv_data_267 : _GEN_2835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2837 = 9'h10c == _GEN_13606 ? phv_data_268 : _GEN_2836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2838 = 9'h10d == _GEN_13606 ? phv_data_269 : _GEN_2837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2839 = 9'h10e == _GEN_13606 ? phv_data_270 : _GEN_2838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2840 = 9'h10f == _GEN_13606 ? phv_data_271 : _GEN_2839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2841 = 9'h110 == _GEN_13606 ? phv_data_272 : _GEN_2840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2842 = 9'h111 == _GEN_13606 ? phv_data_273 : _GEN_2841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2843 = 9'h112 == _GEN_13606 ? phv_data_274 : _GEN_2842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2844 = 9'h113 == _GEN_13606 ? phv_data_275 : _GEN_2843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2845 = 9'h114 == _GEN_13606 ? phv_data_276 : _GEN_2844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2846 = 9'h115 == _GEN_13606 ? phv_data_277 : _GEN_2845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2847 = 9'h116 == _GEN_13606 ? phv_data_278 : _GEN_2846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2848 = 9'h117 == _GEN_13606 ? phv_data_279 : _GEN_2847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2849 = 9'h118 == _GEN_13606 ? phv_data_280 : _GEN_2848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2850 = 9'h119 == _GEN_13606 ? phv_data_281 : _GEN_2849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2851 = 9'h11a == _GEN_13606 ? phv_data_282 : _GEN_2850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2852 = 9'h11b == _GEN_13606 ? phv_data_283 : _GEN_2851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2853 = 9'h11c == _GEN_13606 ? phv_data_284 : _GEN_2852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2854 = 9'h11d == _GEN_13606 ? phv_data_285 : _GEN_2853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2855 = 9'h11e == _GEN_13606 ? phv_data_286 : _GEN_2854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2856 = 9'h11f == _GEN_13606 ? phv_data_287 : _GEN_2855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2857 = 9'h120 == _GEN_13606 ? phv_data_288 : _GEN_2856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2858 = 9'h121 == _GEN_13606 ? phv_data_289 : _GEN_2857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2859 = 9'h122 == _GEN_13606 ? phv_data_290 : _GEN_2858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2860 = 9'h123 == _GEN_13606 ? phv_data_291 : _GEN_2859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2861 = 9'h124 == _GEN_13606 ? phv_data_292 : _GEN_2860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2862 = 9'h125 == _GEN_13606 ? phv_data_293 : _GEN_2861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2863 = 9'h126 == _GEN_13606 ? phv_data_294 : _GEN_2862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2864 = 9'h127 == _GEN_13606 ? phv_data_295 : _GEN_2863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2865 = 9'h128 == _GEN_13606 ? phv_data_296 : _GEN_2864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2866 = 9'h129 == _GEN_13606 ? phv_data_297 : _GEN_2865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2867 = 9'h12a == _GEN_13606 ? phv_data_298 : _GEN_2866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2868 = 9'h12b == _GEN_13606 ? phv_data_299 : _GEN_2867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2869 = 9'h12c == _GEN_13606 ? phv_data_300 : _GEN_2868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2870 = 9'h12d == _GEN_13606 ? phv_data_301 : _GEN_2869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2871 = 9'h12e == _GEN_13606 ? phv_data_302 : _GEN_2870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2872 = 9'h12f == _GEN_13606 ? phv_data_303 : _GEN_2871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2873 = 9'h130 == _GEN_13606 ? phv_data_304 : _GEN_2872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2874 = 9'h131 == _GEN_13606 ? phv_data_305 : _GEN_2873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2875 = 9'h132 == _GEN_13606 ? phv_data_306 : _GEN_2874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2876 = 9'h133 == _GEN_13606 ? phv_data_307 : _GEN_2875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2877 = 9'h134 == _GEN_13606 ? phv_data_308 : _GEN_2876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2878 = 9'h135 == _GEN_13606 ? phv_data_309 : _GEN_2877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2879 = 9'h136 == _GEN_13606 ? phv_data_310 : _GEN_2878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2880 = 9'h137 == _GEN_13606 ? phv_data_311 : _GEN_2879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2881 = 9'h138 == _GEN_13606 ? phv_data_312 : _GEN_2880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2882 = 9'h139 == _GEN_13606 ? phv_data_313 : _GEN_2881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2883 = 9'h13a == _GEN_13606 ? phv_data_314 : _GEN_2882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2884 = 9'h13b == _GEN_13606 ? phv_data_315 : _GEN_2883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2885 = 9'h13c == _GEN_13606 ? phv_data_316 : _GEN_2884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2886 = 9'h13d == _GEN_13606 ? phv_data_317 : _GEN_2885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2887 = 9'h13e == _GEN_13606 ? phv_data_318 : _GEN_2886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2888 = 9'h13f == _GEN_13606 ? phv_data_319 : _GEN_2887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2889 = 9'h140 == _GEN_13606 ? phv_data_320 : _GEN_2888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2890 = 9'h141 == _GEN_13606 ? phv_data_321 : _GEN_2889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2891 = 9'h142 == _GEN_13606 ? phv_data_322 : _GEN_2890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2892 = 9'h143 == _GEN_13606 ? phv_data_323 : _GEN_2891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2893 = 9'h144 == _GEN_13606 ? phv_data_324 : _GEN_2892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2894 = 9'h145 == _GEN_13606 ? phv_data_325 : _GEN_2893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2895 = 9'h146 == _GEN_13606 ? phv_data_326 : _GEN_2894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2896 = 9'h147 == _GEN_13606 ? phv_data_327 : _GEN_2895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2897 = 9'h148 == _GEN_13606 ? phv_data_328 : _GEN_2896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2898 = 9'h149 == _GEN_13606 ? phv_data_329 : _GEN_2897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2899 = 9'h14a == _GEN_13606 ? phv_data_330 : _GEN_2898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2900 = 9'h14b == _GEN_13606 ? phv_data_331 : _GEN_2899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2901 = 9'h14c == _GEN_13606 ? phv_data_332 : _GEN_2900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2902 = 9'h14d == _GEN_13606 ? phv_data_333 : _GEN_2901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2903 = 9'h14e == _GEN_13606 ? phv_data_334 : _GEN_2902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2904 = 9'h14f == _GEN_13606 ? phv_data_335 : _GEN_2903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2905 = 9'h150 == _GEN_13606 ? phv_data_336 : _GEN_2904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2906 = 9'h151 == _GEN_13606 ? phv_data_337 : _GEN_2905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2907 = 9'h152 == _GEN_13606 ? phv_data_338 : _GEN_2906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2908 = 9'h153 == _GEN_13606 ? phv_data_339 : _GEN_2907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2909 = 9'h154 == _GEN_13606 ? phv_data_340 : _GEN_2908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2910 = 9'h155 == _GEN_13606 ? phv_data_341 : _GEN_2909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2911 = 9'h156 == _GEN_13606 ? phv_data_342 : _GEN_2910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2912 = 9'h157 == _GEN_13606 ? phv_data_343 : _GEN_2911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2913 = 9'h158 == _GEN_13606 ? phv_data_344 : _GEN_2912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2914 = 9'h159 == _GEN_13606 ? phv_data_345 : _GEN_2913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2915 = 9'h15a == _GEN_13606 ? phv_data_346 : _GEN_2914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2916 = 9'h15b == _GEN_13606 ? phv_data_347 : _GEN_2915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2917 = 9'h15c == _GEN_13606 ? phv_data_348 : _GEN_2916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2918 = 9'h15d == _GEN_13606 ? phv_data_349 : _GEN_2917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2919 = 9'h15e == _GEN_13606 ? phv_data_350 : _GEN_2918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2920 = 9'h15f == _GEN_13606 ? phv_data_351 : _GEN_2919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2921 = 9'h160 == _GEN_13606 ? phv_data_352 : _GEN_2920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2922 = 9'h161 == _GEN_13606 ? phv_data_353 : _GEN_2921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2923 = 9'h162 == _GEN_13606 ? phv_data_354 : _GEN_2922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2924 = 9'h163 == _GEN_13606 ? phv_data_355 : _GEN_2923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2925 = 9'h164 == _GEN_13606 ? phv_data_356 : _GEN_2924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2926 = 9'h165 == _GEN_13606 ? phv_data_357 : _GEN_2925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2927 = 9'h166 == _GEN_13606 ? phv_data_358 : _GEN_2926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2928 = 9'h167 == _GEN_13606 ? phv_data_359 : _GEN_2927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2929 = 9'h168 == _GEN_13606 ? phv_data_360 : _GEN_2928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2930 = 9'h169 == _GEN_13606 ? phv_data_361 : _GEN_2929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2931 = 9'h16a == _GEN_13606 ? phv_data_362 : _GEN_2930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2932 = 9'h16b == _GEN_13606 ? phv_data_363 : _GEN_2931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2933 = 9'h16c == _GEN_13606 ? phv_data_364 : _GEN_2932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2934 = 9'h16d == _GEN_13606 ? phv_data_365 : _GEN_2933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2935 = 9'h16e == _GEN_13606 ? phv_data_366 : _GEN_2934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2936 = 9'h16f == _GEN_13606 ? phv_data_367 : _GEN_2935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2937 = 9'h170 == _GEN_13606 ? phv_data_368 : _GEN_2936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2938 = 9'h171 == _GEN_13606 ? phv_data_369 : _GEN_2937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2939 = 9'h172 == _GEN_13606 ? phv_data_370 : _GEN_2938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2940 = 9'h173 == _GEN_13606 ? phv_data_371 : _GEN_2939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2941 = 9'h174 == _GEN_13606 ? phv_data_372 : _GEN_2940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2942 = 9'h175 == _GEN_13606 ? phv_data_373 : _GEN_2941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2943 = 9'h176 == _GEN_13606 ? phv_data_374 : _GEN_2942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2944 = 9'h177 == _GEN_13606 ? phv_data_375 : _GEN_2943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2945 = 9'h178 == _GEN_13606 ? phv_data_376 : _GEN_2944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2946 = 9'h179 == _GEN_13606 ? phv_data_377 : _GEN_2945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2947 = 9'h17a == _GEN_13606 ? phv_data_378 : _GEN_2946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2948 = 9'h17b == _GEN_13606 ? phv_data_379 : _GEN_2947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2949 = 9'h17c == _GEN_13606 ? phv_data_380 : _GEN_2948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2950 = 9'h17d == _GEN_13606 ? phv_data_381 : _GEN_2949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2951 = 9'h17e == _GEN_13606 ? phv_data_382 : _GEN_2950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2952 = 9'h17f == _GEN_13606 ? phv_data_383 : _GEN_2951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2953 = 9'h180 == _GEN_13606 ? phv_data_384 : _GEN_2952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2954 = 9'h181 == _GEN_13606 ? phv_data_385 : _GEN_2953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2955 = 9'h182 == _GEN_13606 ? phv_data_386 : _GEN_2954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2956 = 9'h183 == _GEN_13606 ? phv_data_387 : _GEN_2955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2957 = 9'h184 == _GEN_13606 ? phv_data_388 : _GEN_2956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2958 = 9'h185 == _GEN_13606 ? phv_data_389 : _GEN_2957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2959 = 9'h186 == _GEN_13606 ? phv_data_390 : _GEN_2958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2960 = 9'h187 == _GEN_13606 ? phv_data_391 : _GEN_2959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2961 = 9'h188 == _GEN_13606 ? phv_data_392 : _GEN_2960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2962 = 9'h189 == _GEN_13606 ? phv_data_393 : _GEN_2961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2963 = 9'h18a == _GEN_13606 ? phv_data_394 : _GEN_2962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2964 = 9'h18b == _GEN_13606 ? phv_data_395 : _GEN_2963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2965 = 9'h18c == _GEN_13606 ? phv_data_396 : _GEN_2964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2966 = 9'h18d == _GEN_13606 ? phv_data_397 : _GEN_2965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2967 = 9'h18e == _GEN_13606 ? phv_data_398 : _GEN_2966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2968 = 9'h18f == _GEN_13606 ? phv_data_399 : _GEN_2967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2969 = 9'h190 == _GEN_13606 ? phv_data_400 : _GEN_2968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2970 = 9'h191 == _GEN_13606 ? phv_data_401 : _GEN_2969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2971 = 9'h192 == _GEN_13606 ? phv_data_402 : _GEN_2970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2972 = 9'h193 == _GEN_13606 ? phv_data_403 : _GEN_2971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2973 = 9'h194 == _GEN_13606 ? phv_data_404 : _GEN_2972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2974 = 9'h195 == _GEN_13606 ? phv_data_405 : _GEN_2973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2975 = 9'h196 == _GEN_13606 ? phv_data_406 : _GEN_2974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2976 = 9'h197 == _GEN_13606 ? phv_data_407 : _GEN_2975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2977 = 9'h198 == _GEN_13606 ? phv_data_408 : _GEN_2976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2978 = 9'h199 == _GEN_13606 ? phv_data_409 : _GEN_2977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2979 = 9'h19a == _GEN_13606 ? phv_data_410 : _GEN_2978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2980 = 9'h19b == _GEN_13606 ? phv_data_411 : _GEN_2979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2981 = 9'h19c == _GEN_13606 ? phv_data_412 : _GEN_2980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2982 = 9'h19d == _GEN_13606 ? phv_data_413 : _GEN_2981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2983 = 9'h19e == _GEN_13606 ? phv_data_414 : _GEN_2982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2984 = 9'h19f == _GEN_13606 ? phv_data_415 : _GEN_2983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2985 = 9'h1a0 == _GEN_13606 ? phv_data_416 : _GEN_2984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2986 = 9'h1a1 == _GEN_13606 ? phv_data_417 : _GEN_2985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2987 = 9'h1a2 == _GEN_13606 ? phv_data_418 : _GEN_2986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2988 = 9'h1a3 == _GEN_13606 ? phv_data_419 : _GEN_2987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2989 = 9'h1a4 == _GEN_13606 ? phv_data_420 : _GEN_2988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2990 = 9'h1a5 == _GEN_13606 ? phv_data_421 : _GEN_2989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2991 = 9'h1a6 == _GEN_13606 ? phv_data_422 : _GEN_2990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2992 = 9'h1a7 == _GEN_13606 ? phv_data_423 : _GEN_2991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2993 = 9'h1a8 == _GEN_13606 ? phv_data_424 : _GEN_2992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2994 = 9'h1a9 == _GEN_13606 ? phv_data_425 : _GEN_2993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2995 = 9'h1aa == _GEN_13606 ? phv_data_426 : _GEN_2994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2996 = 9'h1ab == _GEN_13606 ? phv_data_427 : _GEN_2995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2997 = 9'h1ac == _GEN_13606 ? phv_data_428 : _GEN_2996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2998 = 9'h1ad == _GEN_13606 ? phv_data_429 : _GEN_2997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2999 = 9'h1ae == _GEN_13606 ? phv_data_430 : _GEN_2998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3000 = 9'h1af == _GEN_13606 ? phv_data_431 : _GEN_2999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3001 = 9'h1b0 == _GEN_13606 ? phv_data_432 : _GEN_3000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3002 = 9'h1b1 == _GEN_13606 ? phv_data_433 : _GEN_3001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3003 = 9'h1b2 == _GEN_13606 ? phv_data_434 : _GEN_3002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3004 = 9'h1b3 == _GEN_13606 ? phv_data_435 : _GEN_3003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3005 = 9'h1b4 == _GEN_13606 ? phv_data_436 : _GEN_3004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3006 = 9'h1b5 == _GEN_13606 ? phv_data_437 : _GEN_3005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3007 = 9'h1b6 == _GEN_13606 ? phv_data_438 : _GEN_3006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3008 = 9'h1b7 == _GEN_13606 ? phv_data_439 : _GEN_3007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3009 = 9'h1b8 == _GEN_13606 ? phv_data_440 : _GEN_3008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3010 = 9'h1b9 == _GEN_13606 ? phv_data_441 : _GEN_3009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3011 = 9'h1ba == _GEN_13606 ? phv_data_442 : _GEN_3010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3012 = 9'h1bb == _GEN_13606 ? phv_data_443 : _GEN_3011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3013 = 9'h1bc == _GEN_13606 ? phv_data_444 : _GEN_3012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3014 = 9'h1bd == _GEN_13606 ? phv_data_445 : _GEN_3013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3015 = 9'h1be == _GEN_13606 ? phv_data_446 : _GEN_3014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3016 = 9'h1bf == _GEN_13606 ? phv_data_447 : _GEN_3015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3017 = 9'h1c0 == _GEN_13606 ? phv_data_448 : _GEN_3016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3018 = 9'h1c1 == _GEN_13606 ? phv_data_449 : _GEN_3017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3019 = 9'h1c2 == _GEN_13606 ? phv_data_450 : _GEN_3018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3020 = 9'h1c3 == _GEN_13606 ? phv_data_451 : _GEN_3019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3021 = 9'h1c4 == _GEN_13606 ? phv_data_452 : _GEN_3020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3022 = 9'h1c5 == _GEN_13606 ? phv_data_453 : _GEN_3021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3023 = 9'h1c6 == _GEN_13606 ? phv_data_454 : _GEN_3022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3024 = 9'h1c7 == _GEN_13606 ? phv_data_455 : _GEN_3023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3025 = 9'h1c8 == _GEN_13606 ? phv_data_456 : _GEN_3024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3026 = 9'h1c9 == _GEN_13606 ? phv_data_457 : _GEN_3025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3027 = 9'h1ca == _GEN_13606 ? phv_data_458 : _GEN_3026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3028 = 9'h1cb == _GEN_13606 ? phv_data_459 : _GEN_3027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3029 = 9'h1cc == _GEN_13606 ? phv_data_460 : _GEN_3028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3030 = 9'h1cd == _GEN_13606 ? phv_data_461 : _GEN_3029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3031 = 9'h1ce == _GEN_13606 ? phv_data_462 : _GEN_3030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3032 = 9'h1cf == _GEN_13606 ? phv_data_463 : _GEN_3031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3033 = 9'h1d0 == _GEN_13606 ? phv_data_464 : _GEN_3032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3034 = 9'h1d1 == _GEN_13606 ? phv_data_465 : _GEN_3033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3035 = 9'h1d2 == _GEN_13606 ? phv_data_466 : _GEN_3034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3036 = 9'h1d3 == _GEN_13606 ? phv_data_467 : _GEN_3035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3037 = 9'h1d4 == _GEN_13606 ? phv_data_468 : _GEN_3036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3038 = 9'h1d5 == _GEN_13606 ? phv_data_469 : _GEN_3037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3039 = 9'h1d6 == _GEN_13606 ? phv_data_470 : _GEN_3038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3040 = 9'h1d7 == _GEN_13606 ? phv_data_471 : _GEN_3039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3041 = 9'h1d8 == _GEN_13606 ? phv_data_472 : _GEN_3040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3042 = 9'h1d9 == _GEN_13606 ? phv_data_473 : _GEN_3041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3043 = 9'h1da == _GEN_13606 ? phv_data_474 : _GEN_3042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3044 = 9'h1db == _GEN_13606 ? phv_data_475 : _GEN_3043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3045 = 9'h1dc == _GEN_13606 ? phv_data_476 : _GEN_3044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3046 = 9'h1dd == _GEN_13606 ? phv_data_477 : _GEN_3045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3047 = 9'h1de == _GEN_13606 ? phv_data_478 : _GEN_3046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3048 = 9'h1df == _GEN_13606 ? phv_data_479 : _GEN_3047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3049 = 9'h1e0 == _GEN_13606 ? phv_data_480 : _GEN_3048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3050 = 9'h1e1 == _GEN_13606 ? phv_data_481 : _GEN_3049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3051 = 9'h1e2 == _GEN_13606 ? phv_data_482 : _GEN_3050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3052 = 9'h1e3 == _GEN_13606 ? phv_data_483 : _GEN_3051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3053 = 9'h1e4 == _GEN_13606 ? phv_data_484 : _GEN_3052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3054 = 9'h1e5 == _GEN_13606 ? phv_data_485 : _GEN_3053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3055 = 9'h1e6 == _GEN_13606 ? phv_data_486 : _GEN_3054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3056 = 9'h1e7 == _GEN_13606 ? phv_data_487 : _GEN_3055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3057 = 9'h1e8 == _GEN_13606 ? phv_data_488 : _GEN_3056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3058 = 9'h1e9 == _GEN_13606 ? phv_data_489 : _GEN_3057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3059 = 9'h1ea == _GEN_13606 ? phv_data_490 : _GEN_3058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3060 = 9'h1eb == _GEN_13606 ? phv_data_491 : _GEN_3059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3061 = 9'h1ec == _GEN_13606 ? phv_data_492 : _GEN_3060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3062 = 9'h1ed == _GEN_13606 ? phv_data_493 : _GEN_3061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3063 = 9'h1ee == _GEN_13606 ? phv_data_494 : _GEN_3062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3064 = 9'h1ef == _GEN_13606 ? phv_data_495 : _GEN_3063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3065 = 9'h1f0 == _GEN_13606 ? phv_data_496 : _GEN_3064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3066 = 9'h1f1 == _GEN_13606 ? phv_data_497 : _GEN_3065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3067 = 9'h1f2 == _GEN_13606 ? phv_data_498 : _GEN_3066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3068 = 9'h1f3 == _GEN_13606 ? phv_data_499 : _GEN_3067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3069 = 9'h1f4 == _GEN_13606 ? phv_data_500 : _GEN_3068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3070 = 9'h1f5 == _GEN_13606 ? phv_data_501 : _GEN_3069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3071 = 9'h1f6 == _GEN_13606 ? phv_data_502 : _GEN_3070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3072 = 9'h1f7 == _GEN_13606 ? phv_data_503 : _GEN_3071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3073 = 9'h1f8 == _GEN_13606 ? phv_data_504 : _GEN_3072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3074 = 9'h1f9 == _GEN_13606 ? phv_data_505 : _GEN_3073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3075 = 9'h1fa == _GEN_13606 ? phv_data_506 : _GEN_3074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3076 = 9'h1fb == _GEN_13606 ? phv_data_507 : _GEN_3075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3077 = 9'h1fc == _GEN_13606 ? phv_data_508 : _GEN_3076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3078 = 9'h1fd == _GEN_13606 ? phv_data_509 : _GEN_3077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3079 = 9'h1fe == _GEN_13606 ? phv_data_510 : _GEN_3078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3080 = 9'h1ff == _GEN_13606 ? phv_data_511 : _GEN_3079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3082 = 8'h1 == _match_key_qbytes_1_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3083 = 8'h2 == _match_key_qbytes_1_T ? phv_data_2 : _GEN_3082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3084 = 8'h3 == _match_key_qbytes_1_T ? phv_data_3 : _GEN_3083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3085 = 8'h4 == _match_key_qbytes_1_T ? phv_data_4 : _GEN_3084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3086 = 8'h5 == _match_key_qbytes_1_T ? phv_data_5 : _GEN_3085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3087 = 8'h6 == _match_key_qbytes_1_T ? phv_data_6 : _GEN_3086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3088 = 8'h7 == _match_key_qbytes_1_T ? phv_data_7 : _GEN_3087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3089 = 8'h8 == _match_key_qbytes_1_T ? phv_data_8 : _GEN_3088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3090 = 8'h9 == _match_key_qbytes_1_T ? phv_data_9 : _GEN_3089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3091 = 8'ha == _match_key_qbytes_1_T ? phv_data_10 : _GEN_3090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3092 = 8'hb == _match_key_qbytes_1_T ? phv_data_11 : _GEN_3091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3093 = 8'hc == _match_key_qbytes_1_T ? phv_data_12 : _GEN_3092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3094 = 8'hd == _match_key_qbytes_1_T ? phv_data_13 : _GEN_3093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3095 = 8'he == _match_key_qbytes_1_T ? phv_data_14 : _GEN_3094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3096 = 8'hf == _match_key_qbytes_1_T ? phv_data_15 : _GEN_3095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3097 = 8'h10 == _match_key_qbytes_1_T ? phv_data_16 : _GEN_3096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3098 = 8'h11 == _match_key_qbytes_1_T ? phv_data_17 : _GEN_3097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3099 = 8'h12 == _match_key_qbytes_1_T ? phv_data_18 : _GEN_3098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3100 = 8'h13 == _match_key_qbytes_1_T ? phv_data_19 : _GEN_3099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3101 = 8'h14 == _match_key_qbytes_1_T ? phv_data_20 : _GEN_3100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3102 = 8'h15 == _match_key_qbytes_1_T ? phv_data_21 : _GEN_3101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3103 = 8'h16 == _match_key_qbytes_1_T ? phv_data_22 : _GEN_3102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3104 = 8'h17 == _match_key_qbytes_1_T ? phv_data_23 : _GEN_3103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3105 = 8'h18 == _match_key_qbytes_1_T ? phv_data_24 : _GEN_3104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3106 = 8'h19 == _match_key_qbytes_1_T ? phv_data_25 : _GEN_3105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3107 = 8'h1a == _match_key_qbytes_1_T ? phv_data_26 : _GEN_3106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3108 = 8'h1b == _match_key_qbytes_1_T ? phv_data_27 : _GEN_3107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3109 = 8'h1c == _match_key_qbytes_1_T ? phv_data_28 : _GEN_3108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3110 = 8'h1d == _match_key_qbytes_1_T ? phv_data_29 : _GEN_3109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3111 = 8'h1e == _match_key_qbytes_1_T ? phv_data_30 : _GEN_3110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3112 = 8'h1f == _match_key_qbytes_1_T ? phv_data_31 : _GEN_3111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3113 = 8'h20 == _match_key_qbytes_1_T ? phv_data_32 : _GEN_3112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3114 = 8'h21 == _match_key_qbytes_1_T ? phv_data_33 : _GEN_3113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3115 = 8'h22 == _match_key_qbytes_1_T ? phv_data_34 : _GEN_3114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3116 = 8'h23 == _match_key_qbytes_1_T ? phv_data_35 : _GEN_3115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3117 = 8'h24 == _match_key_qbytes_1_T ? phv_data_36 : _GEN_3116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3118 = 8'h25 == _match_key_qbytes_1_T ? phv_data_37 : _GEN_3117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3119 = 8'h26 == _match_key_qbytes_1_T ? phv_data_38 : _GEN_3118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3120 = 8'h27 == _match_key_qbytes_1_T ? phv_data_39 : _GEN_3119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3121 = 8'h28 == _match_key_qbytes_1_T ? phv_data_40 : _GEN_3120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3122 = 8'h29 == _match_key_qbytes_1_T ? phv_data_41 : _GEN_3121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3123 = 8'h2a == _match_key_qbytes_1_T ? phv_data_42 : _GEN_3122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3124 = 8'h2b == _match_key_qbytes_1_T ? phv_data_43 : _GEN_3123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3125 = 8'h2c == _match_key_qbytes_1_T ? phv_data_44 : _GEN_3124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3126 = 8'h2d == _match_key_qbytes_1_T ? phv_data_45 : _GEN_3125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3127 = 8'h2e == _match_key_qbytes_1_T ? phv_data_46 : _GEN_3126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3128 = 8'h2f == _match_key_qbytes_1_T ? phv_data_47 : _GEN_3127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3129 = 8'h30 == _match_key_qbytes_1_T ? phv_data_48 : _GEN_3128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3130 = 8'h31 == _match_key_qbytes_1_T ? phv_data_49 : _GEN_3129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3131 = 8'h32 == _match_key_qbytes_1_T ? phv_data_50 : _GEN_3130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3132 = 8'h33 == _match_key_qbytes_1_T ? phv_data_51 : _GEN_3131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3133 = 8'h34 == _match_key_qbytes_1_T ? phv_data_52 : _GEN_3132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3134 = 8'h35 == _match_key_qbytes_1_T ? phv_data_53 : _GEN_3133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3135 = 8'h36 == _match_key_qbytes_1_T ? phv_data_54 : _GEN_3134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3136 = 8'h37 == _match_key_qbytes_1_T ? phv_data_55 : _GEN_3135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3137 = 8'h38 == _match_key_qbytes_1_T ? phv_data_56 : _GEN_3136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3138 = 8'h39 == _match_key_qbytes_1_T ? phv_data_57 : _GEN_3137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3139 = 8'h3a == _match_key_qbytes_1_T ? phv_data_58 : _GEN_3138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3140 = 8'h3b == _match_key_qbytes_1_T ? phv_data_59 : _GEN_3139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3141 = 8'h3c == _match_key_qbytes_1_T ? phv_data_60 : _GEN_3140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3142 = 8'h3d == _match_key_qbytes_1_T ? phv_data_61 : _GEN_3141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3143 = 8'h3e == _match_key_qbytes_1_T ? phv_data_62 : _GEN_3142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3144 = 8'h3f == _match_key_qbytes_1_T ? phv_data_63 : _GEN_3143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3145 = 8'h40 == _match_key_qbytes_1_T ? phv_data_64 : _GEN_3144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3146 = 8'h41 == _match_key_qbytes_1_T ? phv_data_65 : _GEN_3145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3147 = 8'h42 == _match_key_qbytes_1_T ? phv_data_66 : _GEN_3146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3148 = 8'h43 == _match_key_qbytes_1_T ? phv_data_67 : _GEN_3147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3149 = 8'h44 == _match_key_qbytes_1_T ? phv_data_68 : _GEN_3148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3150 = 8'h45 == _match_key_qbytes_1_T ? phv_data_69 : _GEN_3149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3151 = 8'h46 == _match_key_qbytes_1_T ? phv_data_70 : _GEN_3150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3152 = 8'h47 == _match_key_qbytes_1_T ? phv_data_71 : _GEN_3151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3153 = 8'h48 == _match_key_qbytes_1_T ? phv_data_72 : _GEN_3152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3154 = 8'h49 == _match_key_qbytes_1_T ? phv_data_73 : _GEN_3153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3155 = 8'h4a == _match_key_qbytes_1_T ? phv_data_74 : _GEN_3154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3156 = 8'h4b == _match_key_qbytes_1_T ? phv_data_75 : _GEN_3155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3157 = 8'h4c == _match_key_qbytes_1_T ? phv_data_76 : _GEN_3156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3158 = 8'h4d == _match_key_qbytes_1_T ? phv_data_77 : _GEN_3157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3159 = 8'h4e == _match_key_qbytes_1_T ? phv_data_78 : _GEN_3158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3160 = 8'h4f == _match_key_qbytes_1_T ? phv_data_79 : _GEN_3159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3161 = 8'h50 == _match_key_qbytes_1_T ? phv_data_80 : _GEN_3160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3162 = 8'h51 == _match_key_qbytes_1_T ? phv_data_81 : _GEN_3161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3163 = 8'h52 == _match_key_qbytes_1_T ? phv_data_82 : _GEN_3162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3164 = 8'h53 == _match_key_qbytes_1_T ? phv_data_83 : _GEN_3163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3165 = 8'h54 == _match_key_qbytes_1_T ? phv_data_84 : _GEN_3164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3166 = 8'h55 == _match_key_qbytes_1_T ? phv_data_85 : _GEN_3165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3167 = 8'h56 == _match_key_qbytes_1_T ? phv_data_86 : _GEN_3166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3168 = 8'h57 == _match_key_qbytes_1_T ? phv_data_87 : _GEN_3167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3169 = 8'h58 == _match_key_qbytes_1_T ? phv_data_88 : _GEN_3168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3170 = 8'h59 == _match_key_qbytes_1_T ? phv_data_89 : _GEN_3169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3171 = 8'h5a == _match_key_qbytes_1_T ? phv_data_90 : _GEN_3170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3172 = 8'h5b == _match_key_qbytes_1_T ? phv_data_91 : _GEN_3171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3173 = 8'h5c == _match_key_qbytes_1_T ? phv_data_92 : _GEN_3172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3174 = 8'h5d == _match_key_qbytes_1_T ? phv_data_93 : _GEN_3173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3175 = 8'h5e == _match_key_qbytes_1_T ? phv_data_94 : _GEN_3174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3176 = 8'h5f == _match_key_qbytes_1_T ? phv_data_95 : _GEN_3175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3177 = 8'h60 == _match_key_qbytes_1_T ? phv_data_96 : _GEN_3176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3178 = 8'h61 == _match_key_qbytes_1_T ? phv_data_97 : _GEN_3177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3179 = 8'h62 == _match_key_qbytes_1_T ? phv_data_98 : _GEN_3178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3180 = 8'h63 == _match_key_qbytes_1_T ? phv_data_99 : _GEN_3179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3181 = 8'h64 == _match_key_qbytes_1_T ? phv_data_100 : _GEN_3180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3182 = 8'h65 == _match_key_qbytes_1_T ? phv_data_101 : _GEN_3181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3183 = 8'h66 == _match_key_qbytes_1_T ? phv_data_102 : _GEN_3182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3184 = 8'h67 == _match_key_qbytes_1_T ? phv_data_103 : _GEN_3183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3185 = 8'h68 == _match_key_qbytes_1_T ? phv_data_104 : _GEN_3184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3186 = 8'h69 == _match_key_qbytes_1_T ? phv_data_105 : _GEN_3185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3187 = 8'h6a == _match_key_qbytes_1_T ? phv_data_106 : _GEN_3186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3188 = 8'h6b == _match_key_qbytes_1_T ? phv_data_107 : _GEN_3187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3189 = 8'h6c == _match_key_qbytes_1_T ? phv_data_108 : _GEN_3188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3190 = 8'h6d == _match_key_qbytes_1_T ? phv_data_109 : _GEN_3189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3191 = 8'h6e == _match_key_qbytes_1_T ? phv_data_110 : _GEN_3190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3192 = 8'h6f == _match_key_qbytes_1_T ? phv_data_111 : _GEN_3191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3193 = 8'h70 == _match_key_qbytes_1_T ? phv_data_112 : _GEN_3192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3194 = 8'h71 == _match_key_qbytes_1_T ? phv_data_113 : _GEN_3193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3195 = 8'h72 == _match_key_qbytes_1_T ? phv_data_114 : _GEN_3194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3196 = 8'h73 == _match_key_qbytes_1_T ? phv_data_115 : _GEN_3195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3197 = 8'h74 == _match_key_qbytes_1_T ? phv_data_116 : _GEN_3196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3198 = 8'h75 == _match_key_qbytes_1_T ? phv_data_117 : _GEN_3197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3199 = 8'h76 == _match_key_qbytes_1_T ? phv_data_118 : _GEN_3198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3200 = 8'h77 == _match_key_qbytes_1_T ? phv_data_119 : _GEN_3199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3201 = 8'h78 == _match_key_qbytes_1_T ? phv_data_120 : _GEN_3200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3202 = 8'h79 == _match_key_qbytes_1_T ? phv_data_121 : _GEN_3201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3203 = 8'h7a == _match_key_qbytes_1_T ? phv_data_122 : _GEN_3202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3204 = 8'h7b == _match_key_qbytes_1_T ? phv_data_123 : _GEN_3203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3205 = 8'h7c == _match_key_qbytes_1_T ? phv_data_124 : _GEN_3204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3206 = 8'h7d == _match_key_qbytes_1_T ? phv_data_125 : _GEN_3205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3207 = 8'h7e == _match_key_qbytes_1_T ? phv_data_126 : _GEN_3206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3208 = 8'h7f == _match_key_qbytes_1_T ? phv_data_127 : _GEN_3207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3209 = 8'h80 == _match_key_qbytes_1_T ? phv_data_128 : _GEN_3208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3210 = 8'h81 == _match_key_qbytes_1_T ? phv_data_129 : _GEN_3209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3211 = 8'h82 == _match_key_qbytes_1_T ? phv_data_130 : _GEN_3210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3212 = 8'h83 == _match_key_qbytes_1_T ? phv_data_131 : _GEN_3211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3213 = 8'h84 == _match_key_qbytes_1_T ? phv_data_132 : _GEN_3212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3214 = 8'h85 == _match_key_qbytes_1_T ? phv_data_133 : _GEN_3213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3215 = 8'h86 == _match_key_qbytes_1_T ? phv_data_134 : _GEN_3214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3216 = 8'h87 == _match_key_qbytes_1_T ? phv_data_135 : _GEN_3215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3217 = 8'h88 == _match_key_qbytes_1_T ? phv_data_136 : _GEN_3216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3218 = 8'h89 == _match_key_qbytes_1_T ? phv_data_137 : _GEN_3217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3219 = 8'h8a == _match_key_qbytes_1_T ? phv_data_138 : _GEN_3218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3220 = 8'h8b == _match_key_qbytes_1_T ? phv_data_139 : _GEN_3219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3221 = 8'h8c == _match_key_qbytes_1_T ? phv_data_140 : _GEN_3220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3222 = 8'h8d == _match_key_qbytes_1_T ? phv_data_141 : _GEN_3221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3223 = 8'h8e == _match_key_qbytes_1_T ? phv_data_142 : _GEN_3222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3224 = 8'h8f == _match_key_qbytes_1_T ? phv_data_143 : _GEN_3223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3225 = 8'h90 == _match_key_qbytes_1_T ? phv_data_144 : _GEN_3224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3226 = 8'h91 == _match_key_qbytes_1_T ? phv_data_145 : _GEN_3225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3227 = 8'h92 == _match_key_qbytes_1_T ? phv_data_146 : _GEN_3226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3228 = 8'h93 == _match_key_qbytes_1_T ? phv_data_147 : _GEN_3227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3229 = 8'h94 == _match_key_qbytes_1_T ? phv_data_148 : _GEN_3228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3230 = 8'h95 == _match_key_qbytes_1_T ? phv_data_149 : _GEN_3229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3231 = 8'h96 == _match_key_qbytes_1_T ? phv_data_150 : _GEN_3230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3232 = 8'h97 == _match_key_qbytes_1_T ? phv_data_151 : _GEN_3231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3233 = 8'h98 == _match_key_qbytes_1_T ? phv_data_152 : _GEN_3232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3234 = 8'h99 == _match_key_qbytes_1_T ? phv_data_153 : _GEN_3233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3235 = 8'h9a == _match_key_qbytes_1_T ? phv_data_154 : _GEN_3234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3236 = 8'h9b == _match_key_qbytes_1_T ? phv_data_155 : _GEN_3235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3237 = 8'h9c == _match_key_qbytes_1_T ? phv_data_156 : _GEN_3236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3238 = 8'h9d == _match_key_qbytes_1_T ? phv_data_157 : _GEN_3237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3239 = 8'h9e == _match_key_qbytes_1_T ? phv_data_158 : _GEN_3238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3240 = 8'h9f == _match_key_qbytes_1_T ? phv_data_159 : _GEN_3239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3241 = 8'ha0 == _match_key_qbytes_1_T ? phv_data_160 : _GEN_3240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3242 = 8'ha1 == _match_key_qbytes_1_T ? phv_data_161 : _GEN_3241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3243 = 8'ha2 == _match_key_qbytes_1_T ? phv_data_162 : _GEN_3242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3244 = 8'ha3 == _match_key_qbytes_1_T ? phv_data_163 : _GEN_3243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3245 = 8'ha4 == _match_key_qbytes_1_T ? phv_data_164 : _GEN_3244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3246 = 8'ha5 == _match_key_qbytes_1_T ? phv_data_165 : _GEN_3245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3247 = 8'ha6 == _match_key_qbytes_1_T ? phv_data_166 : _GEN_3246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3248 = 8'ha7 == _match_key_qbytes_1_T ? phv_data_167 : _GEN_3247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3249 = 8'ha8 == _match_key_qbytes_1_T ? phv_data_168 : _GEN_3248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3250 = 8'ha9 == _match_key_qbytes_1_T ? phv_data_169 : _GEN_3249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3251 = 8'haa == _match_key_qbytes_1_T ? phv_data_170 : _GEN_3250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3252 = 8'hab == _match_key_qbytes_1_T ? phv_data_171 : _GEN_3251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3253 = 8'hac == _match_key_qbytes_1_T ? phv_data_172 : _GEN_3252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3254 = 8'had == _match_key_qbytes_1_T ? phv_data_173 : _GEN_3253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3255 = 8'hae == _match_key_qbytes_1_T ? phv_data_174 : _GEN_3254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3256 = 8'haf == _match_key_qbytes_1_T ? phv_data_175 : _GEN_3255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3257 = 8'hb0 == _match_key_qbytes_1_T ? phv_data_176 : _GEN_3256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3258 = 8'hb1 == _match_key_qbytes_1_T ? phv_data_177 : _GEN_3257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3259 = 8'hb2 == _match_key_qbytes_1_T ? phv_data_178 : _GEN_3258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3260 = 8'hb3 == _match_key_qbytes_1_T ? phv_data_179 : _GEN_3259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3261 = 8'hb4 == _match_key_qbytes_1_T ? phv_data_180 : _GEN_3260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3262 = 8'hb5 == _match_key_qbytes_1_T ? phv_data_181 : _GEN_3261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3263 = 8'hb6 == _match_key_qbytes_1_T ? phv_data_182 : _GEN_3262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3264 = 8'hb7 == _match_key_qbytes_1_T ? phv_data_183 : _GEN_3263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3265 = 8'hb8 == _match_key_qbytes_1_T ? phv_data_184 : _GEN_3264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3266 = 8'hb9 == _match_key_qbytes_1_T ? phv_data_185 : _GEN_3265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3267 = 8'hba == _match_key_qbytes_1_T ? phv_data_186 : _GEN_3266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3268 = 8'hbb == _match_key_qbytes_1_T ? phv_data_187 : _GEN_3267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3269 = 8'hbc == _match_key_qbytes_1_T ? phv_data_188 : _GEN_3268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3270 = 8'hbd == _match_key_qbytes_1_T ? phv_data_189 : _GEN_3269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3271 = 8'hbe == _match_key_qbytes_1_T ? phv_data_190 : _GEN_3270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3272 = 8'hbf == _match_key_qbytes_1_T ? phv_data_191 : _GEN_3271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3273 = 8'hc0 == _match_key_qbytes_1_T ? phv_data_192 : _GEN_3272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3274 = 8'hc1 == _match_key_qbytes_1_T ? phv_data_193 : _GEN_3273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3275 = 8'hc2 == _match_key_qbytes_1_T ? phv_data_194 : _GEN_3274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3276 = 8'hc3 == _match_key_qbytes_1_T ? phv_data_195 : _GEN_3275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3277 = 8'hc4 == _match_key_qbytes_1_T ? phv_data_196 : _GEN_3276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3278 = 8'hc5 == _match_key_qbytes_1_T ? phv_data_197 : _GEN_3277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3279 = 8'hc6 == _match_key_qbytes_1_T ? phv_data_198 : _GEN_3278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3280 = 8'hc7 == _match_key_qbytes_1_T ? phv_data_199 : _GEN_3279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3281 = 8'hc8 == _match_key_qbytes_1_T ? phv_data_200 : _GEN_3280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3282 = 8'hc9 == _match_key_qbytes_1_T ? phv_data_201 : _GEN_3281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3283 = 8'hca == _match_key_qbytes_1_T ? phv_data_202 : _GEN_3282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3284 = 8'hcb == _match_key_qbytes_1_T ? phv_data_203 : _GEN_3283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3285 = 8'hcc == _match_key_qbytes_1_T ? phv_data_204 : _GEN_3284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3286 = 8'hcd == _match_key_qbytes_1_T ? phv_data_205 : _GEN_3285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3287 = 8'hce == _match_key_qbytes_1_T ? phv_data_206 : _GEN_3286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3288 = 8'hcf == _match_key_qbytes_1_T ? phv_data_207 : _GEN_3287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3289 = 8'hd0 == _match_key_qbytes_1_T ? phv_data_208 : _GEN_3288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3290 = 8'hd1 == _match_key_qbytes_1_T ? phv_data_209 : _GEN_3289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3291 = 8'hd2 == _match_key_qbytes_1_T ? phv_data_210 : _GEN_3290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3292 = 8'hd3 == _match_key_qbytes_1_T ? phv_data_211 : _GEN_3291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3293 = 8'hd4 == _match_key_qbytes_1_T ? phv_data_212 : _GEN_3292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3294 = 8'hd5 == _match_key_qbytes_1_T ? phv_data_213 : _GEN_3293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3295 = 8'hd6 == _match_key_qbytes_1_T ? phv_data_214 : _GEN_3294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3296 = 8'hd7 == _match_key_qbytes_1_T ? phv_data_215 : _GEN_3295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3297 = 8'hd8 == _match_key_qbytes_1_T ? phv_data_216 : _GEN_3296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3298 = 8'hd9 == _match_key_qbytes_1_T ? phv_data_217 : _GEN_3297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3299 = 8'hda == _match_key_qbytes_1_T ? phv_data_218 : _GEN_3298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3300 = 8'hdb == _match_key_qbytes_1_T ? phv_data_219 : _GEN_3299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3301 = 8'hdc == _match_key_qbytes_1_T ? phv_data_220 : _GEN_3300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3302 = 8'hdd == _match_key_qbytes_1_T ? phv_data_221 : _GEN_3301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3303 = 8'hde == _match_key_qbytes_1_T ? phv_data_222 : _GEN_3302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3304 = 8'hdf == _match_key_qbytes_1_T ? phv_data_223 : _GEN_3303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3305 = 8'he0 == _match_key_qbytes_1_T ? phv_data_224 : _GEN_3304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3306 = 8'he1 == _match_key_qbytes_1_T ? phv_data_225 : _GEN_3305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3307 = 8'he2 == _match_key_qbytes_1_T ? phv_data_226 : _GEN_3306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3308 = 8'he3 == _match_key_qbytes_1_T ? phv_data_227 : _GEN_3307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3309 = 8'he4 == _match_key_qbytes_1_T ? phv_data_228 : _GEN_3308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3310 = 8'he5 == _match_key_qbytes_1_T ? phv_data_229 : _GEN_3309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3311 = 8'he6 == _match_key_qbytes_1_T ? phv_data_230 : _GEN_3310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3312 = 8'he7 == _match_key_qbytes_1_T ? phv_data_231 : _GEN_3311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3313 = 8'he8 == _match_key_qbytes_1_T ? phv_data_232 : _GEN_3312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3314 = 8'he9 == _match_key_qbytes_1_T ? phv_data_233 : _GEN_3313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3315 = 8'hea == _match_key_qbytes_1_T ? phv_data_234 : _GEN_3314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3316 = 8'heb == _match_key_qbytes_1_T ? phv_data_235 : _GEN_3315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3317 = 8'hec == _match_key_qbytes_1_T ? phv_data_236 : _GEN_3316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3318 = 8'hed == _match_key_qbytes_1_T ? phv_data_237 : _GEN_3317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3319 = 8'hee == _match_key_qbytes_1_T ? phv_data_238 : _GEN_3318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3320 = 8'hef == _match_key_qbytes_1_T ? phv_data_239 : _GEN_3319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3321 = 8'hf0 == _match_key_qbytes_1_T ? phv_data_240 : _GEN_3320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3322 = 8'hf1 == _match_key_qbytes_1_T ? phv_data_241 : _GEN_3321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3323 = 8'hf2 == _match_key_qbytes_1_T ? phv_data_242 : _GEN_3322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3324 = 8'hf3 == _match_key_qbytes_1_T ? phv_data_243 : _GEN_3323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3325 = 8'hf4 == _match_key_qbytes_1_T ? phv_data_244 : _GEN_3324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3326 = 8'hf5 == _match_key_qbytes_1_T ? phv_data_245 : _GEN_3325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3327 = 8'hf6 == _match_key_qbytes_1_T ? phv_data_246 : _GEN_3326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3328 = 8'hf7 == _match_key_qbytes_1_T ? phv_data_247 : _GEN_3327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3329 = 8'hf8 == _match_key_qbytes_1_T ? phv_data_248 : _GEN_3328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3330 = 8'hf9 == _match_key_qbytes_1_T ? phv_data_249 : _GEN_3329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3331 = 8'hfa == _match_key_qbytes_1_T ? phv_data_250 : _GEN_3330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3332 = 8'hfb == _match_key_qbytes_1_T ? phv_data_251 : _GEN_3331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3333 = 8'hfc == _match_key_qbytes_1_T ? phv_data_252 : _GEN_3332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3334 = 8'hfd == _match_key_qbytes_1_T ? phv_data_253 : _GEN_3333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3335 = 8'hfe == _match_key_qbytes_1_T ? phv_data_254 : _GEN_3334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3336 = 8'hff == _match_key_qbytes_1_T ? phv_data_255 : _GEN_3335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_13862 = {{1'd0}, _match_key_qbytes_1_T}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3337 = 9'h100 == _GEN_13862 ? phv_data_256 : _GEN_3336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3338 = 9'h101 == _GEN_13862 ? phv_data_257 : _GEN_3337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3339 = 9'h102 == _GEN_13862 ? phv_data_258 : _GEN_3338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3340 = 9'h103 == _GEN_13862 ? phv_data_259 : _GEN_3339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3341 = 9'h104 == _GEN_13862 ? phv_data_260 : _GEN_3340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3342 = 9'h105 == _GEN_13862 ? phv_data_261 : _GEN_3341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3343 = 9'h106 == _GEN_13862 ? phv_data_262 : _GEN_3342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3344 = 9'h107 == _GEN_13862 ? phv_data_263 : _GEN_3343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3345 = 9'h108 == _GEN_13862 ? phv_data_264 : _GEN_3344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3346 = 9'h109 == _GEN_13862 ? phv_data_265 : _GEN_3345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3347 = 9'h10a == _GEN_13862 ? phv_data_266 : _GEN_3346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3348 = 9'h10b == _GEN_13862 ? phv_data_267 : _GEN_3347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3349 = 9'h10c == _GEN_13862 ? phv_data_268 : _GEN_3348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3350 = 9'h10d == _GEN_13862 ? phv_data_269 : _GEN_3349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3351 = 9'h10e == _GEN_13862 ? phv_data_270 : _GEN_3350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3352 = 9'h10f == _GEN_13862 ? phv_data_271 : _GEN_3351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3353 = 9'h110 == _GEN_13862 ? phv_data_272 : _GEN_3352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3354 = 9'h111 == _GEN_13862 ? phv_data_273 : _GEN_3353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3355 = 9'h112 == _GEN_13862 ? phv_data_274 : _GEN_3354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3356 = 9'h113 == _GEN_13862 ? phv_data_275 : _GEN_3355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3357 = 9'h114 == _GEN_13862 ? phv_data_276 : _GEN_3356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3358 = 9'h115 == _GEN_13862 ? phv_data_277 : _GEN_3357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3359 = 9'h116 == _GEN_13862 ? phv_data_278 : _GEN_3358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3360 = 9'h117 == _GEN_13862 ? phv_data_279 : _GEN_3359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3361 = 9'h118 == _GEN_13862 ? phv_data_280 : _GEN_3360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3362 = 9'h119 == _GEN_13862 ? phv_data_281 : _GEN_3361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3363 = 9'h11a == _GEN_13862 ? phv_data_282 : _GEN_3362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3364 = 9'h11b == _GEN_13862 ? phv_data_283 : _GEN_3363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3365 = 9'h11c == _GEN_13862 ? phv_data_284 : _GEN_3364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3366 = 9'h11d == _GEN_13862 ? phv_data_285 : _GEN_3365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3367 = 9'h11e == _GEN_13862 ? phv_data_286 : _GEN_3366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3368 = 9'h11f == _GEN_13862 ? phv_data_287 : _GEN_3367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3369 = 9'h120 == _GEN_13862 ? phv_data_288 : _GEN_3368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3370 = 9'h121 == _GEN_13862 ? phv_data_289 : _GEN_3369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3371 = 9'h122 == _GEN_13862 ? phv_data_290 : _GEN_3370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3372 = 9'h123 == _GEN_13862 ? phv_data_291 : _GEN_3371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3373 = 9'h124 == _GEN_13862 ? phv_data_292 : _GEN_3372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3374 = 9'h125 == _GEN_13862 ? phv_data_293 : _GEN_3373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3375 = 9'h126 == _GEN_13862 ? phv_data_294 : _GEN_3374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3376 = 9'h127 == _GEN_13862 ? phv_data_295 : _GEN_3375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3377 = 9'h128 == _GEN_13862 ? phv_data_296 : _GEN_3376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3378 = 9'h129 == _GEN_13862 ? phv_data_297 : _GEN_3377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3379 = 9'h12a == _GEN_13862 ? phv_data_298 : _GEN_3378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3380 = 9'h12b == _GEN_13862 ? phv_data_299 : _GEN_3379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3381 = 9'h12c == _GEN_13862 ? phv_data_300 : _GEN_3380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3382 = 9'h12d == _GEN_13862 ? phv_data_301 : _GEN_3381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3383 = 9'h12e == _GEN_13862 ? phv_data_302 : _GEN_3382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3384 = 9'h12f == _GEN_13862 ? phv_data_303 : _GEN_3383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3385 = 9'h130 == _GEN_13862 ? phv_data_304 : _GEN_3384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3386 = 9'h131 == _GEN_13862 ? phv_data_305 : _GEN_3385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3387 = 9'h132 == _GEN_13862 ? phv_data_306 : _GEN_3386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3388 = 9'h133 == _GEN_13862 ? phv_data_307 : _GEN_3387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3389 = 9'h134 == _GEN_13862 ? phv_data_308 : _GEN_3388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3390 = 9'h135 == _GEN_13862 ? phv_data_309 : _GEN_3389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3391 = 9'h136 == _GEN_13862 ? phv_data_310 : _GEN_3390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3392 = 9'h137 == _GEN_13862 ? phv_data_311 : _GEN_3391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3393 = 9'h138 == _GEN_13862 ? phv_data_312 : _GEN_3392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3394 = 9'h139 == _GEN_13862 ? phv_data_313 : _GEN_3393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3395 = 9'h13a == _GEN_13862 ? phv_data_314 : _GEN_3394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3396 = 9'h13b == _GEN_13862 ? phv_data_315 : _GEN_3395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3397 = 9'h13c == _GEN_13862 ? phv_data_316 : _GEN_3396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3398 = 9'h13d == _GEN_13862 ? phv_data_317 : _GEN_3397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3399 = 9'h13e == _GEN_13862 ? phv_data_318 : _GEN_3398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3400 = 9'h13f == _GEN_13862 ? phv_data_319 : _GEN_3399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3401 = 9'h140 == _GEN_13862 ? phv_data_320 : _GEN_3400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3402 = 9'h141 == _GEN_13862 ? phv_data_321 : _GEN_3401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3403 = 9'h142 == _GEN_13862 ? phv_data_322 : _GEN_3402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3404 = 9'h143 == _GEN_13862 ? phv_data_323 : _GEN_3403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3405 = 9'h144 == _GEN_13862 ? phv_data_324 : _GEN_3404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3406 = 9'h145 == _GEN_13862 ? phv_data_325 : _GEN_3405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3407 = 9'h146 == _GEN_13862 ? phv_data_326 : _GEN_3406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3408 = 9'h147 == _GEN_13862 ? phv_data_327 : _GEN_3407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3409 = 9'h148 == _GEN_13862 ? phv_data_328 : _GEN_3408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3410 = 9'h149 == _GEN_13862 ? phv_data_329 : _GEN_3409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3411 = 9'h14a == _GEN_13862 ? phv_data_330 : _GEN_3410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3412 = 9'h14b == _GEN_13862 ? phv_data_331 : _GEN_3411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3413 = 9'h14c == _GEN_13862 ? phv_data_332 : _GEN_3412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3414 = 9'h14d == _GEN_13862 ? phv_data_333 : _GEN_3413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3415 = 9'h14e == _GEN_13862 ? phv_data_334 : _GEN_3414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3416 = 9'h14f == _GEN_13862 ? phv_data_335 : _GEN_3415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3417 = 9'h150 == _GEN_13862 ? phv_data_336 : _GEN_3416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3418 = 9'h151 == _GEN_13862 ? phv_data_337 : _GEN_3417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3419 = 9'h152 == _GEN_13862 ? phv_data_338 : _GEN_3418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3420 = 9'h153 == _GEN_13862 ? phv_data_339 : _GEN_3419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3421 = 9'h154 == _GEN_13862 ? phv_data_340 : _GEN_3420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3422 = 9'h155 == _GEN_13862 ? phv_data_341 : _GEN_3421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3423 = 9'h156 == _GEN_13862 ? phv_data_342 : _GEN_3422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3424 = 9'h157 == _GEN_13862 ? phv_data_343 : _GEN_3423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3425 = 9'h158 == _GEN_13862 ? phv_data_344 : _GEN_3424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3426 = 9'h159 == _GEN_13862 ? phv_data_345 : _GEN_3425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3427 = 9'h15a == _GEN_13862 ? phv_data_346 : _GEN_3426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3428 = 9'h15b == _GEN_13862 ? phv_data_347 : _GEN_3427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3429 = 9'h15c == _GEN_13862 ? phv_data_348 : _GEN_3428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3430 = 9'h15d == _GEN_13862 ? phv_data_349 : _GEN_3429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3431 = 9'h15e == _GEN_13862 ? phv_data_350 : _GEN_3430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3432 = 9'h15f == _GEN_13862 ? phv_data_351 : _GEN_3431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3433 = 9'h160 == _GEN_13862 ? phv_data_352 : _GEN_3432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3434 = 9'h161 == _GEN_13862 ? phv_data_353 : _GEN_3433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3435 = 9'h162 == _GEN_13862 ? phv_data_354 : _GEN_3434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3436 = 9'h163 == _GEN_13862 ? phv_data_355 : _GEN_3435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3437 = 9'h164 == _GEN_13862 ? phv_data_356 : _GEN_3436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3438 = 9'h165 == _GEN_13862 ? phv_data_357 : _GEN_3437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3439 = 9'h166 == _GEN_13862 ? phv_data_358 : _GEN_3438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3440 = 9'h167 == _GEN_13862 ? phv_data_359 : _GEN_3439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3441 = 9'h168 == _GEN_13862 ? phv_data_360 : _GEN_3440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3442 = 9'h169 == _GEN_13862 ? phv_data_361 : _GEN_3441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3443 = 9'h16a == _GEN_13862 ? phv_data_362 : _GEN_3442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3444 = 9'h16b == _GEN_13862 ? phv_data_363 : _GEN_3443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3445 = 9'h16c == _GEN_13862 ? phv_data_364 : _GEN_3444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3446 = 9'h16d == _GEN_13862 ? phv_data_365 : _GEN_3445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3447 = 9'h16e == _GEN_13862 ? phv_data_366 : _GEN_3446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3448 = 9'h16f == _GEN_13862 ? phv_data_367 : _GEN_3447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3449 = 9'h170 == _GEN_13862 ? phv_data_368 : _GEN_3448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3450 = 9'h171 == _GEN_13862 ? phv_data_369 : _GEN_3449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3451 = 9'h172 == _GEN_13862 ? phv_data_370 : _GEN_3450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3452 = 9'h173 == _GEN_13862 ? phv_data_371 : _GEN_3451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3453 = 9'h174 == _GEN_13862 ? phv_data_372 : _GEN_3452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3454 = 9'h175 == _GEN_13862 ? phv_data_373 : _GEN_3453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3455 = 9'h176 == _GEN_13862 ? phv_data_374 : _GEN_3454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3456 = 9'h177 == _GEN_13862 ? phv_data_375 : _GEN_3455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3457 = 9'h178 == _GEN_13862 ? phv_data_376 : _GEN_3456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3458 = 9'h179 == _GEN_13862 ? phv_data_377 : _GEN_3457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3459 = 9'h17a == _GEN_13862 ? phv_data_378 : _GEN_3458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3460 = 9'h17b == _GEN_13862 ? phv_data_379 : _GEN_3459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3461 = 9'h17c == _GEN_13862 ? phv_data_380 : _GEN_3460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3462 = 9'h17d == _GEN_13862 ? phv_data_381 : _GEN_3461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3463 = 9'h17e == _GEN_13862 ? phv_data_382 : _GEN_3462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3464 = 9'h17f == _GEN_13862 ? phv_data_383 : _GEN_3463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3465 = 9'h180 == _GEN_13862 ? phv_data_384 : _GEN_3464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3466 = 9'h181 == _GEN_13862 ? phv_data_385 : _GEN_3465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3467 = 9'h182 == _GEN_13862 ? phv_data_386 : _GEN_3466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3468 = 9'h183 == _GEN_13862 ? phv_data_387 : _GEN_3467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3469 = 9'h184 == _GEN_13862 ? phv_data_388 : _GEN_3468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3470 = 9'h185 == _GEN_13862 ? phv_data_389 : _GEN_3469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3471 = 9'h186 == _GEN_13862 ? phv_data_390 : _GEN_3470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3472 = 9'h187 == _GEN_13862 ? phv_data_391 : _GEN_3471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3473 = 9'h188 == _GEN_13862 ? phv_data_392 : _GEN_3472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3474 = 9'h189 == _GEN_13862 ? phv_data_393 : _GEN_3473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3475 = 9'h18a == _GEN_13862 ? phv_data_394 : _GEN_3474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3476 = 9'h18b == _GEN_13862 ? phv_data_395 : _GEN_3475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3477 = 9'h18c == _GEN_13862 ? phv_data_396 : _GEN_3476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3478 = 9'h18d == _GEN_13862 ? phv_data_397 : _GEN_3477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3479 = 9'h18e == _GEN_13862 ? phv_data_398 : _GEN_3478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3480 = 9'h18f == _GEN_13862 ? phv_data_399 : _GEN_3479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3481 = 9'h190 == _GEN_13862 ? phv_data_400 : _GEN_3480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3482 = 9'h191 == _GEN_13862 ? phv_data_401 : _GEN_3481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3483 = 9'h192 == _GEN_13862 ? phv_data_402 : _GEN_3482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3484 = 9'h193 == _GEN_13862 ? phv_data_403 : _GEN_3483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3485 = 9'h194 == _GEN_13862 ? phv_data_404 : _GEN_3484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3486 = 9'h195 == _GEN_13862 ? phv_data_405 : _GEN_3485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3487 = 9'h196 == _GEN_13862 ? phv_data_406 : _GEN_3486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3488 = 9'h197 == _GEN_13862 ? phv_data_407 : _GEN_3487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3489 = 9'h198 == _GEN_13862 ? phv_data_408 : _GEN_3488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3490 = 9'h199 == _GEN_13862 ? phv_data_409 : _GEN_3489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3491 = 9'h19a == _GEN_13862 ? phv_data_410 : _GEN_3490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3492 = 9'h19b == _GEN_13862 ? phv_data_411 : _GEN_3491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3493 = 9'h19c == _GEN_13862 ? phv_data_412 : _GEN_3492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3494 = 9'h19d == _GEN_13862 ? phv_data_413 : _GEN_3493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3495 = 9'h19e == _GEN_13862 ? phv_data_414 : _GEN_3494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3496 = 9'h19f == _GEN_13862 ? phv_data_415 : _GEN_3495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3497 = 9'h1a0 == _GEN_13862 ? phv_data_416 : _GEN_3496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3498 = 9'h1a1 == _GEN_13862 ? phv_data_417 : _GEN_3497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3499 = 9'h1a2 == _GEN_13862 ? phv_data_418 : _GEN_3498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3500 = 9'h1a3 == _GEN_13862 ? phv_data_419 : _GEN_3499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3501 = 9'h1a4 == _GEN_13862 ? phv_data_420 : _GEN_3500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3502 = 9'h1a5 == _GEN_13862 ? phv_data_421 : _GEN_3501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3503 = 9'h1a6 == _GEN_13862 ? phv_data_422 : _GEN_3502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3504 = 9'h1a7 == _GEN_13862 ? phv_data_423 : _GEN_3503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3505 = 9'h1a8 == _GEN_13862 ? phv_data_424 : _GEN_3504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3506 = 9'h1a9 == _GEN_13862 ? phv_data_425 : _GEN_3505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3507 = 9'h1aa == _GEN_13862 ? phv_data_426 : _GEN_3506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3508 = 9'h1ab == _GEN_13862 ? phv_data_427 : _GEN_3507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3509 = 9'h1ac == _GEN_13862 ? phv_data_428 : _GEN_3508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3510 = 9'h1ad == _GEN_13862 ? phv_data_429 : _GEN_3509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3511 = 9'h1ae == _GEN_13862 ? phv_data_430 : _GEN_3510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3512 = 9'h1af == _GEN_13862 ? phv_data_431 : _GEN_3511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3513 = 9'h1b0 == _GEN_13862 ? phv_data_432 : _GEN_3512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3514 = 9'h1b1 == _GEN_13862 ? phv_data_433 : _GEN_3513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3515 = 9'h1b2 == _GEN_13862 ? phv_data_434 : _GEN_3514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3516 = 9'h1b3 == _GEN_13862 ? phv_data_435 : _GEN_3515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3517 = 9'h1b4 == _GEN_13862 ? phv_data_436 : _GEN_3516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3518 = 9'h1b5 == _GEN_13862 ? phv_data_437 : _GEN_3517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3519 = 9'h1b6 == _GEN_13862 ? phv_data_438 : _GEN_3518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3520 = 9'h1b7 == _GEN_13862 ? phv_data_439 : _GEN_3519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3521 = 9'h1b8 == _GEN_13862 ? phv_data_440 : _GEN_3520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3522 = 9'h1b9 == _GEN_13862 ? phv_data_441 : _GEN_3521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3523 = 9'h1ba == _GEN_13862 ? phv_data_442 : _GEN_3522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3524 = 9'h1bb == _GEN_13862 ? phv_data_443 : _GEN_3523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3525 = 9'h1bc == _GEN_13862 ? phv_data_444 : _GEN_3524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3526 = 9'h1bd == _GEN_13862 ? phv_data_445 : _GEN_3525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3527 = 9'h1be == _GEN_13862 ? phv_data_446 : _GEN_3526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3528 = 9'h1bf == _GEN_13862 ? phv_data_447 : _GEN_3527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3529 = 9'h1c0 == _GEN_13862 ? phv_data_448 : _GEN_3528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3530 = 9'h1c1 == _GEN_13862 ? phv_data_449 : _GEN_3529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3531 = 9'h1c2 == _GEN_13862 ? phv_data_450 : _GEN_3530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3532 = 9'h1c3 == _GEN_13862 ? phv_data_451 : _GEN_3531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3533 = 9'h1c4 == _GEN_13862 ? phv_data_452 : _GEN_3532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3534 = 9'h1c5 == _GEN_13862 ? phv_data_453 : _GEN_3533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3535 = 9'h1c6 == _GEN_13862 ? phv_data_454 : _GEN_3534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3536 = 9'h1c7 == _GEN_13862 ? phv_data_455 : _GEN_3535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3537 = 9'h1c8 == _GEN_13862 ? phv_data_456 : _GEN_3536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3538 = 9'h1c9 == _GEN_13862 ? phv_data_457 : _GEN_3537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3539 = 9'h1ca == _GEN_13862 ? phv_data_458 : _GEN_3538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3540 = 9'h1cb == _GEN_13862 ? phv_data_459 : _GEN_3539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3541 = 9'h1cc == _GEN_13862 ? phv_data_460 : _GEN_3540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3542 = 9'h1cd == _GEN_13862 ? phv_data_461 : _GEN_3541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3543 = 9'h1ce == _GEN_13862 ? phv_data_462 : _GEN_3542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3544 = 9'h1cf == _GEN_13862 ? phv_data_463 : _GEN_3543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3545 = 9'h1d0 == _GEN_13862 ? phv_data_464 : _GEN_3544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3546 = 9'h1d1 == _GEN_13862 ? phv_data_465 : _GEN_3545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3547 = 9'h1d2 == _GEN_13862 ? phv_data_466 : _GEN_3546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3548 = 9'h1d3 == _GEN_13862 ? phv_data_467 : _GEN_3547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3549 = 9'h1d4 == _GEN_13862 ? phv_data_468 : _GEN_3548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3550 = 9'h1d5 == _GEN_13862 ? phv_data_469 : _GEN_3549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3551 = 9'h1d6 == _GEN_13862 ? phv_data_470 : _GEN_3550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3552 = 9'h1d7 == _GEN_13862 ? phv_data_471 : _GEN_3551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3553 = 9'h1d8 == _GEN_13862 ? phv_data_472 : _GEN_3552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3554 = 9'h1d9 == _GEN_13862 ? phv_data_473 : _GEN_3553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3555 = 9'h1da == _GEN_13862 ? phv_data_474 : _GEN_3554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3556 = 9'h1db == _GEN_13862 ? phv_data_475 : _GEN_3555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3557 = 9'h1dc == _GEN_13862 ? phv_data_476 : _GEN_3556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3558 = 9'h1dd == _GEN_13862 ? phv_data_477 : _GEN_3557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3559 = 9'h1de == _GEN_13862 ? phv_data_478 : _GEN_3558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3560 = 9'h1df == _GEN_13862 ? phv_data_479 : _GEN_3559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3561 = 9'h1e0 == _GEN_13862 ? phv_data_480 : _GEN_3560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3562 = 9'h1e1 == _GEN_13862 ? phv_data_481 : _GEN_3561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3563 = 9'h1e2 == _GEN_13862 ? phv_data_482 : _GEN_3562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3564 = 9'h1e3 == _GEN_13862 ? phv_data_483 : _GEN_3563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3565 = 9'h1e4 == _GEN_13862 ? phv_data_484 : _GEN_3564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3566 = 9'h1e5 == _GEN_13862 ? phv_data_485 : _GEN_3565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3567 = 9'h1e6 == _GEN_13862 ? phv_data_486 : _GEN_3566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3568 = 9'h1e7 == _GEN_13862 ? phv_data_487 : _GEN_3567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3569 = 9'h1e8 == _GEN_13862 ? phv_data_488 : _GEN_3568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3570 = 9'h1e9 == _GEN_13862 ? phv_data_489 : _GEN_3569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3571 = 9'h1ea == _GEN_13862 ? phv_data_490 : _GEN_3570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3572 = 9'h1eb == _GEN_13862 ? phv_data_491 : _GEN_3571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3573 = 9'h1ec == _GEN_13862 ? phv_data_492 : _GEN_3572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3574 = 9'h1ed == _GEN_13862 ? phv_data_493 : _GEN_3573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3575 = 9'h1ee == _GEN_13862 ? phv_data_494 : _GEN_3574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3576 = 9'h1ef == _GEN_13862 ? phv_data_495 : _GEN_3575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3577 = 9'h1f0 == _GEN_13862 ? phv_data_496 : _GEN_3576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3578 = 9'h1f1 == _GEN_13862 ? phv_data_497 : _GEN_3577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3579 = 9'h1f2 == _GEN_13862 ? phv_data_498 : _GEN_3578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3580 = 9'h1f3 == _GEN_13862 ? phv_data_499 : _GEN_3579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3581 = 9'h1f4 == _GEN_13862 ? phv_data_500 : _GEN_3580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3582 = 9'h1f5 == _GEN_13862 ? phv_data_501 : _GEN_3581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3583 = 9'h1f6 == _GEN_13862 ? phv_data_502 : _GEN_3582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3584 = 9'h1f7 == _GEN_13862 ? phv_data_503 : _GEN_3583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3585 = 9'h1f8 == _GEN_13862 ? phv_data_504 : _GEN_3584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3586 = 9'h1f9 == _GEN_13862 ? phv_data_505 : _GEN_3585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3587 = 9'h1fa == _GEN_13862 ? phv_data_506 : _GEN_3586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3588 = 9'h1fb == _GEN_13862 ? phv_data_507 : _GEN_3587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3589 = 9'h1fc == _GEN_13862 ? phv_data_508 : _GEN_3588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3590 = 9'h1fd == _GEN_13862 ? phv_data_509 : _GEN_3589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3591 = 9'h1fe == _GEN_13862 ? phv_data_510 : _GEN_3590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3592 = 9'h1ff == _GEN_13862 ? phv_data_511 : _GEN_3591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3594 = 8'h1 == _match_key_qbytes_1_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3595 = 8'h2 == _match_key_qbytes_1_T_1 ? phv_data_2 : _GEN_3594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3596 = 8'h3 == _match_key_qbytes_1_T_1 ? phv_data_3 : _GEN_3595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3597 = 8'h4 == _match_key_qbytes_1_T_1 ? phv_data_4 : _GEN_3596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3598 = 8'h5 == _match_key_qbytes_1_T_1 ? phv_data_5 : _GEN_3597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3599 = 8'h6 == _match_key_qbytes_1_T_1 ? phv_data_6 : _GEN_3598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3600 = 8'h7 == _match_key_qbytes_1_T_1 ? phv_data_7 : _GEN_3599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3601 = 8'h8 == _match_key_qbytes_1_T_1 ? phv_data_8 : _GEN_3600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3602 = 8'h9 == _match_key_qbytes_1_T_1 ? phv_data_9 : _GEN_3601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3603 = 8'ha == _match_key_qbytes_1_T_1 ? phv_data_10 : _GEN_3602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3604 = 8'hb == _match_key_qbytes_1_T_1 ? phv_data_11 : _GEN_3603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3605 = 8'hc == _match_key_qbytes_1_T_1 ? phv_data_12 : _GEN_3604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3606 = 8'hd == _match_key_qbytes_1_T_1 ? phv_data_13 : _GEN_3605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3607 = 8'he == _match_key_qbytes_1_T_1 ? phv_data_14 : _GEN_3606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3608 = 8'hf == _match_key_qbytes_1_T_1 ? phv_data_15 : _GEN_3607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3609 = 8'h10 == _match_key_qbytes_1_T_1 ? phv_data_16 : _GEN_3608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3610 = 8'h11 == _match_key_qbytes_1_T_1 ? phv_data_17 : _GEN_3609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3611 = 8'h12 == _match_key_qbytes_1_T_1 ? phv_data_18 : _GEN_3610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3612 = 8'h13 == _match_key_qbytes_1_T_1 ? phv_data_19 : _GEN_3611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3613 = 8'h14 == _match_key_qbytes_1_T_1 ? phv_data_20 : _GEN_3612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3614 = 8'h15 == _match_key_qbytes_1_T_1 ? phv_data_21 : _GEN_3613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3615 = 8'h16 == _match_key_qbytes_1_T_1 ? phv_data_22 : _GEN_3614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3616 = 8'h17 == _match_key_qbytes_1_T_1 ? phv_data_23 : _GEN_3615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3617 = 8'h18 == _match_key_qbytes_1_T_1 ? phv_data_24 : _GEN_3616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3618 = 8'h19 == _match_key_qbytes_1_T_1 ? phv_data_25 : _GEN_3617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3619 = 8'h1a == _match_key_qbytes_1_T_1 ? phv_data_26 : _GEN_3618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3620 = 8'h1b == _match_key_qbytes_1_T_1 ? phv_data_27 : _GEN_3619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3621 = 8'h1c == _match_key_qbytes_1_T_1 ? phv_data_28 : _GEN_3620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3622 = 8'h1d == _match_key_qbytes_1_T_1 ? phv_data_29 : _GEN_3621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3623 = 8'h1e == _match_key_qbytes_1_T_1 ? phv_data_30 : _GEN_3622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3624 = 8'h1f == _match_key_qbytes_1_T_1 ? phv_data_31 : _GEN_3623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3625 = 8'h20 == _match_key_qbytes_1_T_1 ? phv_data_32 : _GEN_3624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3626 = 8'h21 == _match_key_qbytes_1_T_1 ? phv_data_33 : _GEN_3625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3627 = 8'h22 == _match_key_qbytes_1_T_1 ? phv_data_34 : _GEN_3626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3628 = 8'h23 == _match_key_qbytes_1_T_1 ? phv_data_35 : _GEN_3627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3629 = 8'h24 == _match_key_qbytes_1_T_1 ? phv_data_36 : _GEN_3628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3630 = 8'h25 == _match_key_qbytes_1_T_1 ? phv_data_37 : _GEN_3629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3631 = 8'h26 == _match_key_qbytes_1_T_1 ? phv_data_38 : _GEN_3630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3632 = 8'h27 == _match_key_qbytes_1_T_1 ? phv_data_39 : _GEN_3631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3633 = 8'h28 == _match_key_qbytes_1_T_1 ? phv_data_40 : _GEN_3632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3634 = 8'h29 == _match_key_qbytes_1_T_1 ? phv_data_41 : _GEN_3633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3635 = 8'h2a == _match_key_qbytes_1_T_1 ? phv_data_42 : _GEN_3634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3636 = 8'h2b == _match_key_qbytes_1_T_1 ? phv_data_43 : _GEN_3635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3637 = 8'h2c == _match_key_qbytes_1_T_1 ? phv_data_44 : _GEN_3636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3638 = 8'h2d == _match_key_qbytes_1_T_1 ? phv_data_45 : _GEN_3637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3639 = 8'h2e == _match_key_qbytes_1_T_1 ? phv_data_46 : _GEN_3638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3640 = 8'h2f == _match_key_qbytes_1_T_1 ? phv_data_47 : _GEN_3639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3641 = 8'h30 == _match_key_qbytes_1_T_1 ? phv_data_48 : _GEN_3640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3642 = 8'h31 == _match_key_qbytes_1_T_1 ? phv_data_49 : _GEN_3641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3643 = 8'h32 == _match_key_qbytes_1_T_1 ? phv_data_50 : _GEN_3642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3644 = 8'h33 == _match_key_qbytes_1_T_1 ? phv_data_51 : _GEN_3643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3645 = 8'h34 == _match_key_qbytes_1_T_1 ? phv_data_52 : _GEN_3644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3646 = 8'h35 == _match_key_qbytes_1_T_1 ? phv_data_53 : _GEN_3645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3647 = 8'h36 == _match_key_qbytes_1_T_1 ? phv_data_54 : _GEN_3646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3648 = 8'h37 == _match_key_qbytes_1_T_1 ? phv_data_55 : _GEN_3647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3649 = 8'h38 == _match_key_qbytes_1_T_1 ? phv_data_56 : _GEN_3648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3650 = 8'h39 == _match_key_qbytes_1_T_1 ? phv_data_57 : _GEN_3649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3651 = 8'h3a == _match_key_qbytes_1_T_1 ? phv_data_58 : _GEN_3650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3652 = 8'h3b == _match_key_qbytes_1_T_1 ? phv_data_59 : _GEN_3651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3653 = 8'h3c == _match_key_qbytes_1_T_1 ? phv_data_60 : _GEN_3652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3654 = 8'h3d == _match_key_qbytes_1_T_1 ? phv_data_61 : _GEN_3653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3655 = 8'h3e == _match_key_qbytes_1_T_1 ? phv_data_62 : _GEN_3654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3656 = 8'h3f == _match_key_qbytes_1_T_1 ? phv_data_63 : _GEN_3655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3657 = 8'h40 == _match_key_qbytes_1_T_1 ? phv_data_64 : _GEN_3656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3658 = 8'h41 == _match_key_qbytes_1_T_1 ? phv_data_65 : _GEN_3657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3659 = 8'h42 == _match_key_qbytes_1_T_1 ? phv_data_66 : _GEN_3658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3660 = 8'h43 == _match_key_qbytes_1_T_1 ? phv_data_67 : _GEN_3659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3661 = 8'h44 == _match_key_qbytes_1_T_1 ? phv_data_68 : _GEN_3660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3662 = 8'h45 == _match_key_qbytes_1_T_1 ? phv_data_69 : _GEN_3661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3663 = 8'h46 == _match_key_qbytes_1_T_1 ? phv_data_70 : _GEN_3662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3664 = 8'h47 == _match_key_qbytes_1_T_1 ? phv_data_71 : _GEN_3663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3665 = 8'h48 == _match_key_qbytes_1_T_1 ? phv_data_72 : _GEN_3664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3666 = 8'h49 == _match_key_qbytes_1_T_1 ? phv_data_73 : _GEN_3665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3667 = 8'h4a == _match_key_qbytes_1_T_1 ? phv_data_74 : _GEN_3666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3668 = 8'h4b == _match_key_qbytes_1_T_1 ? phv_data_75 : _GEN_3667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3669 = 8'h4c == _match_key_qbytes_1_T_1 ? phv_data_76 : _GEN_3668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3670 = 8'h4d == _match_key_qbytes_1_T_1 ? phv_data_77 : _GEN_3669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3671 = 8'h4e == _match_key_qbytes_1_T_1 ? phv_data_78 : _GEN_3670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3672 = 8'h4f == _match_key_qbytes_1_T_1 ? phv_data_79 : _GEN_3671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3673 = 8'h50 == _match_key_qbytes_1_T_1 ? phv_data_80 : _GEN_3672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3674 = 8'h51 == _match_key_qbytes_1_T_1 ? phv_data_81 : _GEN_3673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3675 = 8'h52 == _match_key_qbytes_1_T_1 ? phv_data_82 : _GEN_3674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3676 = 8'h53 == _match_key_qbytes_1_T_1 ? phv_data_83 : _GEN_3675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3677 = 8'h54 == _match_key_qbytes_1_T_1 ? phv_data_84 : _GEN_3676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3678 = 8'h55 == _match_key_qbytes_1_T_1 ? phv_data_85 : _GEN_3677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3679 = 8'h56 == _match_key_qbytes_1_T_1 ? phv_data_86 : _GEN_3678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3680 = 8'h57 == _match_key_qbytes_1_T_1 ? phv_data_87 : _GEN_3679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3681 = 8'h58 == _match_key_qbytes_1_T_1 ? phv_data_88 : _GEN_3680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3682 = 8'h59 == _match_key_qbytes_1_T_1 ? phv_data_89 : _GEN_3681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3683 = 8'h5a == _match_key_qbytes_1_T_1 ? phv_data_90 : _GEN_3682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3684 = 8'h5b == _match_key_qbytes_1_T_1 ? phv_data_91 : _GEN_3683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3685 = 8'h5c == _match_key_qbytes_1_T_1 ? phv_data_92 : _GEN_3684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3686 = 8'h5d == _match_key_qbytes_1_T_1 ? phv_data_93 : _GEN_3685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3687 = 8'h5e == _match_key_qbytes_1_T_1 ? phv_data_94 : _GEN_3686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3688 = 8'h5f == _match_key_qbytes_1_T_1 ? phv_data_95 : _GEN_3687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3689 = 8'h60 == _match_key_qbytes_1_T_1 ? phv_data_96 : _GEN_3688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3690 = 8'h61 == _match_key_qbytes_1_T_1 ? phv_data_97 : _GEN_3689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3691 = 8'h62 == _match_key_qbytes_1_T_1 ? phv_data_98 : _GEN_3690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3692 = 8'h63 == _match_key_qbytes_1_T_1 ? phv_data_99 : _GEN_3691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3693 = 8'h64 == _match_key_qbytes_1_T_1 ? phv_data_100 : _GEN_3692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3694 = 8'h65 == _match_key_qbytes_1_T_1 ? phv_data_101 : _GEN_3693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3695 = 8'h66 == _match_key_qbytes_1_T_1 ? phv_data_102 : _GEN_3694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3696 = 8'h67 == _match_key_qbytes_1_T_1 ? phv_data_103 : _GEN_3695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3697 = 8'h68 == _match_key_qbytes_1_T_1 ? phv_data_104 : _GEN_3696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3698 = 8'h69 == _match_key_qbytes_1_T_1 ? phv_data_105 : _GEN_3697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3699 = 8'h6a == _match_key_qbytes_1_T_1 ? phv_data_106 : _GEN_3698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3700 = 8'h6b == _match_key_qbytes_1_T_1 ? phv_data_107 : _GEN_3699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3701 = 8'h6c == _match_key_qbytes_1_T_1 ? phv_data_108 : _GEN_3700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3702 = 8'h6d == _match_key_qbytes_1_T_1 ? phv_data_109 : _GEN_3701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3703 = 8'h6e == _match_key_qbytes_1_T_1 ? phv_data_110 : _GEN_3702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3704 = 8'h6f == _match_key_qbytes_1_T_1 ? phv_data_111 : _GEN_3703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3705 = 8'h70 == _match_key_qbytes_1_T_1 ? phv_data_112 : _GEN_3704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3706 = 8'h71 == _match_key_qbytes_1_T_1 ? phv_data_113 : _GEN_3705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3707 = 8'h72 == _match_key_qbytes_1_T_1 ? phv_data_114 : _GEN_3706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3708 = 8'h73 == _match_key_qbytes_1_T_1 ? phv_data_115 : _GEN_3707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3709 = 8'h74 == _match_key_qbytes_1_T_1 ? phv_data_116 : _GEN_3708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3710 = 8'h75 == _match_key_qbytes_1_T_1 ? phv_data_117 : _GEN_3709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3711 = 8'h76 == _match_key_qbytes_1_T_1 ? phv_data_118 : _GEN_3710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3712 = 8'h77 == _match_key_qbytes_1_T_1 ? phv_data_119 : _GEN_3711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3713 = 8'h78 == _match_key_qbytes_1_T_1 ? phv_data_120 : _GEN_3712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3714 = 8'h79 == _match_key_qbytes_1_T_1 ? phv_data_121 : _GEN_3713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3715 = 8'h7a == _match_key_qbytes_1_T_1 ? phv_data_122 : _GEN_3714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3716 = 8'h7b == _match_key_qbytes_1_T_1 ? phv_data_123 : _GEN_3715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3717 = 8'h7c == _match_key_qbytes_1_T_1 ? phv_data_124 : _GEN_3716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3718 = 8'h7d == _match_key_qbytes_1_T_1 ? phv_data_125 : _GEN_3717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3719 = 8'h7e == _match_key_qbytes_1_T_1 ? phv_data_126 : _GEN_3718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3720 = 8'h7f == _match_key_qbytes_1_T_1 ? phv_data_127 : _GEN_3719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3721 = 8'h80 == _match_key_qbytes_1_T_1 ? phv_data_128 : _GEN_3720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3722 = 8'h81 == _match_key_qbytes_1_T_1 ? phv_data_129 : _GEN_3721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3723 = 8'h82 == _match_key_qbytes_1_T_1 ? phv_data_130 : _GEN_3722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3724 = 8'h83 == _match_key_qbytes_1_T_1 ? phv_data_131 : _GEN_3723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3725 = 8'h84 == _match_key_qbytes_1_T_1 ? phv_data_132 : _GEN_3724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3726 = 8'h85 == _match_key_qbytes_1_T_1 ? phv_data_133 : _GEN_3725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3727 = 8'h86 == _match_key_qbytes_1_T_1 ? phv_data_134 : _GEN_3726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3728 = 8'h87 == _match_key_qbytes_1_T_1 ? phv_data_135 : _GEN_3727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3729 = 8'h88 == _match_key_qbytes_1_T_1 ? phv_data_136 : _GEN_3728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3730 = 8'h89 == _match_key_qbytes_1_T_1 ? phv_data_137 : _GEN_3729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3731 = 8'h8a == _match_key_qbytes_1_T_1 ? phv_data_138 : _GEN_3730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3732 = 8'h8b == _match_key_qbytes_1_T_1 ? phv_data_139 : _GEN_3731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3733 = 8'h8c == _match_key_qbytes_1_T_1 ? phv_data_140 : _GEN_3732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3734 = 8'h8d == _match_key_qbytes_1_T_1 ? phv_data_141 : _GEN_3733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3735 = 8'h8e == _match_key_qbytes_1_T_1 ? phv_data_142 : _GEN_3734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3736 = 8'h8f == _match_key_qbytes_1_T_1 ? phv_data_143 : _GEN_3735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3737 = 8'h90 == _match_key_qbytes_1_T_1 ? phv_data_144 : _GEN_3736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3738 = 8'h91 == _match_key_qbytes_1_T_1 ? phv_data_145 : _GEN_3737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3739 = 8'h92 == _match_key_qbytes_1_T_1 ? phv_data_146 : _GEN_3738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3740 = 8'h93 == _match_key_qbytes_1_T_1 ? phv_data_147 : _GEN_3739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3741 = 8'h94 == _match_key_qbytes_1_T_1 ? phv_data_148 : _GEN_3740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3742 = 8'h95 == _match_key_qbytes_1_T_1 ? phv_data_149 : _GEN_3741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3743 = 8'h96 == _match_key_qbytes_1_T_1 ? phv_data_150 : _GEN_3742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3744 = 8'h97 == _match_key_qbytes_1_T_1 ? phv_data_151 : _GEN_3743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3745 = 8'h98 == _match_key_qbytes_1_T_1 ? phv_data_152 : _GEN_3744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3746 = 8'h99 == _match_key_qbytes_1_T_1 ? phv_data_153 : _GEN_3745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3747 = 8'h9a == _match_key_qbytes_1_T_1 ? phv_data_154 : _GEN_3746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3748 = 8'h9b == _match_key_qbytes_1_T_1 ? phv_data_155 : _GEN_3747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3749 = 8'h9c == _match_key_qbytes_1_T_1 ? phv_data_156 : _GEN_3748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3750 = 8'h9d == _match_key_qbytes_1_T_1 ? phv_data_157 : _GEN_3749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3751 = 8'h9e == _match_key_qbytes_1_T_1 ? phv_data_158 : _GEN_3750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3752 = 8'h9f == _match_key_qbytes_1_T_1 ? phv_data_159 : _GEN_3751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3753 = 8'ha0 == _match_key_qbytes_1_T_1 ? phv_data_160 : _GEN_3752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3754 = 8'ha1 == _match_key_qbytes_1_T_1 ? phv_data_161 : _GEN_3753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3755 = 8'ha2 == _match_key_qbytes_1_T_1 ? phv_data_162 : _GEN_3754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3756 = 8'ha3 == _match_key_qbytes_1_T_1 ? phv_data_163 : _GEN_3755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3757 = 8'ha4 == _match_key_qbytes_1_T_1 ? phv_data_164 : _GEN_3756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3758 = 8'ha5 == _match_key_qbytes_1_T_1 ? phv_data_165 : _GEN_3757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3759 = 8'ha6 == _match_key_qbytes_1_T_1 ? phv_data_166 : _GEN_3758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3760 = 8'ha7 == _match_key_qbytes_1_T_1 ? phv_data_167 : _GEN_3759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3761 = 8'ha8 == _match_key_qbytes_1_T_1 ? phv_data_168 : _GEN_3760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3762 = 8'ha9 == _match_key_qbytes_1_T_1 ? phv_data_169 : _GEN_3761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3763 = 8'haa == _match_key_qbytes_1_T_1 ? phv_data_170 : _GEN_3762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3764 = 8'hab == _match_key_qbytes_1_T_1 ? phv_data_171 : _GEN_3763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3765 = 8'hac == _match_key_qbytes_1_T_1 ? phv_data_172 : _GEN_3764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3766 = 8'had == _match_key_qbytes_1_T_1 ? phv_data_173 : _GEN_3765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3767 = 8'hae == _match_key_qbytes_1_T_1 ? phv_data_174 : _GEN_3766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3768 = 8'haf == _match_key_qbytes_1_T_1 ? phv_data_175 : _GEN_3767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3769 = 8'hb0 == _match_key_qbytes_1_T_1 ? phv_data_176 : _GEN_3768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3770 = 8'hb1 == _match_key_qbytes_1_T_1 ? phv_data_177 : _GEN_3769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3771 = 8'hb2 == _match_key_qbytes_1_T_1 ? phv_data_178 : _GEN_3770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3772 = 8'hb3 == _match_key_qbytes_1_T_1 ? phv_data_179 : _GEN_3771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3773 = 8'hb4 == _match_key_qbytes_1_T_1 ? phv_data_180 : _GEN_3772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3774 = 8'hb5 == _match_key_qbytes_1_T_1 ? phv_data_181 : _GEN_3773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3775 = 8'hb6 == _match_key_qbytes_1_T_1 ? phv_data_182 : _GEN_3774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3776 = 8'hb7 == _match_key_qbytes_1_T_1 ? phv_data_183 : _GEN_3775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3777 = 8'hb8 == _match_key_qbytes_1_T_1 ? phv_data_184 : _GEN_3776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3778 = 8'hb9 == _match_key_qbytes_1_T_1 ? phv_data_185 : _GEN_3777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3779 = 8'hba == _match_key_qbytes_1_T_1 ? phv_data_186 : _GEN_3778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3780 = 8'hbb == _match_key_qbytes_1_T_1 ? phv_data_187 : _GEN_3779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3781 = 8'hbc == _match_key_qbytes_1_T_1 ? phv_data_188 : _GEN_3780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3782 = 8'hbd == _match_key_qbytes_1_T_1 ? phv_data_189 : _GEN_3781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3783 = 8'hbe == _match_key_qbytes_1_T_1 ? phv_data_190 : _GEN_3782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3784 = 8'hbf == _match_key_qbytes_1_T_1 ? phv_data_191 : _GEN_3783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3785 = 8'hc0 == _match_key_qbytes_1_T_1 ? phv_data_192 : _GEN_3784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3786 = 8'hc1 == _match_key_qbytes_1_T_1 ? phv_data_193 : _GEN_3785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3787 = 8'hc2 == _match_key_qbytes_1_T_1 ? phv_data_194 : _GEN_3786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3788 = 8'hc3 == _match_key_qbytes_1_T_1 ? phv_data_195 : _GEN_3787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3789 = 8'hc4 == _match_key_qbytes_1_T_1 ? phv_data_196 : _GEN_3788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3790 = 8'hc5 == _match_key_qbytes_1_T_1 ? phv_data_197 : _GEN_3789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3791 = 8'hc6 == _match_key_qbytes_1_T_1 ? phv_data_198 : _GEN_3790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3792 = 8'hc7 == _match_key_qbytes_1_T_1 ? phv_data_199 : _GEN_3791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3793 = 8'hc8 == _match_key_qbytes_1_T_1 ? phv_data_200 : _GEN_3792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3794 = 8'hc9 == _match_key_qbytes_1_T_1 ? phv_data_201 : _GEN_3793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3795 = 8'hca == _match_key_qbytes_1_T_1 ? phv_data_202 : _GEN_3794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3796 = 8'hcb == _match_key_qbytes_1_T_1 ? phv_data_203 : _GEN_3795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3797 = 8'hcc == _match_key_qbytes_1_T_1 ? phv_data_204 : _GEN_3796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3798 = 8'hcd == _match_key_qbytes_1_T_1 ? phv_data_205 : _GEN_3797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3799 = 8'hce == _match_key_qbytes_1_T_1 ? phv_data_206 : _GEN_3798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3800 = 8'hcf == _match_key_qbytes_1_T_1 ? phv_data_207 : _GEN_3799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3801 = 8'hd0 == _match_key_qbytes_1_T_1 ? phv_data_208 : _GEN_3800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3802 = 8'hd1 == _match_key_qbytes_1_T_1 ? phv_data_209 : _GEN_3801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3803 = 8'hd2 == _match_key_qbytes_1_T_1 ? phv_data_210 : _GEN_3802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3804 = 8'hd3 == _match_key_qbytes_1_T_1 ? phv_data_211 : _GEN_3803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3805 = 8'hd4 == _match_key_qbytes_1_T_1 ? phv_data_212 : _GEN_3804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3806 = 8'hd5 == _match_key_qbytes_1_T_1 ? phv_data_213 : _GEN_3805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3807 = 8'hd6 == _match_key_qbytes_1_T_1 ? phv_data_214 : _GEN_3806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3808 = 8'hd7 == _match_key_qbytes_1_T_1 ? phv_data_215 : _GEN_3807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3809 = 8'hd8 == _match_key_qbytes_1_T_1 ? phv_data_216 : _GEN_3808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3810 = 8'hd9 == _match_key_qbytes_1_T_1 ? phv_data_217 : _GEN_3809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3811 = 8'hda == _match_key_qbytes_1_T_1 ? phv_data_218 : _GEN_3810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3812 = 8'hdb == _match_key_qbytes_1_T_1 ? phv_data_219 : _GEN_3811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3813 = 8'hdc == _match_key_qbytes_1_T_1 ? phv_data_220 : _GEN_3812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3814 = 8'hdd == _match_key_qbytes_1_T_1 ? phv_data_221 : _GEN_3813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3815 = 8'hde == _match_key_qbytes_1_T_1 ? phv_data_222 : _GEN_3814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3816 = 8'hdf == _match_key_qbytes_1_T_1 ? phv_data_223 : _GEN_3815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3817 = 8'he0 == _match_key_qbytes_1_T_1 ? phv_data_224 : _GEN_3816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3818 = 8'he1 == _match_key_qbytes_1_T_1 ? phv_data_225 : _GEN_3817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3819 = 8'he2 == _match_key_qbytes_1_T_1 ? phv_data_226 : _GEN_3818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3820 = 8'he3 == _match_key_qbytes_1_T_1 ? phv_data_227 : _GEN_3819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3821 = 8'he4 == _match_key_qbytes_1_T_1 ? phv_data_228 : _GEN_3820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3822 = 8'he5 == _match_key_qbytes_1_T_1 ? phv_data_229 : _GEN_3821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3823 = 8'he6 == _match_key_qbytes_1_T_1 ? phv_data_230 : _GEN_3822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3824 = 8'he7 == _match_key_qbytes_1_T_1 ? phv_data_231 : _GEN_3823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3825 = 8'he8 == _match_key_qbytes_1_T_1 ? phv_data_232 : _GEN_3824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3826 = 8'he9 == _match_key_qbytes_1_T_1 ? phv_data_233 : _GEN_3825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3827 = 8'hea == _match_key_qbytes_1_T_1 ? phv_data_234 : _GEN_3826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3828 = 8'heb == _match_key_qbytes_1_T_1 ? phv_data_235 : _GEN_3827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3829 = 8'hec == _match_key_qbytes_1_T_1 ? phv_data_236 : _GEN_3828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3830 = 8'hed == _match_key_qbytes_1_T_1 ? phv_data_237 : _GEN_3829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3831 = 8'hee == _match_key_qbytes_1_T_1 ? phv_data_238 : _GEN_3830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3832 = 8'hef == _match_key_qbytes_1_T_1 ? phv_data_239 : _GEN_3831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3833 = 8'hf0 == _match_key_qbytes_1_T_1 ? phv_data_240 : _GEN_3832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3834 = 8'hf1 == _match_key_qbytes_1_T_1 ? phv_data_241 : _GEN_3833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3835 = 8'hf2 == _match_key_qbytes_1_T_1 ? phv_data_242 : _GEN_3834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3836 = 8'hf3 == _match_key_qbytes_1_T_1 ? phv_data_243 : _GEN_3835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3837 = 8'hf4 == _match_key_qbytes_1_T_1 ? phv_data_244 : _GEN_3836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3838 = 8'hf5 == _match_key_qbytes_1_T_1 ? phv_data_245 : _GEN_3837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3839 = 8'hf6 == _match_key_qbytes_1_T_1 ? phv_data_246 : _GEN_3838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3840 = 8'hf7 == _match_key_qbytes_1_T_1 ? phv_data_247 : _GEN_3839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3841 = 8'hf8 == _match_key_qbytes_1_T_1 ? phv_data_248 : _GEN_3840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3842 = 8'hf9 == _match_key_qbytes_1_T_1 ? phv_data_249 : _GEN_3841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3843 = 8'hfa == _match_key_qbytes_1_T_1 ? phv_data_250 : _GEN_3842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3844 = 8'hfb == _match_key_qbytes_1_T_1 ? phv_data_251 : _GEN_3843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3845 = 8'hfc == _match_key_qbytes_1_T_1 ? phv_data_252 : _GEN_3844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3846 = 8'hfd == _match_key_qbytes_1_T_1 ? phv_data_253 : _GEN_3845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3847 = 8'hfe == _match_key_qbytes_1_T_1 ? phv_data_254 : _GEN_3846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3848 = 8'hff == _match_key_qbytes_1_T_1 ? phv_data_255 : _GEN_3847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_14118 = {{1'd0}, _match_key_qbytes_1_T_1}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3849 = 9'h100 == _GEN_14118 ? phv_data_256 : _GEN_3848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3850 = 9'h101 == _GEN_14118 ? phv_data_257 : _GEN_3849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3851 = 9'h102 == _GEN_14118 ? phv_data_258 : _GEN_3850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3852 = 9'h103 == _GEN_14118 ? phv_data_259 : _GEN_3851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3853 = 9'h104 == _GEN_14118 ? phv_data_260 : _GEN_3852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3854 = 9'h105 == _GEN_14118 ? phv_data_261 : _GEN_3853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3855 = 9'h106 == _GEN_14118 ? phv_data_262 : _GEN_3854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3856 = 9'h107 == _GEN_14118 ? phv_data_263 : _GEN_3855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3857 = 9'h108 == _GEN_14118 ? phv_data_264 : _GEN_3856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3858 = 9'h109 == _GEN_14118 ? phv_data_265 : _GEN_3857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3859 = 9'h10a == _GEN_14118 ? phv_data_266 : _GEN_3858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3860 = 9'h10b == _GEN_14118 ? phv_data_267 : _GEN_3859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3861 = 9'h10c == _GEN_14118 ? phv_data_268 : _GEN_3860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3862 = 9'h10d == _GEN_14118 ? phv_data_269 : _GEN_3861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3863 = 9'h10e == _GEN_14118 ? phv_data_270 : _GEN_3862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3864 = 9'h10f == _GEN_14118 ? phv_data_271 : _GEN_3863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3865 = 9'h110 == _GEN_14118 ? phv_data_272 : _GEN_3864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3866 = 9'h111 == _GEN_14118 ? phv_data_273 : _GEN_3865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3867 = 9'h112 == _GEN_14118 ? phv_data_274 : _GEN_3866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3868 = 9'h113 == _GEN_14118 ? phv_data_275 : _GEN_3867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3869 = 9'h114 == _GEN_14118 ? phv_data_276 : _GEN_3868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3870 = 9'h115 == _GEN_14118 ? phv_data_277 : _GEN_3869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3871 = 9'h116 == _GEN_14118 ? phv_data_278 : _GEN_3870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3872 = 9'h117 == _GEN_14118 ? phv_data_279 : _GEN_3871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3873 = 9'h118 == _GEN_14118 ? phv_data_280 : _GEN_3872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3874 = 9'h119 == _GEN_14118 ? phv_data_281 : _GEN_3873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3875 = 9'h11a == _GEN_14118 ? phv_data_282 : _GEN_3874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3876 = 9'h11b == _GEN_14118 ? phv_data_283 : _GEN_3875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3877 = 9'h11c == _GEN_14118 ? phv_data_284 : _GEN_3876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3878 = 9'h11d == _GEN_14118 ? phv_data_285 : _GEN_3877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3879 = 9'h11e == _GEN_14118 ? phv_data_286 : _GEN_3878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3880 = 9'h11f == _GEN_14118 ? phv_data_287 : _GEN_3879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3881 = 9'h120 == _GEN_14118 ? phv_data_288 : _GEN_3880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3882 = 9'h121 == _GEN_14118 ? phv_data_289 : _GEN_3881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3883 = 9'h122 == _GEN_14118 ? phv_data_290 : _GEN_3882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3884 = 9'h123 == _GEN_14118 ? phv_data_291 : _GEN_3883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3885 = 9'h124 == _GEN_14118 ? phv_data_292 : _GEN_3884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3886 = 9'h125 == _GEN_14118 ? phv_data_293 : _GEN_3885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3887 = 9'h126 == _GEN_14118 ? phv_data_294 : _GEN_3886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3888 = 9'h127 == _GEN_14118 ? phv_data_295 : _GEN_3887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3889 = 9'h128 == _GEN_14118 ? phv_data_296 : _GEN_3888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3890 = 9'h129 == _GEN_14118 ? phv_data_297 : _GEN_3889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3891 = 9'h12a == _GEN_14118 ? phv_data_298 : _GEN_3890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3892 = 9'h12b == _GEN_14118 ? phv_data_299 : _GEN_3891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3893 = 9'h12c == _GEN_14118 ? phv_data_300 : _GEN_3892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3894 = 9'h12d == _GEN_14118 ? phv_data_301 : _GEN_3893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3895 = 9'h12e == _GEN_14118 ? phv_data_302 : _GEN_3894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3896 = 9'h12f == _GEN_14118 ? phv_data_303 : _GEN_3895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3897 = 9'h130 == _GEN_14118 ? phv_data_304 : _GEN_3896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3898 = 9'h131 == _GEN_14118 ? phv_data_305 : _GEN_3897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3899 = 9'h132 == _GEN_14118 ? phv_data_306 : _GEN_3898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3900 = 9'h133 == _GEN_14118 ? phv_data_307 : _GEN_3899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3901 = 9'h134 == _GEN_14118 ? phv_data_308 : _GEN_3900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3902 = 9'h135 == _GEN_14118 ? phv_data_309 : _GEN_3901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3903 = 9'h136 == _GEN_14118 ? phv_data_310 : _GEN_3902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3904 = 9'h137 == _GEN_14118 ? phv_data_311 : _GEN_3903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3905 = 9'h138 == _GEN_14118 ? phv_data_312 : _GEN_3904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3906 = 9'h139 == _GEN_14118 ? phv_data_313 : _GEN_3905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3907 = 9'h13a == _GEN_14118 ? phv_data_314 : _GEN_3906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3908 = 9'h13b == _GEN_14118 ? phv_data_315 : _GEN_3907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3909 = 9'h13c == _GEN_14118 ? phv_data_316 : _GEN_3908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3910 = 9'h13d == _GEN_14118 ? phv_data_317 : _GEN_3909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3911 = 9'h13e == _GEN_14118 ? phv_data_318 : _GEN_3910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3912 = 9'h13f == _GEN_14118 ? phv_data_319 : _GEN_3911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3913 = 9'h140 == _GEN_14118 ? phv_data_320 : _GEN_3912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3914 = 9'h141 == _GEN_14118 ? phv_data_321 : _GEN_3913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3915 = 9'h142 == _GEN_14118 ? phv_data_322 : _GEN_3914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3916 = 9'h143 == _GEN_14118 ? phv_data_323 : _GEN_3915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3917 = 9'h144 == _GEN_14118 ? phv_data_324 : _GEN_3916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3918 = 9'h145 == _GEN_14118 ? phv_data_325 : _GEN_3917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3919 = 9'h146 == _GEN_14118 ? phv_data_326 : _GEN_3918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3920 = 9'h147 == _GEN_14118 ? phv_data_327 : _GEN_3919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3921 = 9'h148 == _GEN_14118 ? phv_data_328 : _GEN_3920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3922 = 9'h149 == _GEN_14118 ? phv_data_329 : _GEN_3921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3923 = 9'h14a == _GEN_14118 ? phv_data_330 : _GEN_3922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3924 = 9'h14b == _GEN_14118 ? phv_data_331 : _GEN_3923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3925 = 9'h14c == _GEN_14118 ? phv_data_332 : _GEN_3924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3926 = 9'h14d == _GEN_14118 ? phv_data_333 : _GEN_3925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3927 = 9'h14e == _GEN_14118 ? phv_data_334 : _GEN_3926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3928 = 9'h14f == _GEN_14118 ? phv_data_335 : _GEN_3927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3929 = 9'h150 == _GEN_14118 ? phv_data_336 : _GEN_3928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3930 = 9'h151 == _GEN_14118 ? phv_data_337 : _GEN_3929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3931 = 9'h152 == _GEN_14118 ? phv_data_338 : _GEN_3930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3932 = 9'h153 == _GEN_14118 ? phv_data_339 : _GEN_3931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3933 = 9'h154 == _GEN_14118 ? phv_data_340 : _GEN_3932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3934 = 9'h155 == _GEN_14118 ? phv_data_341 : _GEN_3933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3935 = 9'h156 == _GEN_14118 ? phv_data_342 : _GEN_3934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3936 = 9'h157 == _GEN_14118 ? phv_data_343 : _GEN_3935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3937 = 9'h158 == _GEN_14118 ? phv_data_344 : _GEN_3936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3938 = 9'h159 == _GEN_14118 ? phv_data_345 : _GEN_3937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3939 = 9'h15a == _GEN_14118 ? phv_data_346 : _GEN_3938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3940 = 9'h15b == _GEN_14118 ? phv_data_347 : _GEN_3939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3941 = 9'h15c == _GEN_14118 ? phv_data_348 : _GEN_3940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3942 = 9'h15d == _GEN_14118 ? phv_data_349 : _GEN_3941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3943 = 9'h15e == _GEN_14118 ? phv_data_350 : _GEN_3942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3944 = 9'h15f == _GEN_14118 ? phv_data_351 : _GEN_3943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3945 = 9'h160 == _GEN_14118 ? phv_data_352 : _GEN_3944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3946 = 9'h161 == _GEN_14118 ? phv_data_353 : _GEN_3945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3947 = 9'h162 == _GEN_14118 ? phv_data_354 : _GEN_3946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3948 = 9'h163 == _GEN_14118 ? phv_data_355 : _GEN_3947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3949 = 9'h164 == _GEN_14118 ? phv_data_356 : _GEN_3948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3950 = 9'h165 == _GEN_14118 ? phv_data_357 : _GEN_3949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3951 = 9'h166 == _GEN_14118 ? phv_data_358 : _GEN_3950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3952 = 9'h167 == _GEN_14118 ? phv_data_359 : _GEN_3951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3953 = 9'h168 == _GEN_14118 ? phv_data_360 : _GEN_3952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3954 = 9'h169 == _GEN_14118 ? phv_data_361 : _GEN_3953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3955 = 9'h16a == _GEN_14118 ? phv_data_362 : _GEN_3954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3956 = 9'h16b == _GEN_14118 ? phv_data_363 : _GEN_3955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3957 = 9'h16c == _GEN_14118 ? phv_data_364 : _GEN_3956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3958 = 9'h16d == _GEN_14118 ? phv_data_365 : _GEN_3957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3959 = 9'h16e == _GEN_14118 ? phv_data_366 : _GEN_3958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3960 = 9'h16f == _GEN_14118 ? phv_data_367 : _GEN_3959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3961 = 9'h170 == _GEN_14118 ? phv_data_368 : _GEN_3960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3962 = 9'h171 == _GEN_14118 ? phv_data_369 : _GEN_3961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3963 = 9'h172 == _GEN_14118 ? phv_data_370 : _GEN_3962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3964 = 9'h173 == _GEN_14118 ? phv_data_371 : _GEN_3963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3965 = 9'h174 == _GEN_14118 ? phv_data_372 : _GEN_3964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3966 = 9'h175 == _GEN_14118 ? phv_data_373 : _GEN_3965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3967 = 9'h176 == _GEN_14118 ? phv_data_374 : _GEN_3966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3968 = 9'h177 == _GEN_14118 ? phv_data_375 : _GEN_3967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3969 = 9'h178 == _GEN_14118 ? phv_data_376 : _GEN_3968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3970 = 9'h179 == _GEN_14118 ? phv_data_377 : _GEN_3969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3971 = 9'h17a == _GEN_14118 ? phv_data_378 : _GEN_3970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3972 = 9'h17b == _GEN_14118 ? phv_data_379 : _GEN_3971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3973 = 9'h17c == _GEN_14118 ? phv_data_380 : _GEN_3972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3974 = 9'h17d == _GEN_14118 ? phv_data_381 : _GEN_3973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3975 = 9'h17e == _GEN_14118 ? phv_data_382 : _GEN_3974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3976 = 9'h17f == _GEN_14118 ? phv_data_383 : _GEN_3975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3977 = 9'h180 == _GEN_14118 ? phv_data_384 : _GEN_3976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3978 = 9'h181 == _GEN_14118 ? phv_data_385 : _GEN_3977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3979 = 9'h182 == _GEN_14118 ? phv_data_386 : _GEN_3978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3980 = 9'h183 == _GEN_14118 ? phv_data_387 : _GEN_3979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3981 = 9'h184 == _GEN_14118 ? phv_data_388 : _GEN_3980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3982 = 9'h185 == _GEN_14118 ? phv_data_389 : _GEN_3981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3983 = 9'h186 == _GEN_14118 ? phv_data_390 : _GEN_3982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3984 = 9'h187 == _GEN_14118 ? phv_data_391 : _GEN_3983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3985 = 9'h188 == _GEN_14118 ? phv_data_392 : _GEN_3984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3986 = 9'h189 == _GEN_14118 ? phv_data_393 : _GEN_3985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3987 = 9'h18a == _GEN_14118 ? phv_data_394 : _GEN_3986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3988 = 9'h18b == _GEN_14118 ? phv_data_395 : _GEN_3987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3989 = 9'h18c == _GEN_14118 ? phv_data_396 : _GEN_3988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3990 = 9'h18d == _GEN_14118 ? phv_data_397 : _GEN_3989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3991 = 9'h18e == _GEN_14118 ? phv_data_398 : _GEN_3990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3992 = 9'h18f == _GEN_14118 ? phv_data_399 : _GEN_3991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3993 = 9'h190 == _GEN_14118 ? phv_data_400 : _GEN_3992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3994 = 9'h191 == _GEN_14118 ? phv_data_401 : _GEN_3993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3995 = 9'h192 == _GEN_14118 ? phv_data_402 : _GEN_3994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3996 = 9'h193 == _GEN_14118 ? phv_data_403 : _GEN_3995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3997 = 9'h194 == _GEN_14118 ? phv_data_404 : _GEN_3996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3998 = 9'h195 == _GEN_14118 ? phv_data_405 : _GEN_3997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3999 = 9'h196 == _GEN_14118 ? phv_data_406 : _GEN_3998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4000 = 9'h197 == _GEN_14118 ? phv_data_407 : _GEN_3999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4001 = 9'h198 == _GEN_14118 ? phv_data_408 : _GEN_4000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4002 = 9'h199 == _GEN_14118 ? phv_data_409 : _GEN_4001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4003 = 9'h19a == _GEN_14118 ? phv_data_410 : _GEN_4002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4004 = 9'h19b == _GEN_14118 ? phv_data_411 : _GEN_4003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4005 = 9'h19c == _GEN_14118 ? phv_data_412 : _GEN_4004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4006 = 9'h19d == _GEN_14118 ? phv_data_413 : _GEN_4005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4007 = 9'h19e == _GEN_14118 ? phv_data_414 : _GEN_4006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4008 = 9'h19f == _GEN_14118 ? phv_data_415 : _GEN_4007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4009 = 9'h1a0 == _GEN_14118 ? phv_data_416 : _GEN_4008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4010 = 9'h1a1 == _GEN_14118 ? phv_data_417 : _GEN_4009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4011 = 9'h1a2 == _GEN_14118 ? phv_data_418 : _GEN_4010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4012 = 9'h1a3 == _GEN_14118 ? phv_data_419 : _GEN_4011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4013 = 9'h1a4 == _GEN_14118 ? phv_data_420 : _GEN_4012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4014 = 9'h1a5 == _GEN_14118 ? phv_data_421 : _GEN_4013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4015 = 9'h1a6 == _GEN_14118 ? phv_data_422 : _GEN_4014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4016 = 9'h1a7 == _GEN_14118 ? phv_data_423 : _GEN_4015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4017 = 9'h1a8 == _GEN_14118 ? phv_data_424 : _GEN_4016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4018 = 9'h1a9 == _GEN_14118 ? phv_data_425 : _GEN_4017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4019 = 9'h1aa == _GEN_14118 ? phv_data_426 : _GEN_4018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4020 = 9'h1ab == _GEN_14118 ? phv_data_427 : _GEN_4019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4021 = 9'h1ac == _GEN_14118 ? phv_data_428 : _GEN_4020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4022 = 9'h1ad == _GEN_14118 ? phv_data_429 : _GEN_4021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4023 = 9'h1ae == _GEN_14118 ? phv_data_430 : _GEN_4022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4024 = 9'h1af == _GEN_14118 ? phv_data_431 : _GEN_4023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4025 = 9'h1b0 == _GEN_14118 ? phv_data_432 : _GEN_4024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4026 = 9'h1b1 == _GEN_14118 ? phv_data_433 : _GEN_4025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4027 = 9'h1b2 == _GEN_14118 ? phv_data_434 : _GEN_4026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4028 = 9'h1b3 == _GEN_14118 ? phv_data_435 : _GEN_4027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4029 = 9'h1b4 == _GEN_14118 ? phv_data_436 : _GEN_4028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4030 = 9'h1b5 == _GEN_14118 ? phv_data_437 : _GEN_4029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4031 = 9'h1b6 == _GEN_14118 ? phv_data_438 : _GEN_4030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4032 = 9'h1b7 == _GEN_14118 ? phv_data_439 : _GEN_4031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4033 = 9'h1b8 == _GEN_14118 ? phv_data_440 : _GEN_4032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4034 = 9'h1b9 == _GEN_14118 ? phv_data_441 : _GEN_4033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4035 = 9'h1ba == _GEN_14118 ? phv_data_442 : _GEN_4034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4036 = 9'h1bb == _GEN_14118 ? phv_data_443 : _GEN_4035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4037 = 9'h1bc == _GEN_14118 ? phv_data_444 : _GEN_4036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4038 = 9'h1bd == _GEN_14118 ? phv_data_445 : _GEN_4037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4039 = 9'h1be == _GEN_14118 ? phv_data_446 : _GEN_4038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4040 = 9'h1bf == _GEN_14118 ? phv_data_447 : _GEN_4039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4041 = 9'h1c0 == _GEN_14118 ? phv_data_448 : _GEN_4040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4042 = 9'h1c1 == _GEN_14118 ? phv_data_449 : _GEN_4041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4043 = 9'h1c2 == _GEN_14118 ? phv_data_450 : _GEN_4042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4044 = 9'h1c3 == _GEN_14118 ? phv_data_451 : _GEN_4043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4045 = 9'h1c4 == _GEN_14118 ? phv_data_452 : _GEN_4044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4046 = 9'h1c5 == _GEN_14118 ? phv_data_453 : _GEN_4045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4047 = 9'h1c6 == _GEN_14118 ? phv_data_454 : _GEN_4046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4048 = 9'h1c7 == _GEN_14118 ? phv_data_455 : _GEN_4047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4049 = 9'h1c8 == _GEN_14118 ? phv_data_456 : _GEN_4048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4050 = 9'h1c9 == _GEN_14118 ? phv_data_457 : _GEN_4049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4051 = 9'h1ca == _GEN_14118 ? phv_data_458 : _GEN_4050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4052 = 9'h1cb == _GEN_14118 ? phv_data_459 : _GEN_4051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4053 = 9'h1cc == _GEN_14118 ? phv_data_460 : _GEN_4052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4054 = 9'h1cd == _GEN_14118 ? phv_data_461 : _GEN_4053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4055 = 9'h1ce == _GEN_14118 ? phv_data_462 : _GEN_4054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4056 = 9'h1cf == _GEN_14118 ? phv_data_463 : _GEN_4055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4057 = 9'h1d0 == _GEN_14118 ? phv_data_464 : _GEN_4056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4058 = 9'h1d1 == _GEN_14118 ? phv_data_465 : _GEN_4057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4059 = 9'h1d2 == _GEN_14118 ? phv_data_466 : _GEN_4058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4060 = 9'h1d3 == _GEN_14118 ? phv_data_467 : _GEN_4059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4061 = 9'h1d4 == _GEN_14118 ? phv_data_468 : _GEN_4060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4062 = 9'h1d5 == _GEN_14118 ? phv_data_469 : _GEN_4061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4063 = 9'h1d6 == _GEN_14118 ? phv_data_470 : _GEN_4062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4064 = 9'h1d7 == _GEN_14118 ? phv_data_471 : _GEN_4063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4065 = 9'h1d8 == _GEN_14118 ? phv_data_472 : _GEN_4064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4066 = 9'h1d9 == _GEN_14118 ? phv_data_473 : _GEN_4065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4067 = 9'h1da == _GEN_14118 ? phv_data_474 : _GEN_4066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4068 = 9'h1db == _GEN_14118 ? phv_data_475 : _GEN_4067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4069 = 9'h1dc == _GEN_14118 ? phv_data_476 : _GEN_4068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4070 = 9'h1dd == _GEN_14118 ? phv_data_477 : _GEN_4069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4071 = 9'h1de == _GEN_14118 ? phv_data_478 : _GEN_4070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4072 = 9'h1df == _GEN_14118 ? phv_data_479 : _GEN_4071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4073 = 9'h1e0 == _GEN_14118 ? phv_data_480 : _GEN_4072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4074 = 9'h1e1 == _GEN_14118 ? phv_data_481 : _GEN_4073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4075 = 9'h1e2 == _GEN_14118 ? phv_data_482 : _GEN_4074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4076 = 9'h1e3 == _GEN_14118 ? phv_data_483 : _GEN_4075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4077 = 9'h1e4 == _GEN_14118 ? phv_data_484 : _GEN_4076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4078 = 9'h1e5 == _GEN_14118 ? phv_data_485 : _GEN_4077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4079 = 9'h1e6 == _GEN_14118 ? phv_data_486 : _GEN_4078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4080 = 9'h1e7 == _GEN_14118 ? phv_data_487 : _GEN_4079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4081 = 9'h1e8 == _GEN_14118 ? phv_data_488 : _GEN_4080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4082 = 9'h1e9 == _GEN_14118 ? phv_data_489 : _GEN_4081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4083 = 9'h1ea == _GEN_14118 ? phv_data_490 : _GEN_4082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4084 = 9'h1eb == _GEN_14118 ? phv_data_491 : _GEN_4083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4085 = 9'h1ec == _GEN_14118 ? phv_data_492 : _GEN_4084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4086 = 9'h1ed == _GEN_14118 ? phv_data_493 : _GEN_4085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4087 = 9'h1ee == _GEN_14118 ? phv_data_494 : _GEN_4086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4088 = 9'h1ef == _GEN_14118 ? phv_data_495 : _GEN_4087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4089 = 9'h1f0 == _GEN_14118 ? phv_data_496 : _GEN_4088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4090 = 9'h1f1 == _GEN_14118 ? phv_data_497 : _GEN_4089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4091 = 9'h1f2 == _GEN_14118 ? phv_data_498 : _GEN_4090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4092 = 9'h1f3 == _GEN_14118 ? phv_data_499 : _GEN_4091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4093 = 9'h1f4 == _GEN_14118 ? phv_data_500 : _GEN_4092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4094 = 9'h1f5 == _GEN_14118 ? phv_data_501 : _GEN_4093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4095 = 9'h1f6 == _GEN_14118 ? phv_data_502 : _GEN_4094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4096 = 9'h1f7 == _GEN_14118 ? phv_data_503 : _GEN_4095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4097 = 9'h1f8 == _GEN_14118 ? phv_data_504 : _GEN_4096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4098 = 9'h1f9 == _GEN_14118 ? phv_data_505 : _GEN_4097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4099 = 9'h1fa == _GEN_14118 ? phv_data_506 : _GEN_4098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4100 = 9'h1fb == _GEN_14118 ? phv_data_507 : _GEN_4099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4101 = 9'h1fc == _GEN_14118 ? phv_data_508 : _GEN_4100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4102 = 9'h1fd == _GEN_14118 ? phv_data_509 : _GEN_4101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4103 = 9'h1fe == _GEN_14118 ? phv_data_510 : _GEN_4102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4104 = 9'h1ff == _GEN_14118 ? phv_data_511 : _GEN_4103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_1_T_3 = {_GEN_3592,_GEN_4104,_GEN_2568,_GEN_3080}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_1 = local_offset_1 < end_offset ? _match_key_qbytes_1_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_2 = 8'h8 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_2_hi = local_offset_2[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_2_T = {match_key_qbytes_2_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_2_T_1 = {match_key_qbytes_2_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_2_T_2 = {match_key_qbytes_2_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_4107 = 8'h1 == _match_key_qbytes_2_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4108 = 8'h2 == _match_key_qbytes_2_T_2 ? phv_data_2 : _GEN_4107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4109 = 8'h3 == _match_key_qbytes_2_T_2 ? phv_data_3 : _GEN_4108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4110 = 8'h4 == _match_key_qbytes_2_T_2 ? phv_data_4 : _GEN_4109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4111 = 8'h5 == _match_key_qbytes_2_T_2 ? phv_data_5 : _GEN_4110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4112 = 8'h6 == _match_key_qbytes_2_T_2 ? phv_data_6 : _GEN_4111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4113 = 8'h7 == _match_key_qbytes_2_T_2 ? phv_data_7 : _GEN_4112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4114 = 8'h8 == _match_key_qbytes_2_T_2 ? phv_data_8 : _GEN_4113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4115 = 8'h9 == _match_key_qbytes_2_T_2 ? phv_data_9 : _GEN_4114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4116 = 8'ha == _match_key_qbytes_2_T_2 ? phv_data_10 : _GEN_4115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4117 = 8'hb == _match_key_qbytes_2_T_2 ? phv_data_11 : _GEN_4116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4118 = 8'hc == _match_key_qbytes_2_T_2 ? phv_data_12 : _GEN_4117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4119 = 8'hd == _match_key_qbytes_2_T_2 ? phv_data_13 : _GEN_4118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4120 = 8'he == _match_key_qbytes_2_T_2 ? phv_data_14 : _GEN_4119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4121 = 8'hf == _match_key_qbytes_2_T_2 ? phv_data_15 : _GEN_4120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4122 = 8'h10 == _match_key_qbytes_2_T_2 ? phv_data_16 : _GEN_4121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4123 = 8'h11 == _match_key_qbytes_2_T_2 ? phv_data_17 : _GEN_4122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4124 = 8'h12 == _match_key_qbytes_2_T_2 ? phv_data_18 : _GEN_4123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4125 = 8'h13 == _match_key_qbytes_2_T_2 ? phv_data_19 : _GEN_4124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4126 = 8'h14 == _match_key_qbytes_2_T_2 ? phv_data_20 : _GEN_4125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4127 = 8'h15 == _match_key_qbytes_2_T_2 ? phv_data_21 : _GEN_4126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4128 = 8'h16 == _match_key_qbytes_2_T_2 ? phv_data_22 : _GEN_4127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4129 = 8'h17 == _match_key_qbytes_2_T_2 ? phv_data_23 : _GEN_4128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4130 = 8'h18 == _match_key_qbytes_2_T_2 ? phv_data_24 : _GEN_4129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4131 = 8'h19 == _match_key_qbytes_2_T_2 ? phv_data_25 : _GEN_4130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4132 = 8'h1a == _match_key_qbytes_2_T_2 ? phv_data_26 : _GEN_4131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4133 = 8'h1b == _match_key_qbytes_2_T_2 ? phv_data_27 : _GEN_4132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4134 = 8'h1c == _match_key_qbytes_2_T_2 ? phv_data_28 : _GEN_4133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4135 = 8'h1d == _match_key_qbytes_2_T_2 ? phv_data_29 : _GEN_4134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4136 = 8'h1e == _match_key_qbytes_2_T_2 ? phv_data_30 : _GEN_4135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4137 = 8'h1f == _match_key_qbytes_2_T_2 ? phv_data_31 : _GEN_4136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4138 = 8'h20 == _match_key_qbytes_2_T_2 ? phv_data_32 : _GEN_4137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4139 = 8'h21 == _match_key_qbytes_2_T_2 ? phv_data_33 : _GEN_4138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4140 = 8'h22 == _match_key_qbytes_2_T_2 ? phv_data_34 : _GEN_4139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4141 = 8'h23 == _match_key_qbytes_2_T_2 ? phv_data_35 : _GEN_4140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4142 = 8'h24 == _match_key_qbytes_2_T_2 ? phv_data_36 : _GEN_4141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4143 = 8'h25 == _match_key_qbytes_2_T_2 ? phv_data_37 : _GEN_4142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4144 = 8'h26 == _match_key_qbytes_2_T_2 ? phv_data_38 : _GEN_4143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4145 = 8'h27 == _match_key_qbytes_2_T_2 ? phv_data_39 : _GEN_4144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4146 = 8'h28 == _match_key_qbytes_2_T_2 ? phv_data_40 : _GEN_4145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4147 = 8'h29 == _match_key_qbytes_2_T_2 ? phv_data_41 : _GEN_4146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4148 = 8'h2a == _match_key_qbytes_2_T_2 ? phv_data_42 : _GEN_4147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4149 = 8'h2b == _match_key_qbytes_2_T_2 ? phv_data_43 : _GEN_4148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4150 = 8'h2c == _match_key_qbytes_2_T_2 ? phv_data_44 : _GEN_4149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4151 = 8'h2d == _match_key_qbytes_2_T_2 ? phv_data_45 : _GEN_4150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4152 = 8'h2e == _match_key_qbytes_2_T_2 ? phv_data_46 : _GEN_4151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4153 = 8'h2f == _match_key_qbytes_2_T_2 ? phv_data_47 : _GEN_4152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4154 = 8'h30 == _match_key_qbytes_2_T_2 ? phv_data_48 : _GEN_4153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4155 = 8'h31 == _match_key_qbytes_2_T_2 ? phv_data_49 : _GEN_4154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4156 = 8'h32 == _match_key_qbytes_2_T_2 ? phv_data_50 : _GEN_4155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4157 = 8'h33 == _match_key_qbytes_2_T_2 ? phv_data_51 : _GEN_4156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4158 = 8'h34 == _match_key_qbytes_2_T_2 ? phv_data_52 : _GEN_4157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4159 = 8'h35 == _match_key_qbytes_2_T_2 ? phv_data_53 : _GEN_4158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4160 = 8'h36 == _match_key_qbytes_2_T_2 ? phv_data_54 : _GEN_4159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4161 = 8'h37 == _match_key_qbytes_2_T_2 ? phv_data_55 : _GEN_4160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4162 = 8'h38 == _match_key_qbytes_2_T_2 ? phv_data_56 : _GEN_4161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4163 = 8'h39 == _match_key_qbytes_2_T_2 ? phv_data_57 : _GEN_4162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4164 = 8'h3a == _match_key_qbytes_2_T_2 ? phv_data_58 : _GEN_4163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4165 = 8'h3b == _match_key_qbytes_2_T_2 ? phv_data_59 : _GEN_4164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4166 = 8'h3c == _match_key_qbytes_2_T_2 ? phv_data_60 : _GEN_4165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4167 = 8'h3d == _match_key_qbytes_2_T_2 ? phv_data_61 : _GEN_4166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4168 = 8'h3e == _match_key_qbytes_2_T_2 ? phv_data_62 : _GEN_4167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4169 = 8'h3f == _match_key_qbytes_2_T_2 ? phv_data_63 : _GEN_4168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4170 = 8'h40 == _match_key_qbytes_2_T_2 ? phv_data_64 : _GEN_4169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4171 = 8'h41 == _match_key_qbytes_2_T_2 ? phv_data_65 : _GEN_4170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4172 = 8'h42 == _match_key_qbytes_2_T_2 ? phv_data_66 : _GEN_4171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4173 = 8'h43 == _match_key_qbytes_2_T_2 ? phv_data_67 : _GEN_4172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4174 = 8'h44 == _match_key_qbytes_2_T_2 ? phv_data_68 : _GEN_4173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4175 = 8'h45 == _match_key_qbytes_2_T_2 ? phv_data_69 : _GEN_4174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4176 = 8'h46 == _match_key_qbytes_2_T_2 ? phv_data_70 : _GEN_4175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4177 = 8'h47 == _match_key_qbytes_2_T_2 ? phv_data_71 : _GEN_4176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4178 = 8'h48 == _match_key_qbytes_2_T_2 ? phv_data_72 : _GEN_4177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4179 = 8'h49 == _match_key_qbytes_2_T_2 ? phv_data_73 : _GEN_4178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4180 = 8'h4a == _match_key_qbytes_2_T_2 ? phv_data_74 : _GEN_4179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4181 = 8'h4b == _match_key_qbytes_2_T_2 ? phv_data_75 : _GEN_4180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4182 = 8'h4c == _match_key_qbytes_2_T_2 ? phv_data_76 : _GEN_4181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4183 = 8'h4d == _match_key_qbytes_2_T_2 ? phv_data_77 : _GEN_4182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4184 = 8'h4e == _match_key_qbytes_2_T_2 ? phv_data_78 : _GEN_4183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4185 = 8'h4f == _match_key_qbytes_2_T_2 ? phv_data_79 : _GEN_4184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4186 = 8'h50 == _match_key_qbytes_2_T_2 ? phv_data_80 : _GEN_4185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4187 = 8'h51 == _match_key_qbytes_2_T_2 ? phv_data_81 : _GEN_4186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4188 = 8'h52 == _match_key_qbytes_2_T_2 ? phv_data_82 : _GEN_4187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4189 = 8'h53 == _match_key_qbytes_2_T_2 ? phv_data_83 : _GEN_4188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4190 = 8'h54 == _match_key_qbytes_2_T_2 ? phv_data_84 : _GEN_4189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4191 = 8'h55 == _match_key_qbytes_2_T_2 ? phv_data_85 : _GEN_4190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4192 = 8'h56 == _match_key_qbytes_2_T_2 ? phv_data_86 : _GEN_4191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4193 = 8'h57 == _match_key_qbytes_2_T_2 ? phv_data_87 : _GEN_4192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4194 = 8'h58 == _match_key_qbytes_2_T_2 ? phv_data_88 : _GEN_4193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4195 = 8'h59 == _match_key_qbytes_2_T_2 ? phv_data_89 : _GEN_4194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4196 = 8'h5a == _match_key_qbytes_2_T_2 ? phv_data_90 : _GEN_4195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4197 = 8'h5b == _match_key_qbytes_2_T_2 ? phv_data_91 : _GEN_4196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4198 = 8'h5c == _match_key_qbytes_2_T_2 ? phv_data_92 : _GEN_4197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4199 = 8'h5d == _match_key_qbytes_2_T_2 ? phv_data_93 : _GEN_4198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4200 = 8'h5e == _match_key_qbytes_2_T_2 ? phv_data_94 : _GEN_4199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4201 = 8'h5f == _match_key_qbytes_2_T_2 ? phv_data_95 : _GEN_4200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4202 = 8'h60 == _match_key_qbytes_2_T_2 ? phv_data_96 : _GEN_4201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4203 = 8'h61 == _match_key_qbytes_2_T_2 ? phv_data_97 : _GEN_4202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4204 = 8'h62 == _match_key_qbytes_2_T_2 ? phv_data_98 : _GEN_4203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4205 = 8'h63 == _match_key_qbytes_2_T_2 ? phv_data_99 : _GEN_4204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4206 = 8'h64 == _match_key_qbytes_2_T_2 ? phv_data_100 : _GEN_4205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4207 = 8'h65 == _match_key_qbytes_2_T_2 ? phv_data_101 : _GEN_4206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4208 = 8'h66 == _match_key_qbytes_2_T_2 ? phv_data_102 : _GEN_4207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4209 = 8'h67 == _match_key_qbytes_2_T_2 ? phv_data_103 : _GEN_4208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4210 = 8'h68 == _match_key_qbytes_2_T_2 ? phv_data_104 : _GEN_4209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4211 = 8'h69 == _match_key_qbytes_2_T_2 ? phv_data_105 : _GEN_4210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4212 = 8'h6a == _match_key_qbytes_2_T_2 ? phv_data_106 : _GEN_4211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4213 = 8'h6b == _match_key_qbytes_2_T_2 ? phv_data_107 : _GEN_4212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4214 = 8'h6c == _match_key_qbytes_2_T_2 ? phv_data_108 : _GEN_4213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4215 = 8'h6d == _match_key_qbytes_2_T_2 ? phv_data_109 : _GEN_4214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4216 = 8'h6e == _match_key_qbytes_2_T_2 ? phv_data_110 : _GEN_4215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4217 = 8'h6f == _match_key_qbytes_2_T_2 ? phv_data_111 : _GEN_4216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4218 = 8'h70 == _match_key_qbytes_2_T_2 ? phv_data_112 : _GEN_4217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4219 = 8'h71 == _match_key_qbytes_2_T_2 ? phv_data_113 : _GEN_4218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4220 = 8'h72 == _match_key_qbytes_2_T_2 ? phv_data_114 : _GEN_4219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4221 = 8'h73 == _match_key_qbytes_2_T_2 ? phv_data_115 : _GEN_4220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4222 = 8'h74 == _match_key_qbytes_2_T_2 ? phv_data_116 : _GEN_4221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4223 = 8'h75 == _match_key_qbytes_2_T_2 ? phv_data_117 : _GEN_4222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4224 = 8'h76 == _match_key_qbytes_2_T_2 ? phv_data_118 : _GEN_4223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4225 = 8'h77 == _match_key_qbytes_2_T_2 ? phv_data_119 : _GEN_4224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4226 = 8'h78 == _match_key_qbytes_2_T_2 ? phv_data_120 : _GEN_4225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4227 = 8'h79 == _match_key_qbytes_2_T_2 ? phv_data_121 : _GEN_4226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4228 = 8'h7a == _match_key_qbytes_2_T_2 ? phv_data_122 : _GEN_4227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4229 = 8'h7b == _match_key_qbytes_2_T_2 ? phv_data_123 : _GEN_4228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4230 = 8'h7c == _match_key_qbytes_2_T_2 ? phv_data_124 : _GEN_4229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4231 = 8'h7d == _match_key_qbytes_2_T_2 ? phv_data_125 : _GEN_4230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4232 = 8'h7e == _match_key_qbytes_2_T_2 ? phv_data_126 : _GEN_4231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4233 = 8'h7f == _match_key_qbytes_2_T_2 ? phv_data_127 : _GEN_4232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4234 = 8'h80 == _match_key_qbytes_2_T_2 ? phv_data_128 : _GEN_4233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4235 = 8'h81 == _match_key_qbytes_2_T_2 ? phv_data_129 : _GEN_4234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4236 = 8'h82 == _match_key_qbytes_2_T_2 ? phv_data_130 : _GEN_4235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4237 = 8'h83 == _match_key_qbytes_2_T_2 ? phv_data_131 : _GEN_4236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4238 = 8'h84 == _match_key_qbytes_2_T_2 ? phv_data_132 : _GEN_4237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4239 = 8'h85 == _match_key_qbytes_2_T_2 ? phv_data_133 : _GEN_4238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4240 = 8'h86 == _match_key_qbytes_2_T_2 ? phv_data_134 : _GEN_4239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4241 = 8'h87 == _match_key_qbytes_2_T_2 ? phv_data_135 : _GEN_4240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4242 = 8'h88 == _match_key_qbytes_2_T_2 ? phv_data_136 : _GEN_4241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4243 = 8'h89 == _match_key_qbytes_2_T_2 ? phv_data_137 : _GEN_4242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4244 = 8'h8a == _match_key_qbytes_2_T_2 ? phv_data_138 : _GEN_4243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4245 = 8'h8b == _match_key_qbytes_2_T_2 ? phv_data_139 : _GEN_4244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4246 = 8'h8c == _match_key_qbytes_2_T_2 ? phv_data_140 : _GEN_4245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4247 = 8'h8d == _match_key_qbytes_2_T_2 ? phv_data_141 : _GEN_4246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4248 = 8'h8e == _match_key_qbytes_2_T_2 ? phv_data_142 : _GEN_4247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4249 = 8'h8f == _match_key_qbytes_2_T_2 ? phv_data_143 : _GEN_4248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4250 = 8'h90 == _match_key_qbytes_2_T_2 ? phv_data_144 : _GEN_4249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4251 = 8'h91 == _match_key_qbytes_2_T_2 ? phv_data_145 : _GEN_4250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4252 = 8'h92 == _match_key_qbytes_2_T_2 ? phv_data_146 : _GEN_4251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4253 = 8'h93 == _match_key_qbytes_2_T_2 ? phv_data_147 : _GEN_4252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4254 = 8'h94 == _match_key_qbytes_2_T_2 ? phv_data_148 : _GEN_4253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4255 = 8'h95 == _match_key_qbytes_2_T_2 ? phv_data_149 : _GEN_4254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4256 = 8'h96 == _match_key_qbytes_2_T_2 ? phv_data_150 : _GEN_4255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4257 = 8'h97 == _match_key_qbytes_2_T_2 ? phv_data_151 : _GEN_4256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4258 = 8'h98 == _match_key_qbytes_2_T_2 ? phv_data_152 : _GEN_4257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4259 = 8'h99 == _match_key_qbytes_2_T_2 ? phv_data_153 : _GEN_4258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4260 = 8'h9a == _match_key_qbytes_2_T_2 ? phv_data_154 : _GEN_4259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4261 = 8'h9b == _match_key_qbytes_2_T_2 ? phv_data_155 : _GEN_4260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4262 = 8'h9c == _match_key_qbytes_2_T_2 ? phv_data_156 : _GEN_4261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4263 = 8'h9d == _match_key_qbytes_2_T_2 ? phv_data_157 : _GEN_4262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4264 = 8'h9e == _match_key_qbytes_2_T_2 ? phv_data_158 : _GEN_4263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4265 = 8'h9f == _match_key_qbytes_2_T_2 ? phv_data_159 : _GEN_4264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4266 = 8'ha0 == _match_key_qbytes_2_T_2 ? phv_data_160 : _GEN_4265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4267 = 8'ha1 == _match_key_qbytes_2_T_2 ? phv_data_161 : _GEN_4266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4268 = 8'ha2 == _match_key_qbytes_2_T_2 ? phv_data_162 : _GEN_4267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4269 = 8'ha3 == _match_key_qbytes_2_T_2 ? phv_data_163 : _GEN_4268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4270 = 8'ha4 == _match_key_qbytes_2_T_2 ? phv_data_164 : _GEN_4269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4271 = 8'ha5 == _match_key_qbytes_2_T_2 ? phv_data_165 : _GEN_4270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4272 = 8'ha6 == _match_key_qbytes_2_T_2 ? phv_data_166 : _GEN_4271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4273 = 8'ha7 == _match_key_qbytes_2_T_2 ? phv_data_167 : _GEN_4272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4274 = 8'ha8 == _match_key_qbytes_2_T_2 ? phv_data_168 : _GEN_4273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4275 = 8'ha9 == _match_key_qbytes_2_T_2 ? phv_data_169 : _GEN_4274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4276 = 8'haa == _match_key_qbytes_2_T_2 ? phv_data_170 : _GEN_4275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4277 = 8'hab == _match_key_qbytes_2_T_2 ? phv_data_171 : _GEN_4276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4278 = 8'hac == _match_key_qbytes_2_T_2 ? phv_data_172 : _GEN_4277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4279 = 8'had == _match_key_qbytes_2_T_2 ? phv_data_173 : _GEN_4278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4280 = 8'hae == _match_key_qbytes_2_T_2 ? phv_data_174 : _GEN_4279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4281 = 8'haf == _match_key_qbytes_2_T_2 ? phv_data_175 : _GEN_4280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4282 = 8'hb0 == _match_key_qbytes_2_T_2 ? phv_data_176 : _GEN_4281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4283 = 8'hb1 == _match_key_qbytes_2_T_2 ? phv_data_177 : _GEN_4282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4284 = 8'hb2 == _match_key_qbytes_2_T_2 ? phv_data_178 : _GEN_4283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4285 = 8'hb3 == _match_key_qbytes_2_T_2 ? phv_data_179 : _GEN_4284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4286 = 8'hb4 == _match_key_qbytes_2_T_2 ? phv_data_180 : _GEN_4285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4287 = 8'hb5 == _match_key_qbytes_2_T_2 ? phv_data_181 : _GEN_4286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4288 = 8'hb6 == _match_key_qbytes_2_T_2 ? phv_data_182 : _GEN_4287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4289 = 8'hb7 == _match_key_qbytes_2_T_2 ? phv_data_183 : _GEN_4288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4290 = 8'hb8 == _match_key_qbytes_2_T_2 ? phv_data_184 : _GEN_4289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4291 = 8'hb9 == _match_key_qbytes_2_T_2 ? phv_data_185 : _GEN_4290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4292 = 8'hba == _match_key_qbytes_2_T_2 ? phv_data_186 : _GEN_4291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4293 = 8'hbb == _match_key_qbytes_2_T_2 ? phv_data_187 : _GEN_4292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4294 = 8'hbc == _match_key_qbytes_2_T_2 ? phv_data_188 : _GEN_4293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4295 = 8'hbd == _match_key_qbytes_2_T_2 ? phv_data_189 : _GEN_4294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4296 = 8'hbe == _match_key_qbytes_2_T_2 ? phv_data_190 : _GEN_4295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4297 = 8'hbf == _match_key_qbytes_2_T_2 ? phv_data_191 : _GEN_4296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4298 = 8'hc0 == _match_key_qbytes_2_T_2 ? phv_data_192 : _GEN_4297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4299 = 8'hc1 == _match_key_qbytes_2_T_2 ? phv_data_193 : _GEN_4298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4300 = 8'hc2 == _match_key_qbytes_2_T_2 ? phv_data_194 : _GEN_4299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4301 = 8'hc3 == _match_key_qbytes_2_T_2 ? phv_data_195 : _GEN_4300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4302 = 8'hc4 == _match_key_qbytes_2_T_2 ? phv_data_196 : _GEN_4301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4303 = 8'hc5 == _match_key_qbytes_2_T_2 ? phv_data_197 : _GEN_4302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4304 = 8'hc6 == _match_key_qbytes_2_T_2 ? phv_data_198 : _GEN_4303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4305 = 8'hc7 == _match_key_qbytes_2_T_2 ? phv_data_199 : _GEN_4304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4306 = 8'hc8 == _match_key_qbytes_2_T_2 ? phv_data_200 : _GEN_4305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4307 = 8'hc9 == _match_key_qbytes_2_T_2 ? phv_data_201 : _GEN_4306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4308 = 8'hca == _match_key_qbytes_2_T_2 ? phv_data_202 : _GEN_4307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4309 = 8'hcb == _match_key_qbytes_2_T_2 ? phv_data_203 : _GEN_4308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4310 = 8'hcc == _match_key_qbytes_2_T_2 ? phv_data_204 : _GEN_4309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4311 = 8'hcd == _match_key_qbytes_2_T_2 ? phv_data_205 : _GEN_4310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4312 = 8'hce == _match_key_qbytes_2_T_2 ? phv_data_206 : _GEN_4311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4313 = 8'hcf == _match_key_qbytes_2_T_2 ? phv_data_207 : _GEN_4312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4314 = 8'hd0 == _match_key_qbytes_2_T_2 ? phv_data_208 : _GEN_4313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4315 = 8'hd1 == _match_key_qbytes_2_T_2 ? phv_data_209 : _GEN_4314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4316 = 8'hd2 == _match_key_qbytes_2_T_2 ? phv_data_210 : _GEN_4315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4317 = 8'hd3 == _match_key_qbytes_2_T_2 ? phv_data_211 : _GEN_4316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4318 = 8'hd4 == _match_key_qbytes_2_T_2 ? phv_data_212 : _GEN_4317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4319 = 8'hd5 == _match_key_qbytes_2_T_2 ? phv_data_213 : _GEN_4318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4320 = 8'hd6 == _match_key_qbytes_2_T_2 ? phv_data_214 : _GEN_4319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4321 = 8'hd7 == _match_key_qbytes_2_T_2 ? phv_data_215 : _GEN_4320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4322 = 8'hd8 == _match_key_qbytes_2_T_2 ? phv_data_216 : _GEN_4321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4323 = 8'hd9 == _match_key_qbytes_2_T_2 ? phv_data_217 : _GEN_4322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4324 = 8'hda == _match_key_qbytes_2_T_2 ? phv_data_218 : _GEN_4323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4325 = 8'hdb == _match_key_qbytes_2_T_2 ? phv_data_219 : _GEN_4324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4326 = 8'hdc == _match_key_qbytes_2_T_2 ? phv_data_220 : _GEN_4325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4327 = 8'hdd == _match_key_qbytes_2_T_2 ? phv_data_221 : _GEN_4326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4328 = 8'hde == _match_key_qbytes_2_T_2 ? phv_data_222 : _GEN_4327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4329 = 8'hdf == _match_key_qbytes_2_T_2 ? phv_data_223 : _GEN_4328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4330 = 8'he0 == _match_key_qbytes_2_T_2 ? phv_data_224 : _GEN_4329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4331 = 8'he1 == _match_key_qbytes_2_T_2 ? phv_data_225 : _GEN_4330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4332 = 8'he2 == _match_key_qbytes_2_T_2 ? phv_data_226 : _GEN_4331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4333 = 8'he3 == _match_key_qbytes_2_T_2 ? phv_data_227 : _GEN_4332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4334 = 8'he4 == _match_key_qbytes_2_T_2 ? phv_data_228 : _GEN_4333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4335 = 8'he5 == _match_key_qbytes_2_T_2 ? phv_data_229 : _GEN_4334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4336 = 8'he6 == _match_key_qbytes_2_T_2 ? phv_data_230 : _GEN_4335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4337 = 8'he7 == _match_key_qbytes_2_T_2 ? phv_data_231 : _GEN_4336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4338 = 8'he8 == _match_key_qbytes_2_T_2 ? phv_data_232 : _GEN_4337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4339 = 8'he9 == _match_key_qbytes_2_T_2 ? phv_data_233 : _GEN_4338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4340 = 8'hea == _match_key_qbytes_2_T_2 ? phv_data_234 : _GEN_4339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4341 = 8'heb == _match_key_qbytes_2_T_2 ? phv_data_235 : _GEN_4340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4342 = 8'hec == _match_key_qbytes_2_T_2 ? phv_data_236 : _GEN_4341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4343 = 8'hed == _match_key_qbytes_2_T_2 ? phv_data_237 : _GEN_4342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4344 = 8'hee == _match_key_qbytes_2_T_2 ? phv_data_238 : _GEN_4343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4345 = 8'hef == _match_key_qbytes_2_T_2 ? phv_data_239 : _GEN_4344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4346 = 8'hf0 == _match_key_qbytes_2_T_2 ? phv_data_240 : _GEN_4345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4347 = 8'hf1 == _match_key_qbytes_2_T_2 ? phv_data_241 : _GEN_4346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4348 = 8'hf2 == _match_key_qbytes_2_T_2 ? phv_data_242 : _GEN_4347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4349 = 8'hf3 == _match_key_qbytes_2_T_2 ? phv_data_243 : _GEN_4348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4350 = 8'hf4 == _match_key_qbytes_2_T_2 ? phv_data_244 : _GEN_4349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4351 = 8'hf5 == _match_key_qbytes_2_T_2 ? phv_data_245 : _GEN_4350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4352 = 8'hf6 == _match_key_qbytes_2_T_2 ? phv_data_246 : _GEN_4351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4353 = 8'hf7 == _match_key_qbytes_2_T_2 ? phv_data_247 : _GEN_4352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4354 = 8'hf8 == _match_key_qbytes_2_T_2 ? phv_data_248 : _GEN_4353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4355 = 8'hf9 == _match_key_qbytes_2_T_2 ? phv_data_249 : _GEN_4354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4356 = 8'hfa == _match_key_qbytes_2_T_2 ? phv_data_250 : _GEN_4355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4357 = 8'hfb == _match_key_qbytes_2_T_2 ? phv_data_251 : _GEN_4356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4358 = 8'hfc == _match_key_qbytes_2_T_2 ? phv_data_252 : _GEN_4357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4359 = 8'hfd == _match_key_qbytes_2_T_2 ? phv_data_253 : _GEN_4358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4360 = 8'hfe == _match_key_qbytes_2_T_2 ? phv_data_254 : _GEN_4359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4361 = 8'hff == _match_key_qbytes_2_T_2 ? phv_data_255 : _GEN_4360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_14374 = {{1'd0}, _match_key_qbytes_2_T_2}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4362 = 9'h100 == _GEN_14374 ? phv_data_256 : _GEN_4361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4363 = 9'h101 == _GEN_14374 ? phv_data_257 : _GEN_4362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4364 = 9'h102 == _GEN_14374 ? phv_data_258 : _GEN_4363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4365 = 9'h103 == _GEN_14374 ? phv_data_259 : _GEN_4364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4366 = 9'h104 == _GEN_14374 ? phv_data_260 : _GEN_4365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4367 = 9'h105 == _GEN_14374 ? phv_data_261 : _GEN_4366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4368 = 9'h106 == _GEN_14374 ? phv_data_262 : _GEN_4367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4369 = 9'h107 == _GEN_14374 ? phv_data_263 : _GEN_4368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4370 = 9'h108 == _GEN_14374 ? phv_data_264 : _GEN_4369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4371 = 9'h109 == _GEN_14374 ? phv_data_265 : _GEN_4370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4372 = 9'h10a == _GEN_14374 ? phv_data_266 : _GEN_4371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4373 = 9'h10b == _GEN_14374 ? phv_data_267 : _GEN_4372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4374 = 9'h10c == _GEN_14374 ? phv_data_268 : _GEN_4373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4375 = 9'h10d == _GEN_14374 ? phv_data_269 : _GEN_4374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4376 = 9'h10e == _GEN_14374 ? phv_data_270 : _GEN_4375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4377 = 9'h10f == _GEN_14374 ? phv_data_271 : _GEN_4376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4378 = 9'h110 == _GEN_14374 ? phv_data_272 : _GEN_4377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4379 = 9'h111 == _GEN_14374 ? phv_data_273 : _GEN_4378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4380 = 9'h112 == _GEN_14374 ? phv_data_274 : _GEN_4379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4381 = 9'h113 == _GEN_14374 ? phv_data_275 : _GEN_4380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4382 = 9'h114 == _GEN_14374 ? phv_data_276 : _GEN_4381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4383 = 9'h115 == _GEN_14374 ? phv_data_277 : _GEN_4382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4384 = 9'h116 == _GEN_14374 ? phv_data_278 : _GEN_4383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4385 = 9'h117 == _GEN_14374 ? phv_data_279 : _GEN_4384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4386 = 9'h118 == _GEN_14374 ? phv_data_280 : _GEN_4385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4387 = 9'h119 == _GEN_14374 ? phv_data_281 : _GEN_4386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4388 = 9'h11a == _GEN_14374 ? phv_data_282 : _GEN_4387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4389 = 9'h11b == _GEN_14374 ? phv_data_283 : _GEN_4388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4390 = 9'h11c == _GEN_14374 ? phv_data_284 : _GEN_4389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4391 = 9'h11d == _GEN_14374 ? phv_data_285 : _GEN_4390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4392 = 9'h11e == _GEN_14374 ? phv_data_286 : _GEN_4391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4393 = 9'h11f == _GEN_14374 ? phv_data_287 : _GEN_4392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4394 = 9'h120 == _GEN_14374 ? phv_data_288 : _GEN_4393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4395 = 9'h121 == _GEN_14374 ? phv_data_289 : _GEN_4394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4396 = 9'h122 == _GEN_14374 ? phv_data_290 : _GEN_4395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4397 = 9'h123 == _GEN_14374 ? phv_data_291 : _GEN_4396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4398 = 9'h124 == _GEN_14374 ? phv_data_292 : _GEN_4397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4399 = 9'h125 == _GEN_14374 ? phv_data_293 : _GEN_4398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4400 = 9'h126 == _GEN_14374 ? phv_data_294 : _GEN_4399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4401 = 9'h127 == _GEN_14374 ? phv_data_295 : _GEN_4400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4402 = 9'h128 == _GEN_14374 ? phv_data_296 : _GEN_4401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4403 = 9'h129 == _GEN_14374 ? phv_data_297 : _GEN_4402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4404 = 9'h12a == _GEN_14374 ? phv_data_298 : _GEN_4403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4405 = 9'h12b == _GEN_14374 ? phv_data_299 : _GEN_4404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4406 = 9'h12c == _GEN_14374 ? phv_data_300 : _GEN_4405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4407 = 9'h12d == _GEN_14374 ? phv_data_301 : _GEN_4406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4408 = 9'h12e == _GEN_14374 ? phv_data_302 : _GEN_4407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4409 = 9'h12f == _GEN_14374 ? phv_data_303 : _GEN_4408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4410 = 9'h130 == _GEN_14374 ? phv_data_304 : _GEN_4409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4411 = 9'h131 == _GEN_14374 ? phv_data_305 : _GEN_4410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4412 = 9'h132 == _GEN_14374 ? phv_data_306 : _GEN_4411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4413 = 9'h133 == _GEN_14374 ? phv_data_307 : _GEN_4412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4414 = 9'h134 == _GEN_14374 ? phv_data_308 : _GEN_4413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4415 = 9'h135 == _GEN_14374 ? phv_data_309 : _GEN_4414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4416 = 9'h136 == _GEN_14374 ? phv_data_310 : _GEN_4415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4417 = 9'h137 == _GEN_14374 ? phv_data_311 : _GEN_4416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4418 = 9'h138 == _GEN_14374 ? phv_data_312 : _GEN_4417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4419 = 9'h139 == _GEN_14374 ? phv_data_313 : _GEN_4418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4420 = 9'h13a == _GEN_14374 ? phv_data_314 : _GEN_4419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4421 = 9'h13b == _GEN_14374 ? phv_data_315 : _GEN_4420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4422 = 9'h13c == _GEN_14374 ? phv_data_316 : _GEN_4421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4423 = 9'h13d == _GEN_14374 ? phv_data_317 : _GEN_4422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4424 = 9'h13e == _GEN_14374 ? phv_data_318 : _GEN_4423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4425 = 9'h13f == _GEN_14374 ? phv_data_319 : _GEN_4424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4426 = 9'h140 == _GEN_14374 ? phv_data_320 : _GEN_4425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4427 = 9'h141 == _GEN_14374 ? phv_data_321 : _GEN_4426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4428 = 9'h142 == _GEN_14374 ? phv_data_322 : _GEN_4427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4429 = 9'h143 == _GEN_14374 ? phv_data_323 : _GEN_4428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4430 = 9'h144 == _GEN_14374 ? phv_data_324 : _GEN_4429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4431 = 9'h145 == _GEN_14374 ? phv_data_325 : _GEN_4430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4432 = 9'h146 == _GEN_14374 ? phv_data_326 : _GEN_4431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4433 = 9'h147 == _GEN_14374 ? phv_data_327 : _GEN_4432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4434 = 9'h148 == _GEN_14374 ? phv_data_328 : _GEN_4433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4435 = 9'h149 == _GEN_14374 ? phv_data_329 : _GEN_4434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4436 = 9'h14a == _GEN_14374 ? phv_data_330 : _GEN_4435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4437 = 9'h14b == _GEN_14374 ? phv_data_331 : _GEN_4436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4438 = 9'h14c == _GEN_14374 ? phv_data_332 : _GEN_4437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4439 = 9'h14d == _GEN_14374 ? phv_data_333 : _GEN_4438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4440 = 9'h14e == _GEN_14374 ? phv_data_334 : _GEN_4439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4441 = 9'h14f == _GEN_14374 ? phv_data_335 : _GEN_4440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4442 = 9'h150 == _GEN_14374 ? phv_data_336 : _GEN_4441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4443 = 9'h151 == _GEN_14374 ? phv_data_337 : _GEN_4442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4444 = 9'h152 == _GEN_14374 ? phv_data_338 : _GEN_4443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4445 = 9'h153 == _GEN_14374 ? phv_data_339 : _GEN_4444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4446 = 9'h154 == _GEN_14374 ? phv_data_340 : _GEN_4445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4447 = 9'h155 == _GEN_14374 ? phv_data_341 : _GEN_4446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4448 = 9'h156 == _GEN_14374 ? phv_data_342 : _GEN_4447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4449 = 9'h157 == _GEN_14374 ? phv_data_343 : _GEN_4448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4450 = 9'h158 == _GEN_14374 ? phv_data_344 : _GEN_4449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4451 = 9'h159 == _GEN_14374 ? phv_data_345 : _GEN_4450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4452 = 9'h15a == _GEN_14374 ? phv_data_346 : _GEN_4451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4453 = 9'h15b == _GEN_14374 ? phv_data_347 : _GEN_4452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4454 = 9'h15c == _GEN_14374 ? phv_data_348 : _GEN_4453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4455 = 9'h15d == _GEN_14374 ? phv_data_349 : _GEN_4454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4456 = 9'h15e == _GEN_14374 ? phv_data_350 : _GEN_4455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4457 = 9'h15f == _GEN_14374 ? phv_data_351 : _GEN_4456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4458 = 9'h160 == _GEN_14374 ? phv_data_352 : _GEN_4457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4459 = 9'h161 == _GEN_14374 ? phv_data_353 : _GEN_4458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4460 = 9'h162 == _GEN_14374 ? phv_data_354 : _GEN_4459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4461 = 9'h163 == _GEN_14374 ? phv_data_355 : _GEN_4460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4462 = 9'h164 == _GEN_14374 ? phv_data_356 : _GEN_4461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4463 = 9'h165 == _GEN_14374 ? phv_data_357 : _GEN_4462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4464 = 9'h166 == _GEN_14374 ? phv_data_358 : _GEN_4463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4465 = 9'h167 == _GEN_14374 ? phv_data_359 : _GEN_4464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4466 = 9'h168 == _GEN_14374 ? phv_data_360 : _GEN_4465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4467 = 9'h169 == _GEN_14374 ? phv_data_361 : _GEN_4466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4468 = 9'h16a == _GEN_14374 ? phv_data_362 : _GEN_4467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4469 = 9'h16b == _GEN_14374 ? phv_data_363 : _GEN_4468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4470 = 9'h16c == _GEN_14374 ? phv_data_364 : _GEN_4469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4471 = 9'h16d == _GEN_14374 ? phv_data_365 : _GEN_4470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4472 = 9'h16e == _GEN_14374 ? phv_data_366 : _GEN_4471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4473 = 9'h16f == _GEN_14374 ? phv_data_367 : _GEN_4472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4474 = 9'h170 == _GEN_14374 ? phv_data_368 : _GEN_4473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4475 = 9'h171 == _GEN_14374 ? phv_data_369 : _GEN_4474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4476 = 9'h172 == _GEN_14374 ? phv_data_370 : _GEN_4475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4477 = 9'h173 == _GEN_14374 ? phv_data_371 : _GEN_4476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4478 = 9'h174 == _GEN_14374 ? phv_data_372 : _GEN_4477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4479 = 9'h175 == _GEN_14374 ? phv_data_373 : _GEN_4478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4480 = 9'h176 == _GEN_14374 ? phv_data_374 : _GEN_4479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4481 = 9'h177 == _GEN_14374 ? phv_data_375 : _GEN_4480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4482 = 9'h178 == _GEN_14374 ? phv_data_376 : _GEN_4481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4483 = 9'h179 == _GEN_14374 ? phv_data_377 : _GEN_4482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4484 = 9'h17a == _GEN_14374 ? phv_data_378 : _GEN_4483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4485 = 9'h17b == _GEN_14374 ? phv_data_379 : _GEN_4484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4486 = 9'h17c == _GEN_14374 ? phv_data_380 : _GEN_4485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4487 = 9'h17d == _GEN_14374 ? phv_data_381 : _GEN_4486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4488 = 9'h17e == _GEN_14374 ? phv_data_382 : _GEN_4487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4489 = 9'h17f == _GEN_14374 ? phv_data_383 : _GEN_4488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4490 = 9'h180 == _GEN_14374 ? phv_data_384 : _GEN_4489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4491 = 9'h181 == _GEN_14374 ? phv_data_385 : _GEN_4490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4492 = 9'h182 == _GEN_14374 ? phv_data_386 : _GEN_4491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4493 = 9'h183 == _GEN_14374 ? phv_data_387 : _GEN_4492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4494 = 9'h184 == _GEN_14374 ? phv_data_388 : _GEN_4493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4495 = 9'h185 == _GEN_14374 ? phv_data_389 : _GEN_4494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4496 = 9'h186 == _GEN_14374 ? phv_data_390 : _GEN_4495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4497 = 9'h187 == _GEN_14374 ? phv_data_391 : _GEN_4496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4498 = 9'h188 == _GEN_14374 ? phv_data_392 : _GEN_4497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4499 = 9'h189 == _GEN_14374 ? phv_data_393 : _GEN_4498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4500 = 9'h18a == _GEN_14374 ? phv_data_394 : _GEN_4499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4501 = 9'h18b == _GEN_14374 ? phv_data_395 : _GEN_4500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4502 = 9'h18c == _GEN_14374 ? phv_data_396 : _GEN_4501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4503 = 9'h18d == _GEN_14374 ? phv_data_397 : _GEN_4502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4504 = 9'h18e == _GEN_14374 ? phv_data_398 : _GEN_4503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4505 = 9'h18f == _GEN_14374 ? phv_data_399 : _GEN_4504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4506 = 9'h190 == _GEN_14374 ? phv_data_400 : _GEN_4505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4507 = 9'h191 == _GEN_14374 ? phv_data_401 : _GEN_4506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4508 = 9'h192 == _GEN_14374 ? phv_data_402 : _GEN_4507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4509 = 9'h193 == _GEN_14374 ? phv_data_403 : _GEN_4508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4510 = 9'h194 == _GEN_14374 ? phv_data_404 : _GEN_4509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4511 = 9'h195 == _GEN_14374 ? phv_data_405 : _GEN_4510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4512 = 9'h196 == _GEN_14374 ? phv_data_406 : _GEN_4511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4513 = 9'h197 == _GEN_14374 ? phv_data_407 : _GEN_4512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4514 = 9'h198 == _GEN_14374 ? phv_data_408 : _GEN_4513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4515 = 9'h199 == _GEN_14374 ? phv_data_409 : _GEN_4514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4516 = 9'h19a == _GEN_14374 ? phv_data_410 : _GEN_4515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4517 = 9'h19b == _GEN_14374 ? phv_data_411 : _GEN_4516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4518 = 9'h19c == _GEN_14374 ? phv_data_412 : _GEN_4517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4519 = 9'h19d == _GEN_14374 ? phv_data_413 : _GEN_4518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4520 = 9'h19e == _GEN_14374 ? phv_data_414 : _GEN_4519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4521 = 9'h19f == _GEN_14374 ? phv_data_415 : _GEN_4520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4522 = 9'h1a0 == _GEN_14374 ? phv_data_416 : _GEN_4521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4523 = 9'h1a1 == _GEN_14374 ? phv_data_417 : _GEN_4522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4524 = 9'h1a2 == _GEN_14374 ? phv_data_418 : _GEN_4523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4525 = 9'h1a3 == _GEN_14374 ? phv_data_419 : _GEN_4524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4526 = 9'h1a4 == _GEN_14374 ? phv_data_420 : _GEN_4525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4527 = 9'h1a5 == _GEN_14374 ? phv_data_421 : _GEN_4526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4528 = 9'h1a6 == _GEN_14374 ? phv_data_422 : _GEN_4527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4529 = 9'h1a7 == _GEN_14374 ? phv_data_423 : _GEN_4528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4530 = 9'h1a8 == _GEN_14374 ? phv_data_424 : _GEN_4529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4531 = 9'h1a9 == _GEN_14374 ? phv_data_425 : _GEN_4530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4532 = 9'h1aa == _GEN_14374 ? phv_data_426 : _GEN_4531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4533 = 9'h1ab == _GEN_14374 ? phv_data_427 : _GEN_4532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4534 = 9'h1ac == _GEN_14374 ? phv_data_428 : _GEN_4533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4535 = 9'h1ad == _GEN_14374 ? phv_data_429 : _GEN_4534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4536 = 9'h1ae == _GEN_14374 ? phv_data_430 : _GEN_4535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4537 = 9'h1af == _GEN_14374 ? phv_data_431 : _GEN_4536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4538 = 9'h1b0 == _GEN_14374 ? phv_data_432 : _GEN_4537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4539 = 9'h1b1 == _GEN_14374 ? phv_data_433 : _GEN_4538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4540 = 9'h1b2 == _GEN_14374 ? phv_data_434 : _GEN_4539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4541 = 9'h1b3 == _GEN_14374 ? phv_data_435 : _GEN_4540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4542 = 9'h1b4 == _GEN_14374 ? phv_data_436 : _GEN_4541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4543 = 9'h1b5 == _GEN_14374 ? phv_data_437 : _GEN_4542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4544 = 9'h1b6 == _GEN_14374 ? phv_data_438 : _GEN_4543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4545 = 9'h1b7 == _GEN_14374 ? phv_data_439 : _GEN_4544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4546 = 9'h1b8 == _GEN_14374 ? phv_data_440 : _GEN_4545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4547 = 9'h1b9 == _GEN_14374 ? phv_data_441 : _GEN_4546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4548 = 9'h1ba == _GEN_14374 ? phv_data_442 : _GEN_4547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4549 = 9'h1bb == _GEN_14374 ? phv_data_443 : _GEN_4548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4550 = 9'h1bc == _GEN_14374 ? phv_data_444 : _GEN_4549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4551 = 9'h1bd == _GEN_14374 ? phv_data_445 : _GEN_4550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4552 = 9'h1be == _GEN_14374 ? phv_data_446 : _GEN_4551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4553 = 9'h1bf == _GEN_14374 ? phv_data_447 : _GEN_4552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4554 = 9'h1c0 == _GEN_14374 ? phv_data_448 : _GEN_4553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4555 = 9'h1c1 == _GEN_14374 ? phv_data_449 : _GEN_4554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4556 = 9'h1c2 == _GEN_14374 ? phv_data_450 : _GEN_4555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4557 = 9'h1c3 == _GEN_14374 ? phv_data_451 : _GEN_4556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4558 = 9'h1c4 == _GEN_14374 ? phv_data_452 : _GEN_4557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4559 = 9'h1c5 == _GEN_14374 ? phv_data_453 : _GEN_4558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4560 = 9'h1c6 == _GEN_14374 ? phv_data_454 : _GEN_4559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4561 = 9'h1c7 == _GEN_14374 ? phv_data_455 : _GEN_4560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4562 = 9'h1c8 == _GEN_14374 ? phv_data_456 : _GEN_4561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4563 = 9'h1c9 == _GEN_14374 ? phv_data_457 : _GEN_4562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4564 = 9'h1ca == _GEN_14374 ? phv_data_458 : _GEN_4563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4565 = 9'h1cb == _GEN_14374 ? phv_data_459 : _GEN_4564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4566 = 9'h1cc == _GEN_14374 ? phv_data_460 : _GEN_4565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4567 = 9'h1cd == _GEN_14374 ? phv_data_461 : _GEN_4566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4568 = 9'h1ce == _GEN_14374 ? phv_data_462 : _GEN_4567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4569 = 9'h1cf == _GEN_14374 ? phv_data_463 : _GEN_4568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4570 = 9'h1d0 == _GEN_14374 ? phv_data_464 : _GEN_4569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4571 = 9'h1d1 == _GEN_14374 ? phv_data_465 : _GEN_4570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4572 = 9'h1d2 == _GEN_14374 ? phv_data_466 : _GEN_4571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4573 = 9'h1d3 == _GEN_14374 ? phv_data_467 : _GEN_4572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4574 = 9'h1d4 == _GEN_14374 ? phv_data_468 : _GEN_4573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4575 = 9'h1d5 == _GEN_14374 ? phv_data_469 : _GEN_4574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4576 = 9'h1d6 == _GEN_14374 ? phv_data_470 : _GEN_4575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4577 = 9'h1d7 == _GEN_14374 ? phv_data_471 : _GEN_4576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4578 = 9'h1d8 == _GEN_14374 ? phv_data_472 : _GEN_4577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4579 = 9'h1d9 == _GEN_14374 ? phv_data_473 : _GEN_4578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4580 = 9'h1da == _GEN_14374 ? phv_data_474 : _GEN_4579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4581 = 9'h1db == _GEN_14374 ? phv_data_475 : _GEN_4580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4582 = 9'h1dc == _GEN_14374 ? phv_data_476 : _GEN_4581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4583 = 9'h1dd == _GEN_14374 ? phv_data_477 : _GEN_4582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4584 = 9'h1de == _GEN_14374 ? phv_data_478 : _GEN_4583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4585 = 9'h1df == _GEN_14374 ? phv_data_479 : _GEN_4584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4586 = 9'h1e0 == _GEN_14374 ? phv_data_480 : _GEN_4585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4587 = 9'h1e1 == _GEN_14374 ? phv_data_481 : _GEN_4586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4588 = 9'h1e2 == _GEN_14374 ? phv_data_482 : _GEN_4587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4589 = 9'h1e3 == _GEN_14374 ? phv_data_483 : _GEN_4588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4590 = 9'h1e4 == _GEN_14374 ? phv_data_484 : _GEN_4589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4591 = 9'h1e5 == _GEN_14374 ? phv_data_485 : _GEN_4590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4592 = 9'h1e6 == _GEN_14374 ? phv_data_486 : _GEN_4591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4593 = 9'h1e7 == _GEN_14374 ? phv_data_487 : _GEN_4592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4594 = 9'h1e8 == _GEN_14374 ? phv_data_488 : _GEN_4593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4595 = 9'h1e9 == _GEN_14374 ? phv_data_489 : _GEN_4594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4596 = 9'h1ea == _GEN_14374 ? phv_data_490 : _GEN_4595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4597 = 9'h1eb == _GEN_14374 ? phv_data_491 : _GEN_4596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4598 = 9'h1ec == _GEN_14374 ? phv_data_492 : _GEN_4597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4599 = 9'h1ed == _GEN_14374 ? phv_data_493 : _GEN_4598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4600 = 9'h1ee == _GEN_14374 ? phv_data_494 : _GEN_4599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4601 = 9'h1ef == _GEN_14374 ? phv_data_495 : _GEN_4600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4602 = 9'h1f0 == _GEN_14374 ? phv_data_496 : _GEN_4601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4603 = 9'h1f1 == _GEN_14374 ? phv_data_497 : _GEN_4602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4604 = 9'h1f2 == _GEN_14374 ? phv_data_498 : _GEN_4603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4605 = 9'h1f3 == _GEN_14374 ? phv_data_499 : _GEN_4604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4606 = 9'h1f4 == _GEN_14374 ? phv_data_500 : _GEN_4605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4607 = 9'h1f5 == _GEN_14374 ? phv_data_501 : _GEN_4606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4608 = 9'h1f6 == _GEN_14374 ? phv_data_502 : _GEN_4607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4609 = 9'h1f7 == _GEN_14374 ? phv_data_503 : _GEN_4608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4610 = 9'h1f8 == _GEN_14374 ? phv_data_504 : _GEN_4609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4611 = 9'h1f9 == _GEN_14374 ? phv_data_505 : _GEN_4610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4612 = 9'h1fa == _GEN_14374 ? phv_data_506 : _GEN_4611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4613 = 9'h1fb == _GEN_14374 ? phv_data_507 : _GEN_4612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4614 = 9'h1fc == _GEN_14374 ? phv_data_508 : _GEN_4613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4615 = 9'h1fd == _GEN_14374 ? phv_data_509 : _GEN_4614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4616 = 9'h1fe == _GEN_14374 ? phv_data_510 : _GEN_4615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4617 = 9'h1ff == _GEN_14374 ? phv_data_511 : _GEN_4616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4619 = 8'h1 == local_offset_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4620 = 8'h2 == local_offset_2 ? phv_data_2 : _GEN_4619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4621 = 8'h3 == local_offset_2 ? phv_data_3 : _GEN_4620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4622 = 8'h4 == local_offset_2 ? phv_data_4 : _GEN_4621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4623 = 8'h5 == local_offset_2 ? phv_data_5 : _GEN_4622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4624 = 8'h6 == local_offset_2 ? phv_data_6 : _GEN_4623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4625 = 8'h7 == local_offset_2 ? phv_data_7 : _GEN_4624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4626 = 8'h8 == local_offset_2 ? phv_data_8 : _GEN_4625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4627 = 8'h9 == local_offset_2 ? phv_data_9 : _GEN_4626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4628 = 8'ha == local_offset_2 ? phv_data_10 : _GEN_4627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4629 = 8'hb == local_offset_2 ? phv_data_11 : _GEN_4628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4630 = 8'hc == local_offset_2 ? phv_data_12 : _GEN_4629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4631 = 8'hd == local_offset_2 ? phv_data_13 : _GEN_4630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4632 = 8'he == local_offset_2 ? phv_data_14 : _GEN_4631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4633 = 8'hf == local_offset_2 ? phv_data_15 : _GEN_4632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4634 = 8'h10 == local_offset_2 ? phv_data_16 : _GEN_4633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4635 = 8'h11 == local_offset_2 ? phv_data_17 : _GEN_4634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4636 = 8'h12 == local_offset_2 ? phv_data_18 : _GEN_4635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4637 = 8'h13 == local_offset_2 ? phv_data_19 : _GEN_4636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4638 = 8'h14 == local_offset_2 ? phv_data_20 : _GEN_4637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4639 = 8'h15 == local_offset_2 ? phv_data_21 : _GEN_4638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4640 = 8'h16 == local_offset_2 ? phv_data_22 : _GEN_4639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4641 = 8'h17 == local_offset_2 ? phv_data_23 : _GEN_4640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4642 = 8'h18 == local_offset_2 ? phv_data_24 : _GEN_4641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4643 = 8'h19 == local_offset_2 ? phv_data_25 : _GEN_4642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4644 = 8'h1a == local_offset_2 ? phv_data_26 : _GEN_4643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4645 = 8'h1b == local_offset_2 ? phv_data_27 : _GEN_4644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4646 = 8'h1c == local_offset_2 ? phv_data_28 : _GEN_4645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4647 = 8'h1d == local_offset_2 ? phv_data_29 : _GEN_4646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4648 = 8'h1e == local_offset_2 ? phv_data_30 : _GEN_4647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4649 = 8'h1f == local_offset_2 ? phv_data_31 : _GEN_4648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4650 = 8'h20 == local_offset_2 ? phv_data_32 : _GEN_4649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4651 = 8'h21 == local_offset_2 ? phv_data_33 : _GEN_4650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4652 = 8'h22 == local_offset_2 ? phv_data_34 : _GEN_4651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4653 = 8'h23 == local_offset_2 ? phv_data_35 : _GEN_4652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4654 = 8'h24 == local_offset_2 ? phv_data_36 : _GEN_4653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4655 = 8'h25 == local_offset_2 ? phv_data_37 : _GEN_4654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4656 = 8'h26 == local_offset_2 ? phv_data_38 : _GEN_4655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4657 = 8'h27 == local_offset_2 ? phv_data_39 : _GEN_4656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4658 = 8'h28 == local_offset_2 ? phv_data_40 : _GEN_4657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4659 = 8'h29 == local_offset_2 ? phv_data_41 : _GEN_4658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4660 = 8'h2a == local_offset_2 ? phv_data_42 : _GEN_4659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4661 = 8'h2b == local_offset_2 ? phv_data_43 : _GEN_4660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4662 = 8'h2c == local_offset_2 ? phv_data_44 : _GEN_4661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4663 = 8'h2d == local_offset_2 ? phv_data_45 : _GEN_4662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4664 = 8'h2e == local_offset_2 ? phv_data_46 : _GEN_4663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4665 = 8'h2f == local_offset_2 ? phv_data_47 : _GEN_4664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4666 = 8'h30 == local_offset_2 ? phv_data_48 : _GEN_4665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4667 = 8'h31 == local_offset_2 ? phv_data_49 : _GEN_4666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4668 = 8'h32 == local_offset_2 ? phv_data_50 : _GEN_4667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4669 = 8'h33 == local_offset_2 ? phv_data_51 : _GEN_4668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4670 = 8'h34 == local_offset_2 ? phv_data_52 : _GEN_4669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4671 = 8'h35 == local_offset_2 ? phv_data_53 : _GEN_4670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4672 = 8'h36 == local_offset_2 ? phv_data_54 : _GEN_4671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4673 = 8'h37 == local_offset_2 ? phv_data_55 : _GEN_4672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4674 = 8'h38 == local_offset_2 ? phv_data_56 : _GEN_4673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4675 = 8'h39 == local_offset_2 ? phv_data_57 : _GEN_4674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4676 = 8'h3a == local_offset_2 ? phv_data_58 : _GEN_4675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4677 = 8'h3b == local_offset_2 ? phv_data_59 : _GEN_4676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4678 = 8'h3c == local_offset_2 ? phv_data_60 : _GEN_4677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4679 = 8'h3d == local_offset_2 ? phv_data_61 : _GEN_4678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4680 = 8'h3e == local_offset_2 ? phv_data_62 : _GEN_4679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4681 = 8'h3f == local_offset_2 ? phv_data_63 : _GEN_4680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4682 = 8'h40 == local_offset_2 ? phv_data_64 : _GEN_4681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4683 = 8'h41 == local_offset_2 ? phv_data_65 : _GEN_4682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4684 = 8'h42 == local_offset_2 ? phv_data_66 : _GEN_4683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4685 = 8'h43 == local_offset_2 ? phv_data_67 : _GEN_4684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4686 = 8'h44 == local_offset_2 ? phv_data_68 : _GEN_4685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4687 = 8'h45 == local_offset_2 ? phv_data_69 : _GEN_4686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4688 = 8'h46 == local_offset_2 ? phv_data_70 : _GEN_4687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4689 = 8'h47 == local_offset_2 ? phv_data_71 : _GEN_4688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4690 = 8'h48 == local_offset_2 ? phv_data_72 : _GEN_4689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4691 = 8'h49 == local_offset_2 ? phv_data_73 : _GEN_4690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4692 = 8'h4a == local_offset_2 ? phv_data_74 : _GEN_4691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4693 = 8'h4b == local_offset_2 ? phv_data_75 : _GEN_4692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4694 = 8'h4c == local_offset_2 ? phv_data_76 : _GEN_4693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4695 = 8'h4d == local_offset_2 ? phv_data_77 : _GEN_4694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4696 = 8'h4e == local_offset_2 ? phv_data_78 : _GEN_4695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4697 = 8'h4f == local_offset_2 ? phv_data_79 : _GEN_4696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4698 = 8'h50 == local_offset_2 ? phv_data_80 : _GEN_4697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4699 = 8'h51 == local_offset_2 ? phv_data_81 : _GEN_4698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4700 = 8'h52 == local_offset_2 ? phv_data_82 : _GEN_4699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4701 = 8'h53 == local_offset_2 ? phv_data_83 : _GEN_4700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4702 = 8'h54 == local_offset_2 ? phv_data_84 : _GEN_4701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4703 = 8'h55 == local_offset_2 ? phv_data_85 : _GEN_4702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4704 = 8'h56 == local_offset_2 ? phv_data_86 : _GEN_4703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4705 = 8'h57 == local_offset_2 ? phv_data_87 : _GEN_4704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4706 = 8'h58 == local_offset_2 ? phv_data_88 : _GEN_4705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4707 = 8'h59 == local_offset_2 ? phv_data_89 : _GEN_4706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4708 = 8'h5a == local_offset_2 ? phv_data_90 : _GEN_4707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4709 = 8'h5b == local_offset_2 ? phv_data_91 : _GEN_4708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4710 = 8'h5c == local_offset_2 ? phv_data_92 : _GEN_4709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4711 = 8'h5d == local_offset_2 ? phv_data_93 : _GEN_4710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4712 = 8'h5e == local_offset_2 ? phv_data_94 : _GEN_4711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4713 = 8'h5f == local_offset_2 ? phv_data_95 : _GEN_4712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4714 = 8'h60 == local_offset_2 ? phv_data_96 : _GEN_4713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4715 = 8'h61 == local_offset_2 ? phv_data_97 : _GEN_4714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4716 = 8'h62 == local_offset_2 ? phv_data_98 : _GEN_4715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4717 = 8'h63 == local_offset_2 ? phv_data_99 : _GEN_4716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4718 = 8'h64 == local_offset_2 ? phv_data_100 : _GEN_4717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4719 = 8'h65 == local_offset_2 ? phv_data_101 : _GEN_4718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4720 = 8'h66 == local_offset_2 ? phv_data_102 : _GEN_4719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4721 = 8'h67 == local_offset_2 ? phv_data_103 : _GEN_4720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4722 = 8'h68 == local_offset_2 ? phv_data_104 : _GEN_4721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4723 = 8'h69 == local_offset_2 ? phv_data_105 : _GEN_4722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4724 = 8'h6a == local_offset_2 ? phv_data_106 : _GEN_4723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4725 = 8'h6b == local_offset_2 ? phv_data_107 : _GEN_4724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4726 = 8'h6c == local_offset_2 ? phv_data_108 : _GEN_4725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4727 = 8'h6d == local_offset_2 ? phv_data_109 : _GEN_4726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4728 = 8'h6e == local_offset_2 ? phv_data_110 : _GEN_4727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4729 = 8'h6f == local_offset_2 ? phv_data_111 : _GEN_4728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4730 = 8'h70 == local_offset_2 ? phv_data_112 : _GEN_4729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4731 = 8'h71 == local_offset_2 ? phv_data_113 : _GEN_4730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4732 = 8'h72 == local_offset_2 ? phv_data_114 : _GEN_4731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4733 = 8'h73 == local_offset_2 ? phv_data_115 : _GEN_4732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4734 = 8'h74 == local_offset_2 ? phv_data_116 : _GEN_4733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4735 = 8'h75 == local_offset_2 ? phv_data_117 : _GEN_4734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4736 = 8'h76 == local_offset_2 ? phv_data_118 : _GEN_4735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4737 = 8'h77 == local_offset_2 ? phv_data_119 : _GEN_4736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4738 = 8'h78 == local_offset_2 ? phv_data_120 : _GEN_4737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4739 = 8'h79 == local_offset_2 ? phv_data_121 : _GEN_4738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4740 = 8'h7a == local_offset_2 ? phv_data_122 : _GEN_4739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4741 = 8'h7b == local_offset_2 ? phv_data_123 : _GEN_4740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4742 = 8'h7c == local_offset_2 ? phv_data_124 : _GEN_4741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4743 = 8'h7d == local_offset_2 ? phv_data_125 : _GEN_4742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4744 = 8'h7e == local_offset_2 ? phv_data_126 : _GEN_4743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4745 = 8'h7f == local_offset_2 ? phv_data_127 : _GEN_4744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4746 = 8'h80 == local_offset_2 ? phv_data_128 : _GEN_4745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4747 = 8'h81 == local_offset_2 ? phv_data_129 : _GEN_4746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4748 = 8'h82 == local_offset_2 ? phv_data_130 : _GEN_4747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4749 = 8'h83 == local_offset_2 ? phv_data_131 : _GEN_4748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4750 = 8'h84 == local_offset_2 ? phv_data_132 : _GEN_4749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4751 = 8'h85 == local_offset_2 ? phv_data_133 : _GEN_4750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4752 = 8'h86 == local_offset_2 ? phv_data_134 : _GEN_4751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4753 = 8'h87 == local_offset_2 ? phv_data_135 : _GEN_4752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4754 = 8'h88 == local_offset_2 ? phv_data_136 : _GEN_4753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4755 = 8'h89 == local_offset_2 ? phv_data_137 : _GEN_4754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4756 = 8'h8a == local_offset_2 ? phv_data_138 : _GEN_4755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4757 = 8'h8b == local_offset_2 ? phv_data_139 : _GEN_4756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4758 = 8'h8c == local_offset_2 ? phv_data_140 : _GEN_4757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4759 = 8'h8d == local_offset_2 ? phv_data_141 : _GEN_4758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4760 = 8'h8e == local_offset_2 ? phv_data_142 : _GEN_4759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4761 = 8'h8f == local_offset_2 ? phv_data_143 : _GEN_4760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4762 = 8'h90 == local_offset_2 ? phv_data_144 : _GEN_4761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4763 = 8'h91 == local_offset_2 ? phv_data_145 : _GEN_4762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4764 = 8'h92 == local_offset_2 ? phv_data_146 : _GEN_4763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4765 = 8'h93 == local_offset_2 ? phv_data_147 : _GEN_4764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4766 = 8'h94 == local_offset_2 ? phv_data_148 : _GEN_4765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4767 = 8'h95 == local_offset_2 ? phv_data_149 : _GEN_4766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4768 = 8'h96 == local_offset_2 ? phv_data_150 : _GEN_4767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4769 = 8'h97 == local_offset_2 ? phv_data_151 : _GEN_4768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4770 = 8'h98 == local_offset_2 ? phv_data_152 : _GEN_4769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4771 = 8'h99 == local_offset_2 ? phv_data_153 : _GEN_4770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4772 = 8'h9a == local_offset_2 ? phv_data_154 : _GEN_4771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4773 = 8'h9b == local_offset_2 ? phv_data_155 : _GEN_4772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4774 = 8'h9c == local_offset_2 ? phv_data_156 : _GEN_4773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4775 = 8'h9d == local_offset_2 ? phv_data_157 : _GEN_4774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4776 = 8'h9e == local_offset_2 ? phv_data_158 : _GEN_4775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4777 = 8'h9f == local_offset_2 ? phv_data_159 : _GEN_4776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4778 = 8'ha0 == local_offset_2 ? phv_data_160 : _GEN_4777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4779 = 8'ha1 == local_offset_2 ? phv_data_161 : _GEN_4778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4780 = 8'ha2 == local_offset_2 ? phv_data_162 : _GEN_4779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4781 = 8'ha3 == local_offset_2 ? phv_data_163 : _GEN_4780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4782 = 8'ha4 == local_offset_2 ? phv_data_164 : _GEN_4781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4783 = 8'ha5 == local_offset_2 ? phv_data_165 : _GEN_4782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4784 = 8'ha6 == local_offset_2 ? phv_data_166 : _GEN_4783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4785 = 8'ha7 == local_offset_2 ? phv_data_167 : _GEN_4784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4786 = 8'ha8 == local_offset_2 ? phv_data_168 : _GEN_4785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4787 = 8'ha9 == local_offset_2 ? phv_data_169 : _GEN_4786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4788 = 8'haa == local_offset_2 ? phv_data_170 : _GEN_4787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4789 = 8'hab == local_offset_2 ? phv_data_171 : _GEN_4788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4790 = 8'hac == local_offset_2 ? phv_data_172 : _GEN_4789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4791 = 8'had == local_offset_2 ? phv_data_173 : _GEN_4790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4792 = 8'hae == local_offset_2 ? phv_data_174 : _GEN_4791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4793 = 8'haf == local_offset_2 ? phv_data_175 : _GEN_4792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4794 = 8'hb0 == local_offset_2 ? phv_data_176 : _GEN_4793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4795 = 8'hb1 == local_offset_2 ? phv_data_177 : _GEN_4794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4796 = 8'hb2 == local_offset_2 ? phv_data_178 : _GEN_4795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4797 = 8'hb3 == local_offset_2 ? phv_data_179 : _GEN_4796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4798 = 8'hb4 == local_offset_2 ? phv_data_180 : _GEN_4797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4799 = 8'hb5 == local_offset_2 ? phv_data_181 : _GEN_4798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4800 = 8'hb6 == local_offset_2 ? phv_data_182 : _GEN_4799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4801 = 8'hb7 == local_offset_2 ? phv_data_183 : _GEN_4800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4802 = 8'hb8 == local_offset_2 ? phv_data_184 : _GEN_4801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4803 = 8'hb9 == local_offset_2 ? phv_data_185 : _GEN_4802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4804 = 8'hba == local_offset_2 ? phv_data_186 : _GEN_4803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4805 = 8'hbb == local_offset_2 ? phv_data_187 : _GEN_4804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4806 = 8'hbc == local_offset_2 ? phv_data_188 : _GEN_4805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4807 = 8'hbd == local_offset_2 ? phv_data_189 : _GEN_4806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4808 = 8'hbe == local_offset_2 ? phv_data_190 : _GEN_4807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4809 = 8'hbf == local_offset_2 ? phv_data_191 : _GEN_4808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4810 = 8'hc0 == local_offset_2 ? phv_data_192 : _GEN_4809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4811 = 8'hc1 == local_offset_2 ? phv_data_193 : _GEN_4810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4812 = 8'hc2 == local_offset_2 ? phv_data_194 : _GEN_4811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4813 = 8'hc3 == local_offset_2 ? phv_data_195 : _GEN_4812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4814 = 8'hc4 == local_offset_2 ? phv_data_196 : _GEN_4813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4815 = 8'hc5 == local_offset_2 ? phv_data_197 : _GEN_4814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4816 = 8'hc6 == local_offset_2 ? phv_data_198 : _GEN_4815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4817 = 8'hc7 == local_offset_2 ? phv_data_199 : _GEN_4816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4818 = 8'hc8 == local_offset_2 ? phv_data_200 : _GEN_4817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4819 = 8'hc9 == local_offset_2 ? phv_data_201 : _GEN_4818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4820 = 8'hca == local_offset_2 ? phv_data_202 : _GEN_4819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4821 = 8'hcb == local_offset_2 ? phv_data_203 : _GEN_4820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4822 = 8'hcc == local_offset_2 ? phv_data_204 : _GEN_4821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4823 = 8'hcd == local_offset_2 ? phv_data_205 : _GEN_4822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4824 = 8'hce == local_offset_2 ? phv_data_206 : _GEN_4823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4825 = 8'hcf == local_offset_2 ? phv_data_207 : _GEN_4824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4826 = 8'hd0 == local_offset_2 ? phv_data_208 : _GEN_4825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4827 = 8'hd1 == local_offset_2 ? phv_data_209 : _GEN_4826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4828 = 8'hd2 == local_offset_2 ? phv_data_210 : _GEN_4827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4829 = 8'hd3 == local_offset_2 ? phv_data_211 : _GEN_4828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4830 = 8'hd4 == local_offset_2 ? phv_data_212 : _GEN_4829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4831 = 8'hd5 == local_offset_2 ? phv_data_213 : _GEN_4830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4832 = 8'hd6 == local_offset_2 ? phv_data_214 : _GEN_4831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4833 = 8'hd7 == local_offset_2 ? phv_data_215 : _GEN_4832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4834 = 8'hd8 == local_offset_2 ? phv_data_216 : _GEN_4833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4835 = 8'hd9 == local_offset_2 ? phv_data_217 : _GEN_4834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4836 = 8'hda == local_offset_2 ? phv_data_218 : _GEN_4835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4837 = 8'hdb == local_offset_2 ? phv_data_219 : _GEN_4836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4838 = 8'hdc == local_offset_2 ? phv_data_220 : _GEN_4837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4839 = 8'hdd == local_offset_2 ? phv_data_221 : _GEN_4838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4840 = 8'hde == local_offset_2 ? phv_data_222 : _GEN_4839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4841 = 8'hdf == local_offset_2 ? phv_data_223 : _GEN_4840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4842 = 8'he0 == local_offset_2 ? phv_data_224 : _GEN_4841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4843 = 8'he1 == local_offset_2 ? phv_data_225 : _GEN_4842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4844 = 8'he2 == local_offset_2 ? phv_data_226 : _GEN_4843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4845 = 8'he3 == local_offset_2 ? phv_data_227 : _GEN_4844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4846 = 8'he4 == local_offset_2 ? phv_data_228 : _GEN_4845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4847 = 8'he5 == local_offset_2 ? phv_data_229 : _GEN_4846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4848 = 8'he6 == local_offset_2 ? phv_data_230 : _GEN_4847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4849 = 8'he7 == local_offset_2 ? phv_data_231 : _GEN_4848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4850 = 8'he8 == local_offset_2 ? phv_data_232 : _GEN_4849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4851 = 8'he9 == local_offset_2 ? phv_data_233 : _GEN_4850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4852 = 8'hea == local_offset_2 ? phv_data_234 : _GEN_4851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4853 = 8'heb == local_offset_2 ? phv_data_235 : _GEN_4852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4854 = 8'hec == local_offset_2 ? phv_data_236 : _GEN_4853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4855 = 8'hed == local_offset_2 ? phv_data_237 : _GEN_4854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4856 = 8'hee == local_offset_2 ? phv_data_238 : _GEN_4855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4857 = 8'hef == local_offset_2 ? phv_data_239 : _GEN_4856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4858 = 8'hf0 == local_offset_2 ? phv_data_240 : _GEN_4857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4859 = 8'hf1 == local_offset_2 ? phv_data_241 : _GEN_4858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4860 = 8'hf2 == local_offset_2 ? phv_data_242 : _GEN_4859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4861 = 8'hf3 == local_offset_2 ? phv_data_243 : _GEN_4860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4862 = 8'hf4 == local_offset_2 ? phv_data_244 : _GEN_4861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4863 = 8'hf5 == local_offset_2 ? phv_data_245 : _GEN_4862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4864 = 8'hf6 == local_offset_2 ? phv_data_246 : _GEN_4863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4865 = 8'hf7 == local_offset_2 ? phv_data_247 : _GEN_4864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4866 = 8'hf8 == local_offset_2 ? phv_data_248 : _GEN_4865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4867 = 8'hf9 == local_offset_2 ? phv_data_249 : _GEN_4866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4868 = 8'hfa == local_offset_2 ? phv_data_250 : _GEN_4867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4869 = 8'hfb == local_offset_2 ? phv_data_251 : _GEN_4868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4870 = 8'hfc == local_offset_2 ? phv_data_252 : _GEN_4869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4871 = 8'hfd == local_offset_2 ? phv_data_253 : _GEN_4870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4872 = 8'hfe == local_offset_2 ? phv_data_254 : _GEN_4871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4873 = 8'hff == local_offset_2 ? phv_data_255 : _GEN_4872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_14630 = {{1'd0}, local_offset_2}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4874 = 9'h100 == _GEN_14630 ? phv_data_256 : _GEN_4873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4875 = 9'h101 == _GEN_14630 ? phv_data_257 : _GEN_4874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4876 = 9'h102 == _GEN_14630 ? phv_data_258 : _GEN_4875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4877 = 9'h103 == _GEN_14630 ? phv_data_259 : _GEN_4876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4878 = 9'h104 == _GEN_14630 ? phv_data_260 : _GEN_4877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4879 = 9'h105 == _GEN_14630 ? phv_data_261 : _GEN_4878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4880 = 9'h106 == _GEN_14630 ? phv_data_262 : _GEN_4879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4881 = 9'h107 == _GEN_14630 ? phv_data_263 : _GEN_4880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4882 = 9'h108 == _GEN_14630 ? phv_data_264 : _GEN_4881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4883 = 9'h109 == _GEN_14630 ? phv_data_265 : _GEN_4882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4884 = 9'h10a == _GEN_14630 ? phv_data_266 : _GEN_4883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4885 = 9'h10b == _GEN_14630 ? phv_data_267 : _GEN_4884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4886 = 9'h10c == _GEN_14630 ? phv_data_268 : _GEN_4885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4887 = 9'h10d == _GEN_14630 ? phv_data_269 : _GEN_4886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4888 = 9'h10e == _GEN_14630 ? phv_data_270 : _GEN_4887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4889 = 9'h10f == _GEN_14630 ? phv_data_271 : _GEN_4888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4890 = 9'h110 == _GEN_14630 ? phv_data_272 : _GEN_4889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4891 = 9'h111 == _GEN_14630 ? phv_data_273 : _GEN_4890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4892 = 9'h112 == _GEN_14630 ? phv_data_274 : _GEN_4891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4893 = 9'h113 == _GEN_14630 ? phv_data_275 : _GEN_4892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4894 = 9'h114 == _GEN_14630 ? phv_data_276 : _GEN_4893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4895 = 9'h115 == _GEN_14630 ? phv_data_277 : _GEN_4894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4896 = 9'h116 == _GEN_14630 ? phv_data_278 : _GEN_4895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4897 = 9'h117 == _GEN_14630 ? phv_data_279 : _GEN_4896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4898 = 9'h118 == _GEN_14630 ? phv_data_280 : _GEN_4897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4899 = 9'h119 == _GEN_14630 ? phv_data_281 : _GEN_4898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4900 = 9'h11a == _GEN_14630 ? phv_data_282 : _GEN_4899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4901 = 9'h11b == _GEN_14630 ? phv_data_283 : _GEN_4900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4902 = 9'h11c == _GEN_14630 ? phv_data_284 : _GEN_4901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4903 = 9'h11d == _GEN_14630 ? phv_data_285 : _GEN_4902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4904 = 9'h11e == _GEN_14630 ? phv_data_286 : _GEN_4903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4905 = 9'h11f == _GEN_14630 ? phv_data_287 : _GEN_4904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4906 = 9'h120 == _GEN_14630 ? phv_data_288 : _GEN_4905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4907 = 9'h121 == _GEN_14630 ? phv_data_289 : _GEN_4906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4908 = 9'h122 == _GEN_14630 ? phv_data_290 : _GEN_4907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4909 = 9'h123 == _GEN_14630 ? phv_data_291 : _GEN_4908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4910 = 9'h124 == _GEN_14630 ? phv_data_292 : _GEN_4909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4911 = 9'h125 == _GEN_14630 ? phv_data_293 : _GEN_4910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4912 = 9'h126 == _GEN_14630 ? phv_data_294 : _GEN_4911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4913 = 9'h127 == _GEN_14630 ? phv_data_295 : _GEN_4912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4914 = 9'h128 == _GEN_14630 ? phv_data_296 : _GEN_4913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4915 = 9'h129 == _GEN_14630 ? phv_data_297 : _GEN_4914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4916 = 9'h12a == _GEN_14630 ? phv_data_298 : _GEN_4915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4917 = 9'h12b == _GEN_14630 ? phv_data_299 : _GEN_4916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4918 = 9'h12c == _GEN_14630 ? phv_data_300 : _GEN_4917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4919 = 9'h12d == _GEN_14630 ? phv_data_301 : _GEN_4918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4920 = 9'h12e == _GEN_14630 ? phv_data_302 : _GEN_4919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4921 = 9'h12f == _GEN_14630 ? phv_data_303 : _GEN_4920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4922 = 9'h130 == _GEN_14630 ? phv_data_304 : _GEN_4921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4923 = 9'h131 == _GEN_14630 ? phv_data_305 : _GEN_4922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4924 = 9'h132 == _GEN_14630 ? phv_data_306 : _GEN_4923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4925 = 9'h133 == _GEN_14630 ? phv_data_307 : _GEN_4924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4926 = 9'h134 == _GEN_14630 ? phv_data_308 : _GEN_4925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4927 = 9'h135 == _GEN_14630 ? phv_data_309 : _GEN_4926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4928 = 9'h136 == _GEN_14630 ? phv_data_310 : _GEN_4927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4929 = 9'h137 == _GEN_14630 ? phv_data_311 : _GEN_4928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4930 = 9'h138 == _GEN_14630 ? phv_data_312 : _GEN_4929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4931 = 9'h139 == _GEN_14630 ? phv_data_313 : _GEN_4930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4932 = 9'h13a == _GEN_14630 ? phv_data_314 : _GEN_4931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4933 = 9'h13b == _GEN_14630 ? phv_data_315 : _GEN_4932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4934 = 9'h13c == _GEN_14630 ? phv_data_316 : _GEN_4933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4935 = 9'h13d == _GEN_14630 ? phv_data_317 : _GEN_4934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4936 = 9'h13e == _GEN_14630 ? phv_data_318 : _GEN_4935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4937 = 9'h13f == _GEN_14630 ? phv_data_319 : _GEN_4936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4938 = 9'h140 == _GEN_14630 ? phv_data_320 : _GEN_4937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4939 = 9'h141 == _GEN_14630 ? phv_data_321 : _GEN_4938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4940 = 9'h142 == _GEN_14630 ? phv_data_322 : _GEN_4939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4941 = 9'h143 == _GEN_14630 ? phv_data_323 : _GEN_4940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4942 = 9'h144 == _GEN_14630 ? phv_data_324 : _GEN_4941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4943 = 9'h145 == _GEN_14630 ? phv_data_325 : _GEN_4942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4944 = 9'h146 == _GEN_14630 ? phv_data_326 : _GEN_4943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4945 = 9'h147 == _GEN_14630 ? phv_data_327 : _GEN_4944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4946 = 9'h148 == _GEN_14630 ? phv_data_328 : _GEN_4945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4947 = 9'h149 == _GEN_14630 ? phv_data_329 : _GEN_4946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4948 = 9'h14a == _GEN_14630 ? phv_data_330 : _GEN_4947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4949 = 9'h14b == _GEN_14630 ? phv_data_331 : _GEN_4948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4950 = 9'h14c == _GEN_14630 ? phv_data_332 : _GEN_4949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4951 = 9'h14d == _GEN_14630 ? phv_data_333 : _GEN_4950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4952 = 9'h14e == _GEN_14630 ? phv_data_334 : _GEN_4951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4953 = 9'h14f == _GEN_14630 ? phv_data_335 : _GEN_4952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4954 = 9'h150 == _GEN_14630 ? phv_data_336 : _GEN_4953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4955 = 9'h151 == _GEN_14630 ? phv_data_337 : _GEN_4954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4956 = 9'h152 == _GEN_14630 ? phv_data_338 : _GEN_4955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4957 = 9'h153 == _GEN_14630 ? phv_data_339 : _GEN_4956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4958 = 9'h154 == _GEN_14630 ? phv_data_340 : _GEN_4957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4959 = 9'h155 == _GEN_14630 ? phv_data_341 : _GEN_4958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4960 = 9'h156 == _GEN_14630 ? phv_data_342 : _GEN_4959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4961 = 9'h157 == _GEN_14630 ? phv_data_343 : _GEN_4960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4962 = 9'h158 == _GEN_14630 ? phv_data_344 : _GEN_4961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4963 = 9'h159 == _GEN_14630 ? phv_data_345 : _GEN_4962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4964 = 9'h15a == _GEN_14630 ? phv_data_346 : _GEN_4963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4965 = 9'h15b == _GEN_14630 ? phv_data_347 : _GEN_4964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4966 = 9'h15c == _GEN_14630 ? phv_data_348 : _GEN_4965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4967 = 9'h15d == _GEN_14630 ? phv_data_349 : _GEN_4966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4968 = 9'h15e == _GEN_14630 ? phv_data_350 : _GEN_4967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4969 = 9'h15f == _GEN_14630 ? phv_data_351 : _GEN_4968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4970 = 9'h160 == _GEN_14630 ? phv_data_352 : _GEN_4969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4971 = 9'h161 == _GEN_14630 ? phv_data_353 : _GEN_4970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4972 = 9'h162 == _GEN_14630 ? phv_data_354 : _GEN_4971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4973 = 9'h163 == _GEN_14630 ? phv_data_355 : _GEN_4972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4974 = 9'h164 == _GEN_14630 ? phv_data_356 : _GEN_4973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4975 = 9'h165 == _GEN_14630 ? phv_data_357 : _GEN_4974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4976 = 9'h166 == _GEN_14630 ? phv_data_358 : _GEN_4975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4977 = 9'h167 == _GEN_14630 ? phv_data_359 : _GEN_4976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4978 = 9'h168 == _GEN_14630 ? phv_data_360 : _GEN_4977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4979 = 9'h169 == _GEN_14630 ? phv_data_361 : _GEN_4978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4980 = 9'h16a == _GEN_14630 ? phv_data_362 : _GEN_4979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4981 = 9'h16b == _GEN_14630 ? phv_data_363 : _GEN_4980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4982 = 9'h16c == _GEN_14630 ? phv_data_364 : _GEN_4981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4983 = 9'h16d == _GEN_14630 ? phv_data_365 : _GEN_4982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4984 = 9'h16e == _GEN_14630 ? phv_data_366 : _GEN_4983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4985 = 9'h16f == _GEN_14630 ? phv_data_367 : _GEN_4984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4986 = 9'h170 == _GEN_14630 ? phv_data_368 : _GEN_4985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4987 = 9'h171 == _GEN_14630 ? phv_data_369 : _GEN_4986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4988 = 9'h172 == _GEN_14630 ? phv_data_370 : _GEN_4987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4989 = 9'h173 == _GEN_14630 ? phv_data_371 : _GEN_4988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4990 = 9'h174 == _GEN_14630 ? phv_data_372 : _GEN_4989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4991 = 9'h175 == _GEN_14630 ? phv_data_373 : _GEN_4990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4992 = 9'h176 == _GEN_14630 ? phv_data_374 : _GEN_4991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4993 = 9'h177 == _GEN_14630 ? phv_data_375 : _GEN_4992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4994 = 9'h178 == _GEN_14630 ? phv_data_376 : _GEN_4993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4995 = 9'h179 == _GEN_14630 ? phv_data_377 : _GEN_4994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4996 = 9'h17a == _GEN_14630 ? phv_data_378 : _GEN_4995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4997 = 9'h17b == _GEN_14630 ? phv_data_379 : _GEN_4996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4998 = 9'h17c == _GEN_14630 ? phv_data_380 : _GEN_4997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4999 = 9'h17d == _GEN_14630 ? phv_data_381 : _GEN_4998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5000 = 9'h17e == _GEN_14630 ? phv_data_382 : _GEN_4999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5001 = 9'h17f == _GEN_14630 ? phv_data_383 : _GEN_5000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5002 = 9'h180 == _GEN_14630 ? phv_data_384 : _GEN_5001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5003 = 9'h181 == _GEN_14630 ? phv_data_385 : _GEN_5002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5004 = 9'h182 == _GEN_14630 ? phv_data_386 : _GEN_5003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5005 = 9'h183 == _GEN_14630 ? phv_data_387 : _GEN_5004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5006 = 9'h184 == _GEN_14630 ? phv_data_388 : _GEN_5005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5007 = 9'h185 == _GEN_14630 ? phv_data_389 : _GEN_5006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5008 = 9'h186 == _GEN_14630 ? phv_data_390 : _GEN_5007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5009 = 9'h187 == _GEN_14630 ? phv_data_391 : _GEN_5008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5010 = 9'h188 == _GEN_14630 ? phv_data_392 : _GEN_5009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5011 = 9'h189 == _GEN_14630 ? phv_data_393 : _GEN_5010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5012 = 9'h18a == _GEN_14630 ? phv_data_394 : _GEN_5011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5013 = 9'h18b == _GEN_14630 ? phv_data_395 : _GEN_5012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5014 = 9'h18c == _GEN_14630 ? phv_data_396 : _GEN_5013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5015 = 9'h18d == _GEN_14630 ? phv_data_397 : _GEN_5014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5016 = 9'h18e == _GEN_14630 ? phv_data_398 : _GEN_5015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5017 = 9'h18f == _GEN_14630 ? phv_data_399 : _GEN_5016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5018 = 9'h190 == _GEN_14630 ? phv_data_400 : _GEN_5017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5019 = 9'h191 == _GEN_14630 ? phv_data_401 : _GEN_5018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5020 = 9'h192 == _GEN_14630 ? phv_data_402 : _GEN_5019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5021 = 9'h193 == _GEN_14630 ? phv_data_403 : _GEN_5020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5022 = 9'h194 == _GEN_14630 ? phv_data_404 : _GEN_5021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5023 = 9'h195 == _GEN_14630 ? phv_data_405 : _GEN_5022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5024 = 9'h196 == _GEN_14630 ? phv_data_406 : _GEN_5023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5025 = 9'h197 == _GEN_14630 ? phv_data_407 : _GEN_5024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5026 = 9'h198 == _GEN_14630 ? phv_data_408 : _GEN_5025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5027 = 9'h199 == _GEN_14630 ? phv_data_409 : _GEN_5026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5028 = 9'h19a == _GEN_14630 ? phv_data_410 : _GEN_5027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5029 = 9'h19b == _GEN_14630 ? phv_data_411 : _GEN_5028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5030 = 9'h19c == _GEN_14630 ? phv_data_412 : _GEN_5029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5031 = 9'h19d == _GEN_14630 ? phv_data_413 : _GEN_5030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5032 = 9'h19e == _GEN_14630 ? phv_data_414 : _GEN_5031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5033 = 9'h19f == _GEN_14630 ? phv_data_415 : _GEN_5032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5034 = 9'h1a0 == _GEN_14630 ? phv_data_416 : _GEN_5033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5035 = 9'h1a1 == _GEN_14630 ? phv_data_417 : _GEN_5034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5036 = 9'h1a2 == _GEN_14630 ? phv_data_418 : _GEN_5035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5037 = 9'h1a3 == _GEN_14630 ? phv_data_419 : _GEN_5036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5038 = 9'h1a4 == _GEN_14630 ? phv_data_420 : _GEN_5037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5039 = 9'h1a5 == _GEN_14630 ? phv_data_421 : _GEN_5038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5040 = 9'h1a6 == _GEN_14630 ? phv_data_422 : _GEN_5039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5041 = 9'h1a7 == _GEN_14630 ? phv_data_423 : _GEN_5040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5042 = 9'h1a8 == _GEN_14630 ? phv_data_424 : _GEN_5041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5043 = 9'h1a9 == _GEN_14630 ? phv_data_425 : _GEN_5042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5044 = 9'h1aa == _GEN_14630 ? phv_data_426 : _GEN_5043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5045 = 9'h1ab == _GEN_14630 ? phv_data_427 : _GEN_5044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5046 = 9'h1ac == _GEN_14630 ? phv_data_428 : _GEN_5045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5047 = 9'h1ad == _GEN_14630 ? phv_data_429 : _GEN_5046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5048 = 9'h1ae == _GEN_14630 ? phv_data_430 : _GEN_5047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5049 = 9'h1af == _GEN_14630 ? phv_data_431 : _GEN_5048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5050 = 9'h1b0 == _GEN_14630 ? phv_data_432 : _GEN_5049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5051 = 9'h1b1 == _GEN_14630 ? phv_data_433 : _GEN_5050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5052 = 9'h1b2 == _GEN_14630 ? phv_data_434 : _GEN_5051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5053 = 9'h1b3 == _GEN_14630 ? phv_data_435 : _GEN_5052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5054 = 9'h1b4 == _GEN_14630 ? phv_data_436 : _GEN_5053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5055 = 9'h1b5 == _GEN_14630 ? phv_data_437 : _GEN_5054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5056 = 9'h1b6 == _GEN_14630 ? phv_data_438 : _GEN_5055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5057 = 9'h1b7 == _GEN_14630 ? phv_data_439 : _GEN_5056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5058 = 9'h1b8 == _GEN_14630 ? phv_data_440 : _GEN_5057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5059 = 9'h1b9 == _GEN_14630 ? phv_data_441 : _GEN_5058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5060 = 9'h1ba == _GEN_14630 ? phv_data_442 : _GEN_5059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5061 = 9'h1bb == _GEN_14630 ? phv_data_443 : _GEN_5060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5062 = 9'h1bc == _GEN_14630 ? phv_data_444 : _GEN_5061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5063 = 9'h1bd == _GEN_14630 ? phv_data_445 : _GEN_5062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5064 = 9'h1be == _GEN_14630 ? phv_data_446 : _GEN_5063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5065 = 9'h1bf == _GEN_14630 ? phv_data_447 : _GEN_5064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5066 = 9'h1c0 == _GEN_14630 ? phv_data_448 : _GEN_5065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5067 = 9'h1c1 == _GEN_14630 ? phv_data_449 : _GEN_5066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5068 = 9'h1c2 == _GEN_14630 ? phv_data_450 : _GEN_5067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5069 = 9'h1c3 == _GEN_14630 ? phv_data_451 : _GEN_5068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5070 = 9'h1c4 == _GEN_14630 ? phv_data_452 : _GEN_5069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5071 = 9'h1c5 == _GEN_14630 ? phv_data_453 : _GEN_5070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5072 = 9'h1c6 == _GEN_14630 ? phv_data_454 : _GEN_5071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5073 = 9'h1c7 == _GEN_14630 ? phv_data_455 : _GEN_5072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5074 = 9'h1c8 == _GEN_14630 ? phv_data_456 : _GEN_5073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5075 = 9'h1c9 == _GEN_14630 ? phv_data_457 : _GEN_5074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5076 = 9'h1ca == _GEN_14630 ? phv_data_458 : _GEN_5075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5077 = 9'h1cb == _GEN_14630 ? phv_data_459 : _GEN_5076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5078 = 9'h1cc == _GEN_14630 ? phv_data_460 : _GEN_5077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5079 = 9'h1cd == _GEN_14630 ? phv_data_461 : _GEN_5078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5080 = 9'h1ce == _GEN_14630 ? phv_data_462 : _GEN_5079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5081 = 9'h1cf == _GEN_14630 ? phv_data_463 : _GEN_5080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5082 = 9'h1d0 == _GEN_14630 ? phv_data_464 : _GEN_5081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5083 = 9'h1d1 == _GEN_14630 ? phv_data_465 : _GEN_5082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5084 = 9'h1d2 == _GEN_14630 ? phv_data_466 : _GEN_5083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5085 = 9'h1d3 == _GEN_14630 ? phv_data_467 : _GEN_5084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5086 = 9'h1d4 == _GEN_14630 ? phv_data_468 : _GEN_5085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5087 = 9'h1d5 == _GEN_14630 ? phv_data_469 : _GEN_5086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5088 = 9'h1d6 == _GEN_14630 ? phv_data_470 : _GEN_5087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5089 = 9'h1d7 == _GEN_14630 ? phv_data_471 : _GEN_5088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5090 = 9'h1d8 == _GEN_14630 ? phv_data_472 : _GEN_5089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5091 = 9'h1d9 == _GEN_14630 ? phv_data_473 : _GEN_5090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5092 = 9'h1da == _GEN_14630 ? phv_data_474 : _GEN_5091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5093 = 9'h1db == _GEN_14630 ? phv_data_475 : _GEN_5092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5094 = 9'h1dc == _GEN_14630 ? phv_data_476 : _GEN_5093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5095 = 9'h1dd == _GEN_14630 ? phv_data_477 : _GEN_5094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5096 = 9'h1de == _GEN_14630 ? phv_data_478 : _GEN_5095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5097 = 9'h1df == _GEN_14630 ? phv_data_479 : _GEN_5096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5098 = 9'h1e0 == _GEN_14630 ? phv_data_480 : _GEN_5097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5099 = 9'h1e1 == _GEN_14630 ? phv_data_481 : _GEN_5098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5100 = 9'h1e2 == _GEN_14630 ? phv_data_482 : _GEN_5099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5101 = 9'h1e3 == _GEN_14630 ? phv_data_483 : _GEN_5100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5102 = 9'h1e4 == _GEN_14630 ? phv_data_484 : _GEN_5101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5103 = 9'h1e5 == _GEN_14630 ? phv_data_485 : _GEN_5102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5104 = 9'h1e6 == _GEN_14630 ? phv_data_486 : _GEN_5103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5105 = 9'h1e7 == _GEN_14630 ? phv_data_487 : _GEN_5104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5106 = 9'h1e8 == _GEN_14630 ? phv_data_488 : _GEN_5105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5107 = 9'h1e9 == _GEN_14630 ? phv_data_489 : _GEN_5106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5108 = 9'h1ea == _GEN_14630 ? phv_data_490 : _GEN_5107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5109 = 9'h1eb == _GEN_14630 ? phv_data_491 : _GEN_5108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5110 = 9'h1ec == _GEN_14630 ? phv_data_492 : _GEN_5109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5111 = 9'h1ed == _GEN_14630 ? phv_data_493 : _GEN_5110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5112 = 9'h1ee == _GEN_14630 ? phv_data_494 : _GEN_5111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5113 = 9'h1ef == _GEN_14630 ? phv_data_495 : _GEN_5112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5114 = 9'h1f0 == _GEN_14630 ? phv_data_496 : _GEN_5113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5115 = 9'h1f1 == _GEN_14630 ? phv_data_497 : _GEN_5114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5116 = 9'h1f2 == _GEN_14630 ? phv_data_498 : _GEN_5115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5117 = 9'h1f3 == _GEN_14630 ? phv_data_499 : _GEN_5116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5118 = 9'h1f4 == _GEN_14630 ? phv_data_500 : _GEN_5117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5119 = 9'h1f5 == _GEN_14630 ? phv_data_501 : _GEN_5118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5120 = 9'h1f6 == _GEN_14630 ? phv_data_502 : _GEN_5119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5121 = 9'h1f7 == _GEN_14630 ? phv_data_503 : _GEN_5120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5122 = 9'h1f8 == _GEN_14630 ? phv_data_504 : _GEN_5121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5123 = 9'h1f9 == _GEN_14630 ? phv_data_505 : _GEN_5122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5124 = 9'h1fa == _GEN_14630 ? phv_data_506 : _GEN_5123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5125 = 9'h1fb == _GEN_14630 ? phv_data_507 : _GEN_5124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5126 = 9'h1fc == _GEN_14630 ? phv_data_508 : _GEN_5125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5127 = 9'h1fd == _GEN_14630 ? phv_data_509 : _GEN_5126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5128 = 9'h1fe == _GEN_14630 ? phv_data_510 : _GEN_5127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5129 = 9'h1ff == _GEN_14630 ? phv_data_511 : _GEN_5128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5131 = 8'h1 == _match_key_qbytes_2_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5132 = 8'h2 == _match_key_qbytes_2_T ? phv_data_2 : _GEN_5131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5133 = 8'h3 == _match_key_qbytes_2_T ? phv_data_3 : _GEN_5132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5134 = 8'h4 == _match_key_qbytes_2_T ? phv_data_4 : _GEN_5133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5135 = 8'h5 == _match_key_qbytes_2_T ? phv_data_5 : _GEN_5134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5136 = 8'h6 == _match_key_qbytes_2_T ? phv_data_6 : _GEN_5135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5137 = 8'h7 == _match_key_qbytes_2_T ? phv_data_7 : _GEN_5136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5138 = 8'h8 == _match_key_qbytes_2_T ? phv_data_8 : _GEN_5137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5139 = 8'h9 == _match_key_qbytes_2_T ? phv_data_9 : _GEN_5138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5140 = 8'ha == _match_key_qbytes_2_T ? phv_data_10 : _GEN_5139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5141 = 8'hb == _match_key_qbytes_2_T ? phv_data_11 : _GEN_5140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5142 = 8'hc == _match_key_qbytes_2_T ? phv_data_12 : _GEN_5141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5143 = 8'hd == _match_key_qbytes_2_T ? phv_data_13 : _GEN_5142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5144 = 8'he == _match_key_qbytes_2_T ? phv_data_14 : _GEN_5143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5145 = 8'hf == _match_key_qbytes_2_T ? phv_data_15 : _GEN_5144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5146 = 8'h10 == _match_key_qbytes_2_T ? phv_data_16 : _GEN_5145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5147 = 8'h11 == _match_key_qbytes_2_T ? phv_data_17 : _GEN_5146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5148 = 8'h12 == _match_key_qbytes_2_T ? phv_data_18 : _GEN_5147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5149 = 8'h13 == _match_key_qbytes_2_T ? phv_data_19 : _GEN_5148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5150 = 8'h14 == _match_key_qbytes_2_T ? phv_data_20 : _GEN_5149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5151 = 8'h15 == _match_key_qbytes_2_T ? phv_data_21 : _GEN_5150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5152 = 8'h16 == _match_key_qbytes_2_T ? phv_data_22 : _GEN_5151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5153 = 8'h17 == _match_key_qbytes_2_T ? phv_data_23 : _GEN_5152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5154 = 8'h18 == _match_key_qbytes_2_T ? phv_data_24 : _GEN_5153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5155 = 8'h19 == _match_key_qbytes_2_T ? phv_data_25 : _GEN_5154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5156 = 8'h1a == _match_key_qbytes_2_T ? phv_data_26 : _GEN_5155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5157 = 8'h1b == _match_key_qbytes_2_T ? phv_data_27 : _GEN_5156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5158 = 8'h1c == _match_key_qbytes_2_T ? phv_data_28 : _GEN_5157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5159 = 8'h1d == _match_key_qbytes_2_T ? phv_data_29 : _GEN_5158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5160 = 8'h1e == _match_key_qbytes_2_T ? phv_data_30 : _GEN_5159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5161 = 8'h1f == _match_key_qbytes_2_T ? phv_data_31 : _GEN_5160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5162 = 8'h20 == _match_key_qbytes_2_T ? phv_data_32 : _GEN_5161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5163 = 8'h21 == _match_key_qbytes_2_T ? phv_data_33 : _GEN_5162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5164 = 8'h22 == _match_key_qbytes_2_T ? phv_data_34 : _GEN_5163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5165 = 8'h23 == _match_key_qbytes_2_T ? phv_data_35 : _GEN_5164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5166 = 8'h24 == _match_key_qbytes_2_T ? phv_data_36 : _GEN_5165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5167 = 8'h25 == _match_key_qbytes_2_T ? phv_data_37 : _GEN_5166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5168 = 8'h26 == _match_key_qbytes_2_T ? phv_data_38 : _GEN_5167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5169 = 8'h27 == _match_key_qbytes_2_T ? phv_data_39 : _GEN_5168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5170 = 8'h28 == _match_key_qbytes_2_T ? phv_data_40 : _GEN_5169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5171 = 8'h29 == _match_key_qbytes_2_T ? phv_data_41 : _GEN_5170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5172 = 8'h2a == _match_key_qbytes_2_T ? phv_data_42 : _GEN_5171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5173 = 8'h2b == _match_key_qbytes_2_T ? phv_data_43 : _GEN_5172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5174 = 8'h2c == _match_key_qbytes_2_T ? phv_data_44 : _GEN_5173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5175 = 8'h2d == _match_key_qbytes_2_T ? phv_data_45 : _GEN_5174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5176 = 8'h2e == _match_key_qbytes_2_T ? phv_data_46 : _GEN_5175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5177 = 8'h2f == _match_key_qbytes_2_T ? phv_data_47 : _GEN_5176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5178 = 8'h30 == _match_key_qbytes_2_T ? phv_data_48 : _GEN_5177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5179 = 8'h31 == _match_key_qbytes_2_T ? phv_data_49 : _GEN_5178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5180 = 8'h32 == _match_key_qbytes_2_T ? phv_data_50 : _GEN_5179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5181 = 8'h33 == _match_key_qbytes_2_T ? phv_data_51 : _GEN_5180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5182 = 8'h34 == _match_key_qbytes_2_T ? phv_data_52 : _GEN_5181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5183 = 8'h35 == _match_key_qbytes_2_T ? phv_data_53 : _GEN_5182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5184 = 8'h36 == _match_key_qbytes_2_T ? phv_data_54 : _GEN_5183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5185 = 8'h37 == _match_key_qbytes_2_T ? phv_data_55 : _GEN_5184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5186 = 8'h38 == _match_key_qbytes_2_T ? phv_data_56 : _GEN_5185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5187 = 8'h39 == _match_key_qbytes_2_T ? phv_data_57 : _GEN_5186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5188 = 8'h3a == _match_key_qbytes_2_T ? phv_data_58 : _GEN_5187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5189 = 8'h3b == _match_key_qbytes_2_T ? phv_data_59 : _GEN_5188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5190 = 8'h3c == _match_key_qbytes_2_T ? phv_data_60 : _GEN_5189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5191 = 8'h3d == _match_key_qbytes_2_T ? phv_data_61 : _GEN_5190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5192 = 8'h3e == _match_key_qbytes_2_T ? phv_data_62 : _GEN_5191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5193 = 8'h3f == _match_key_qbytes_2_T ? phv_data_63 : _GEN_5192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5194 = 8'h40 == _match_key_qbytes_2_T ? phv_data_64 : _GEN_5193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5195 = 8'h41 == _match_key_qbytes_2_T ? phv_data_65 : _GEN_5194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5196 = 8'h42 == _match_key_qbytes_2_T ? phv_data_66 : _GEN_5195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5197 = 8'h43 == _match_key_qbytes_2_T ? phv_data_67 : _GEN_5196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5198 = 8'h44 == _match_key_qbytes_2_T ? phv_data_68 : _GEN_5197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5199 = 8'h45 == _match_key_qbytes_2_T ? phv_data_69 : _GEN_5198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5200 = 8'h46 == _match_key_qbytes_2_T ? phv_data_70 : _GEN_5199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5201 = 8'h47 == _match_key_qbytes_2_T ? phv_data_71 : _GEN_5200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5202 = 8'h48 == _match_key_qbytes_2_T ? phv_data_72 : _GEN_5201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5203 = 8'h49 == _match_key_qbytes_2_T ? phv_data_73 : _GEN_5202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5204 = 8'h4a == _match_key_qbytes_2_T ? phv_data_74 : _GEN_5203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5205 = 8'h4b == _match_key_qbytes_2_T ? phv_data_75 : _GEN_5204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5206 = 8'h4c == _match_key_qbytes_2_T ? phv_data_76 : _GEN_5205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5207 = 8'h4d == _match_key_qbytes_2_T ? phv_data_77 : _GEN_5206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5208 = 8'h4e == _match_key_qbytes_2_T ? phv_data_78 : _GEN_5207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5209 = 8'h4f == _match_key_qbytes_2_T ? phv_data_79 : _GEN_5208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5210 = 8'h50 == _match_key_qbytes_2_T ? phv_data_80 : _GEN_5209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5211 = 8'h51 == _match_key_qbytes_2_T ? phv_data_81 : _GEN_5210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5212 = 8'h52 == _match_key_qbytes_2_T ? phv_data_82 : _GEN_5211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5213 = 8'h53 == _match_key_qbytes_2_T ? phv_data_83 : _GEN_5212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5214 = 8'h54 == _match_key_qbytes_2_T ? phv_data_84 : _GEN_5213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5215 = 8'h55 == _match_key_qbytes_2_T ? phv_data_85 : _GEN_5214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5216 = 8'h56 == _match_key_qbytes_2_T ? phv_data_86 : _GEN_5215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5217 = 8'h57 == _match_key_qbytes_2_T ? phv_data_87 : _GEN_5216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5218 = 8'h58 == _match_key_qbytes_2_T ? phv_data_88 : _GEN_5217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5219 = 8'h59 == _match_key_qbytes_2_T ? phv_data_89 : _GEN_5218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5220 = 8'h5a == _match_key_qbytes_2_T ? phv_data_90 : _GEN_5219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5221 = 8'h5b == _match_key_qbytes_2_T ? phv_data_91 : _GEN_5220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5222 = 8'h5c == _match_key_qbytes_2_T ? phv_data_92 : _GEN_5221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5223 = 8'h5d == _match_key_qbytes_2_T ? phv_data_93 : _GEN_5222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5224 = 8'h5e == _match_key_qbytes_2_T ? phv_data_94 : _GEN_5223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5225 = 8'h5f == _match_key_qbytes_2_T ? phv_data_95 : _GEN_5224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5226 = 8'h60 == _match_key_qbytes_2_T ? phv_data_96 : _GEN_5225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5227 = 8'h61 == _match_key_qbytes_2_T ? phv_data_97 : _GEN_5226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5228 = 8'h62 == _match_key_qbytes_2_T ? phv_data_98 : _GEN_5227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5229 = 8'h63 == _match_key_qbytes_2_T ? phv_data_99 : _GEN_5228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5230 = 8'h64 == _match_key_qbytes_2_T ? phv_data_100 : _GEN_5229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5231 = 8'h65 == _match_key_qbytes_2_T ? phv_data_101 : _GEN_5230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5232 = 8'h66 == _match_key_qbytes_2_T ? phv_data_102 : _GEN_5231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5233 = 8'h67 == _match_key_qbytes_2_T ? phv_data_103 : _GEN_5232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5234 = 8'h68 == _match_key_qbytes_2_T ? phv_data_104 : _GEN_5233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5235 = 8'h69 == _match_key_qbytes_2_T ? phv_data_105 : _GEN_5234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5236 = 8'h6a == _match_key_qbytes_2_T ? phv_data_106 : _GEN_5235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5237 = 8'h6b == _match_key_qbytes_2_T ? phv_data_107 : _GEN_5236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5238 = 8'h6c == _match_key_qbytes_2_T ? phv_data_108 : _GEN_5237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5239 = 8'h6d == _match_key_qbytes_2_T ? phv_data_109 : _GEN_5238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5240 = 8'h6e == _match_key_qbytes_2_T ? phv_data_110 : _GEN_5239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5241 = 8'h6f == _match_key_qbytes_2_T ? phv_data_111 : _GEN_5240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5242 = 8'h70 == _match_key_qbytes_2_T ? phv_data_112 : _GEN_5241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5243 = 8'h71 == _match_key_qbytes_2_T ? phv_data_113 : _GEN_5242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5244 = 8'h72 == _match_key_qbytes_2_T ? phv_data_114 : _GEN_5243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5245 = 8'h73 == _match_key_qbytes_2_T ? phv_data_115 : _GEN_5244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5246 = 8'h74 == _match_key_qbytes_2_T ? phv_data_116 : _GEN_5245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5247 = 8'h75 == _match_key_qbytes_2_T ? phv_data_117 : _GEN_5246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5248 = 8'h76 == _match_key_qbytes_2_T ? phv_data_118 : _GEN_5247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5249 = 8'h77 == _match_key_qbytes_2_T ? phv_data_119 : _GEN_5248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5250 = 8'h78 == _match_key_qbytes_2_T ? phv_data_120 : _GEN_5249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5251 = 8'h79 == _match_key_qbytes_2_T ? phv_data_121 : _GEN_5250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5252 = 8'h7a == _match_key_qbytes_2_T ? phv_data_122 : _GEN_5251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5253 = 8'h7b == _match_key_qbytes_2_T ? phv_data_123 : _GEN_5252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5254 = 8'h7c == _match_key_qbytes_2_T ? phv_data_124 : _GEN_5253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5255 = 8'h7d == _match_key_qbytes_2_T ? phv_data_125 : _GEN_5254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5256 = 8'h7e == _match_key_qbytes_2_T ? phv_data_126 : _GEN_5255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5257 = 8'h7f == _match_key_qbytes_2_T ? phv_data_127 : _GEN_5256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5258 = 8'h80 == _match_key_qbytes_2_T ? phv_data_128 : _GEN_5257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5259 = 8'h81 == _match_key_qbytes_2_T ? phv_data_129 : _GEN_5258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5260 = 8'h82 == _match_key_qbytes_2_T ? phv_data_130 : _GEN_5259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5261 = 8'h83 == _match_key_qbytes_2_T ? phv_data_131 : _GEN_5260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5262 = 8'h84 == _match_key_qbytes_2_T ? phv_data_132 : _GEN_5261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5263 = 8'h85 == _match_key_qbytes_2_T ? phv_data_133 : _GEN_5262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5264 = 8'h86 == _match_key_qbytes_2_T ? phv_data_134 : _GEN_5263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5265 = 8'h87 == _match_key_qbytes_2_T ? phv_data_135 : _GEN_5264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5266 = 8'h88 == _match_key_qbytes_2_T ? phv_data_136 : _GEN_5265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5267 = 8'h89 == _match_key_qbytes_2_T ? phv_data_137 : _GEN_5266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5268 = 8'h8a == _match_key_qbytes_2_T ? phv_data_138 : _GEN_5267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5269 = 8'h8b == _match_key_qbytes_2_T ? phv_data_139 : _GEN_5268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5270 = 8'h8c == _match_key_qbytes_2_T ? phv_data_140 : _GEN_5269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5271 = 8'h8d == _match_key_qbytes_2_T ? phv_data_141 : _GEN_5270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5272 = 8'h8e == _match_key_qbytes_2_T ? phv_data_142 : _GEN_5271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5273 = 8'h8f == _match_key_qbytes_2_T ? phv_data_143 : _GEN_5272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5274 = 8'h90 == _match_key_qbytes_2_T ? phv_data_144 : _GEN_5273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5275 = 8'h91 == _match_key_qbytes_2_T ? phv_data_145 : _GEN_5274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5276 = 8'h92 == _match_key_qbytes_2_T ? phv_data_146 : _GEN_5275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5277 = 8'h93 == _match_key_qbytes_2_T ? phv_data_147 : _GEN_5276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5278 = 8'h94 == _match_key_qbytes_2_T ? phv_data_148 : _GEN_5277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5279 = 8'h95 == _match_key_qbytes_2_T ? phv_data_149 : _GEN_5278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5280 = 8'h96 == _match_key_qbytes_2_T ? phv_data_150 : _GEN_5279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5281 = 8'h97 == _match_key_qbytes_2_T ? phv_data_151 : _GEN_5280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5282 = 8'h98 == _match_key_qbytes_2_T ? phv_data_152 : _GEN_5281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5283 = 8'h99 == _match_key_qbytes_2_T ? phv_data_153 : _GEN_5282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5284 = 8'h9a == _match_key_qbytes_2_T ? phv_data_154 : _GEN_5283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5285 = 8'h9b == _match_key_qbytes_2_T ? phv_data_155 : _GEN_5284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5286 = 8'h9c == _match_key_qbytes_2_T ? phv_data_156 : _GEN_5285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5287 = 8'h9d == _match_key_qbytes_2_T ? phv_data_157 : _GEN_5286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5288 = 8'h9e == _match_key_qbytes_2_T ? phv_data_158 : _GEN_5287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5289 = 8'h9f == _match_key_qbytes_2_T ? phv_data_159 : _GEN_5288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5290 = 8'ha0 == _match_key_qbytes_2_T ? phv_data_160 : _GEN_5289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5291 = 8'ha1 == _match_key_qbytes_2_T ? phv_data_161 : _GEN_5290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5292 = 8'ha2 == _match_key_qbytes_2_T ? phv_data_162 : _GEN_5291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5293 = 8'ha3 == _match_key_qbytes_2_T ? phv_data_163 : _GEN_5292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5294 = 8'ha4 == _match_key_qbytes_2_T ? phv_data_164 : _GEN_5293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5295 = 8'ha5 == _match_key_qbytes_2_T ? phv_data_165 : _GEN_5294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5296 = 8'ha6 == _match_key_qbytes_2_T ? phv_data_166 : _GEN_5295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5297 = 8'ha7 == _match_key_qbytes_2_T ? phv_data_167 : _GEN_5296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5298 = 8'ha8 == _match_key_qbytes_2_T ? phv_data_168 : _GEN_5297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5299 = 8'ha9 == _match_key_qbytes_2_T ? phv_data_169 : _GEN_5298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5300 = 8'haa == _match_key_qbytes_2_T ? phv_data_170 : _GEN_5299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5301 = 8'hab == _match_key_qbytes_2_T ? phv_data_171 : _GEN_5300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5302 = 8'hac == _match_key_qbytes_2_T ? phv_data_172 : _GEN_5301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5303 = 8'had == _match_key_qbytes_2_T ? phv_data_173 : _GEN_5302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5304 = 8'hae == _match_key_qbytes_2_T ? phv_data_174 : _GEN_5303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5305 = 8'haf == _match_key_qbytes_2_T ? phv_data_175 : _GEN_5304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5306 = 8'hb0 == _match_key_qbytes_2_T ? phv_data_176 : _GEN_5305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5307 = 8'hb1 == _match_key_qbytes_2_T ? phv_data_177 : _GEN_5306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5308 = 8'hb2 == _match_key_qbytes_2_T ? phv_data_178 : _GEN_5307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5309 = 8'hb3 == _match_key_qbytes_2_T ? phv_data_179 : _GEN_5308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5310 = 8'hb4 == _match_key_qbytes_2_T ? phv_data_180 : _GEN_5309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5311 = 8'hb5 == _match_key_qbytes_2_T ? phv_data_181 : _GEN_5310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5312 = 8'hb6 == _match_key_qbytes_2_T ? phv_data_182 : _GEN_5311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5313 = 8'hb7 == _match_key_qbytes_2_T ? phv_data_183 : _GEN_5312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5314 = 8'hb8 == _match_key_qbytes_2_T ? phv_data_184 : _GEN_5313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5315 = 8'hb9 == _match_key_qbytes_2_T ? phv_data_185 : _GEN_5314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5316 = 8'hba == _match_key_qbytes_2_T ? phv_data_186 : _GEN_5315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5317 = 8'hbb == _match_key_qbytes_2_T ? phv_data_187 : _GEN_5316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5318 = 8'hbc == _match_key_qbytes_2_T ? phv_data_188 : _GEN_5317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5319 = 8'hbd == _match_key_qbytes_2_T ? phv_data_189 : _GEN_5318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5320 = 8'hbe == _match_key_qbytes_2_T ? phv_data_190 : _GEN_5319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5321 = 8'hbf == _match_key_qbytes_2_T ? phv_data_191 : _GEN_5320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5322 = 8'hc0 == _match_key_qbytes_2_T ? phv_data_192 : _GEN_5321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5323 = 8'hc1 == _match_key_qbytes_2_T ? phv_data_193 : _GEN_5322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5324 = 8'hc2 == _match_key_qbytes_2_T ? phv_data_194 : _GEN_5323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5325 = 8'hc3 == _match_key_qbytes_2_T ? phv_data_195 : _GEN_5324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5326 = 8'hc4 == _match_key_qbytes_2_T ? phv_data_196 : _GEN_5325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5327 = 8'hc5 == _match_key_qbytes_2_T ? phv_data_197 : _GEN_5326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5328 = 8'hc6 == _match_key_qbytes_2_T ? phv_data_198 : _GEN_5327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5329 = 8'hc7 == _match_key_qbytes_2_T ? phv_data_199 : _GEN_5328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5330 = 8'hc8 == _match_key_qbytes_2_T ? phv_data_200 : _GEN_5329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5331 = 8'hc9 == _match_key_qbytes_2_T ? phv_data_201 : _GEN_5330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5332 = 8'hca == _match_key_qbytes_2_T ? phv_data_202 : _GEN_5331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5333 = 8'hcb == _match_key_qbytes_2_T ? phv_data_203 : _GEN_5332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5334 = 8'hcc == _match_key_qbytes_2_T ? phv_data_204 : _GEN_5333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5335 = 8'hcd == _match_key_qbytes_2_T ? phv_data_205 : _GEN_5334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5336 = 8'hce == _match_key_qbytes_2_T ? phv_data_206 : _GEN_5335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5337 = 8'hcf == _match_key_qbytes_2_T ? phv_data_207 : _GEN_5336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5338 = 8'hd0 == _match_key_qbytes_2_T ? phv_data_208 : _GEN_5337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5339 = 8'hd1 == _match_key_qbytes_2_T ? phv_data_209 : _GEN_5338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5340 = 8'hd2 == _match_key_qbytes_2_T ? phv_data_210 : _GEN_5339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5341 = 8'hd3 == _match_key_qbytes_2_T ? phv_data_211 : _GEN_5340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5342 = 8'hd4 == _match_key_qbytes_2_T ? phv_data_212 : _GEN_5341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5343 = 8'hd5 == _match_key_qbytes_2_T ? phv_data_213 : _GEN_5342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5344 = 8'hd6 == _match_key_qbytes_2_T ? phv_data_214 : _GEN_5343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5345 = 8'hd7 == _match_key_qbytes_2_T ? phv_data_215 : _GEN_5344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5346 = 8'hd8 == _match_key_qbytes_2_T ? phv_data_216 : _GEN_5345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5347 = 8'hd9 == _match_key_qbytes_2_T ? phv_data_217 : _GEN_5346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5348 = 8'hda == _match_key_qbytes_2_T ? phv_data_218 : _GEN_5347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5349 = 8'hdb == _match_key_qbytes_2_T ? phv_data_219 : _GEN_5348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5350 = 8'hdc == _match_key_qbytes_2_T ? phv_data_220 : _GEN_5349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5351 = 8'hdd == _match_key_qbytes_2_T ? phv_data_221 : _GEN_5350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5352 = 8'hde == _match_key_qbytes_2_T ? phv_data_222 : _GEN_5351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5353 = 8'hdf == _match_key_qbytes_2_T ? phv_data_223 : _GEN_5352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5354 = 8'he0 == _match_key_qbytes_2_T ? phv_data_224 : _GEN_5353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5355 = 8'he1 == _match_key_qbytes_2_T ? phv_data_225 : _GEN_5354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5356 = 8'he2 == _match_key_qbytes_2_T ? phv_data_226 : _GEN_5355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5357 = 8'he3 == _match_key_qbytes_2_T ? phv_data_227 : _GEN_5356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5358 = 8'he4 == _match_key_qbytes_2_T ? phv_data_228 : _GEN_5357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5359 = 8'he5 == _match_key_qbytes_2_T ? phv_data_229 : _GEN_5358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5360 = 8'he6 == _match_key_qbytes_2_T ? phv_data_230 : _GEN_5359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5361 = 8'he7 == _match_key_qbytes_2_T ? phv_data_231 : _GEN_5360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5362 = 8'he8 == _match_key_qbytes_2_T ? phv_data_232 : _GEN_5361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5363 = 8'he9 == _match_key_qbytes_2_T ? phv_data_233 : _GEN_5362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5364 = 8'hea == _match_key_qbytes_2_T ? phv_data_234 : _GEN_5363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5365 = 8'heb == _match_key_qbytes_2_T ? phv_data_235 : _GEN_5364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5366 = 8'hec == _match_key_qbytes_2_T ? phv_data_236 : _GEN_5365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5367 = 8'hed == _match_key_qbytes_2_T ? phv_data_237 : _GEN_5366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5368 = 8'hee == _match_key_qbytes_2_T ? phv_data_238 : _GEN_5367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5369 = 8'hef == _match_key_qbytes_2_T ? phv_data_239 : _GEN_5368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5370 = 8'hf0 == _match_key_qbytes_2_T ? phv_data_240 : _GEN_5369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5371 = 8'hf1 == _match_key_qbytes_2_T ? phv_data_241 : _GEN_5370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5372 = 8'hf2 == _match_key_qbytes_2_T ? phv_data_242 : _GEN_5371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5373 = 8'hf3 == _match_key_qbytes_2_T ? phv_data_243 : _GEN_5372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5374 = 8'hf4 == _match_key_qbytes_2_T ? phv_data_244 : _GEN_5373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5375 = 8'hf5 == _match_key_qbytes_2_T ? phv_data_245 : _GEN_5374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5376 = 8'hf6 == _match_key_qbytes_2_T ? phv_data_246 : _GEN_5375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5377 = 8'hf7 == _match_key_qbytes_2_T ? phv_data_247 : _GEN_5376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5378 = 8'hf8 == _match_key_qbytes_2_T ? phv_data_248 : _GEN_5377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5379 = 8'hf9 == _match_key_qbytes_2_T ? phv_data_249 : _GEN_5378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5380 = 8'hfa == _match_key_qbytes_2_T ? phv_data_250 : _GEN_5379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5381 = 8'hfb == _match_key_qbytes_2_T ? phv_data_251 : _GEN_5380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5382 = 8'hfc == _match_key_qbytes_2_T ? phv_data_252 : _GEN_5381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5383 = 8'hfd == _match_key_qbytes_2_T ? phv_data_253 : _GEN_5382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5384 = 8'hfe == _match_key_qbytes_2_T ? phv_data_254 : _GEN_5383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5385 = 8'hff == _match_key_qbytes_2_T ? phv_data_255 : _GEN_5384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_14886 = {{1'd0}, _match_key_qbytes_2_T}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5386 = 9'h100 == _GEN_14886 ? phv_data_256 : _GEN_5385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5387 = 9'h101 == _GEN_14886 ? phv_data_257 : _GEN_5386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5388 = 9'h102 == _GEN_14886 ? phv_data_258 : _GEN_5387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5389 = 9'h103 == _GEN_14886 ? phv_data_259 : _GEN_5388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5390 = 9'h104 == _GEN_14886 ? phv_data_260 : _GEN_5389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5391 = 9'h105 == _GEN_14886 ? phv_data_261 : _GEN_5390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5392 = 9'h106 == _GEN_14886 ? phv_data_262 : _GEN_5391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5393 = 9'h107 == _GEN_14886 ? phv_data_263 : _GEN_5392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5394 = 9'h108 == _GEN_14886 ? phv_data_264 : _GEN_5393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5395 = 9'h109 == _GEN_14886 ? phv_data_265 : _GEN_5394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5396 = 9'h10a == _GEN_14886 ? phv_data_266 : _GEN_5395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5397 = 9'h10b == _GEN_14886 ? phv_data_267 : _GEN_5396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5398 = 9'h10c == _GEN_14886 ? phv_data_268 : _GEN_5397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5399 = 9'h10d == _GEN_14886 ? phv_data_269 : _GEN_5398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5400 = 9'h10e == _GEN_14886 ? phv_data_270 : _GEN_5399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5401 = 9'h10f == _GEN_14886 ? phv_data_271 : _GEN_5400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5402 = 9'h110 == _GEN_14886 ? phv_data_272 : _GEN_5401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5403 = 9'h111 == _GEN_14886 ? phv_data_273 : _GEN_5402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5404 = 9'h112 == _GEN_14886 ? phv_data_274 : _GEN_5403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5405 = 9'h113 == _GEN_14886 ? phv_data_275 : _GEN_5404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5406 = 9'h114 == _GEN_14886 ? phv_data_276 : _GEN_5405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5407 = 9'h115 == _GEN_14886 ? phv_data_277 : _GEN_5406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5408 = 9'h116 == _GEN_14886 ? phv_data_278 : _GEN_5407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5409 = 9'h117 == _GEN_14886 ? phv_data_279 : _GEN_5408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5410 = 9'h118 == _GEN_14886 ? phv_data_280 : _GEN_5409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5411 = 9'h119 == _GEN_14886 ? phv_data_281 : _GEN_5410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5412 = 9'h11a == _GEN_14886 ? phv_data_282 : _GEN_5411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5413 = 9'h11b == _GEN_14886 ? phv_data_283 : _GEN_5412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5414 = 9'h11c == _GEN_14886 ? phv_data_284 : _GEN_5413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5415 = 9'h11d == _GEN_14886 ? phv_data_285 : _GEN_5414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5416 = 9'h11e == _GEN_14886 ? phv_data_286 : _GEN_5415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5417 = 9'h11f == _GEN_14886 ? phv_data_287 : _GEN_5416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5418 = 9'h120 == _GEN_14886 ? phv_data_288 : _GEN_5417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5419 = 9'h121 == _GEN_14886 ? phv_data_289 : _GEN_5418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5420 = 9'h122 == _GEN_14886 ? phv_data_290 : _GEN_5419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5421 = 9'h123 == _GEN_14886 ? phv_data_291 : _GEN_5420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5422 = 9'h124 == _GEN_14886 ? phv_data_292 : _GEN_5421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5423 = 9'h125 == _GEN_14886 ? phv_data_293 : _GEN_5422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5424 = 9'h126 == _GEN_14886 ? phv_data_294 : _GEN_5423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5425 = 9'h127 == _GEN_14886 ? phv_data_295 : _GEN_5424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5426 = 9'h128 == _GEN_14886 ? phv_data_296 : _GEN_5425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5427 = 9'h129 == _GEN_14886 ? phv_data_297 : _GEN_5426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5428 = 9'h12a == _GEN_14886 ? phv_data_298 : _GEN_5427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5429 = 9'h12b == _GEN_14886 ? phv_data_299 : _GEN_5428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5430 = 9'h12c == _GEN_14886 ? phv_data_300 : _GEN_5429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5431 = 9'h12d == _GEN_14886 ? phv_data_301 : _GEN_5430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5432 = 9'h12e == _GEN_14886 ? phv_data_302 : _GEN_5431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5433 = 9'h12f == _GEN_14886 ? phv_data_303 : _GEN_5432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5434 = 9'h130 == _GEN_14886 ? phv_data_304 : _GEN_5433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5435 = 9'h131 == _GEN_14886 ? phv_data_305 : _GEN_5434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5436 = 9'h132 == _GEN_14886 ? phv_data_306 : _GEN_5435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5437 = 9'h133 == _GEN_14886 ? phv_data_307 : _GEN_5436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5438 = 9'h134 == _GEN_14886 ? phv_data_308 : _GEN_5437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5439 = 9'h135 == _GEN_14886 ? phv_data_309 : _GEN_5438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5440 = 9'h136 == _GEN_14886 ? phv_data_310 : _GEN_5439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5441 = 9'h137 == _GEN_14886 ? phv_data_311 : _GEN_5440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5442 = 9'h138 == _GEN_14886 ? phv_data_312 : _GEN_5441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5443 = 9'h139 == _GEN_14886 ? phv_data_313 : _GEN_5442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5444 = 9'h13a == _GEN_14886 ? phv_data_314 : _GEN_5443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5445 = 9'h13b == _GEN_14886 ? phv_data_315 : _GEN_5444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5446 = 9'h13c == _GEN_14886 ? phv_data_316 : _GEN_5445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5447 = 9'h13d == _GEN_14886 ? phv_data_317 : _GEN_5446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5448 = 9'h13e == _GEN_14886 ? phv_data_318 : _GEN_5447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5449 = 9'h13f == _GEN_14886 ? phv_data_319 : _GEN_5448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5450 = 9'h140 == _GEN_14886 ? phv_data_320 : _GEN_5449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5451 = 9'h141 == _GEN_14886 ? phv_data_321 : _GEN_5450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5452 = 9'h142 == _GEN_14886 ? phv_data_322 : _GEN_5451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5453 = 9'h143 == _GEN_14886 ? phv_data_323 : _GEN_5452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5454 = 9'h144 == _GEN_14886 ? phv_data_324 : _GEN_5453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5455 = 9'h145 == _GEN_14886 ? phv_data_325 : _GEN_5454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5456 = 9'h146 == _GEN_14886 ? phv_data_326 : _GEN_5455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5457 = 9'h147 == _GEN_14886 ? phv_data_327 : _GEN_5456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5458 = 9'h148 == _GEN_14886 ? phv_data_328 : _GEN_5457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5459 = 9'h149 == _GEN_14886 ? phv_data_329 : _GEN_5458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5460 = 9'h14a == _GEN_14886 ? phv_data_330 : _GEN_5459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5461 = 9'h14b == _GEN_14886 ? phv_data_331 : _GEN_5460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5462 = 9'h14c == _GEN_14886 ? phv_data_332 : _GEN_5461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5463 = 9'h14d == _GEN_14886 ? phv_data_333 : _GEN_5462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5464 = 9'h14e == _GEN_14886 ? phv_data_334 : _GEN_5463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5465 = 9'h14f == _GEN_14886 ? phv_data_335 : _GEN_5464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5466 = 9'h150 == _GEN_14886 ? phv_data_336 : _GEN_5465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5467 = 9'h151 == _GEN_14886 ? phv_data_337 : _GEN_5466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5468 = 9'h152 == _GEN_14886 ? phv_data_338 : _GEN_5467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5469 = 9'h153 == _GEN_14886 ? phv_data_339 : _GEN_5468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5470 = 9'h154 == _GEN_14886 ? phv_data_340 : _GEN_5469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5471 = 9'h155 == _GEN_14886 ? phv_data_341 : _GEN_5470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5472 = 9'h156 == _GEN_14886 ? phv_data_342 : _GEN_5471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5473 = 9'h157 == _GEN_14886 ? phv_data_343 : _GEN_5472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5474 = 9'h158 == _GEN_14886 ? phv_data_344 : _GEN_5473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5475 = 9'h159 == _GEN_14886 ? phv_data_345 : _GEN_5474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5476 = 9'h15a == _GEN_14886 ? phv_data_346 : _GEN_5475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5477 = 9'h15b == _GEN_14886 ? phv_data_347 : _GEN_5476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5478 = 9'h15c == _GEN_14886 ? phv_data_348 : _GEN_5477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5479 = 9'h15d == _GEN_14886 ? phv_data_349 : _GEN_5478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5480 = 9'h15e == _GEN_14886 ? phv_data_350 : _GEN_5479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5481 = 9'h15f == _GEN_14886 ? phv_data_351 : _GEN_5480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5482 = 9'h160 == _GEN_14886 ? phv_data_352 : _GEN_5481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5483 = 9'h161 == _GEN_14886 ? phv_data_353 : _GEN_5482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5484 = 9'h162 == _GEN_14886 ? phv_data_354 : _GEN_5483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5485 = 9'h163 == _GEN_14886 ? phv_data_355 : _GEN_5484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5486 = 9'h164 == _GEN_14886 ? phv_data_356 : _GEN_5485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5487 = 9'h165 == _GEN_14886 ? phv_data_357 : _GEN_5486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5488 = 9'h166 == _GEN_14886 ? phv_data_358 : _GEN_5487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5489 = 9'h167 == _GEN_14886 ? phv_data_359 : _GEN_5488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5490 = 9'h168 == _GEN_14886 ? phv_data_360 : _GEN_5489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5491 = 9'h169 == _GEN_14886 ? phv_data_361 : _GEN_5490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5492 = 9'h16a == _GEN_14886 ? phv_data_362 : _GEN_5491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5493 = 9'h16b == _GEN_14886 ? phv_data_363 : _GEN_5492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5494 = 9'h16c == _GEN_14886 ? phv_data_364 : _GEN_5493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5495 = 9'h16d == _GEN_14886 ? phv_data_365 : _GEN_5494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5496 = 9'h16e == _GEN_14886 ? phv_data_366 : _GEN_5495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5497 = 9'h16f == _GEN_14886 ? phv_data_367 : _GEN_5496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5498 = 9'h170 == _GEN_14886 ? phv_data_368 : _GEN_5497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5499 = 9'h171 == _GEN_14886 ? phv_data_369 : _GEN_5498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5500 = 9'h172 == _GEN_14886 ? phv_data_370 : _GEN_5499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5501 = 9'h173 == _GEN_14886 ? phv_data_371 : _GEN_5500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5502 = 9'h174 == _GEN_14886 ? phv_data_372 : _GEN_5501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5503 = 9'h175 == _GEN_14886 ? phv_data_373 : _GEN_5502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5504 = 9'h176 == _GEN_14886 ? phv_data_374 : _GEN_5503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5505 = 9'h177 == _GEN_14886 ? phv_data_375 : _GEN_5504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5506 = 9'h178 == _GEN_14886 ? phv_data_376 : _GEN_5505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5507 = 9'h179 == _GEN_14886 ? phv_data_377 : _GEN_5506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5508 = 9'h17a == _GEN_14886 ? phv_data_378 : _GEN_5507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5509 = 9'h17b == _GEN_14886 ? phv_data_379 : _GEN_5508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5510 = 9'h17c == _GEN_14886 ? phv_data_380 : _GEN_5509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5511 = 9'h17d == _GEN_14886 ? phv_data_381 : _GEN_5510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5512 = 9'h17e == _GEN_14886 ? phv_data_382 : _GEN_5511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5513 = 9'h17f == _GEN_14886 ? phv_data_383 : _GEN_5512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5514 = 9'h180 == _GEN_14886 ? phv_data_384 : _GEN_5513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5515 = 9'h181 == _GEN_14886 ? phv_data_385 : _GEN_5514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5516 = 9'h182 == _GEN_14886 ? phv_data_386 : _GEN_5515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5517 = 9'h183 == _GEN_14886 ? phv_data_387 : _GEN_5516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5518 = 9'h184 == _GEN_14886 ? phv_data_388 : _GEN_5517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5519 = 9'h185 == _GEN_14886 ? phv_data_389 : _GEN_5518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5520 = 9'h186 == _GEN_14886 ? phv_data_390 : _GEN_5519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5521 = 9'h187 == _GEN_14886 ? phv_data_391 : _GEN_5520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5522 = 9'h188 == _GEN_14886 ? phv_data_392 : _GEN_5521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5523 = 9'h189 == _GEN_14886 ? phv_data_393 : _GEN_5522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5524 = 9'h18a == _GEN_14886 ? phv_data_394 : _GEN_5523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5525 = 9'h18b == _GEN_14886 ? phv_data_395 : _GEN_5524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5526 = 9'h18c == _GEN_14886 ? phv_data_396 : _GEN_5525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5527 = 9'h18d == _GEN_14886 ? phv_data_397 : _GEN_5526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5528 = 9'h18e == _GEN_14886 ? phv_data_398 : _GEN_5527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5529 = 9'h18f == _GEN_14886 ? phv_data_399 : _GEN_5528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5530 = 9'h190 == _GEN_14886 ? phv_data_400 : _GEN_5529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5531 = 9'h191 == _GEN_14886 ? phv_data_401 : _GEN_5530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5532 = 9'h192 == _GEN_14886 ? phv_data_402 : _GEN_5531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5533 = 9'h193 == _GEN_14886 ? phv_data_403 : _GEN_5532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5534 = 9'h194 == _GEN_14886 ? phv_data_404 : _GEN_5533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5535 = 9'h195 == _GEN_14886 ? phv_data_405 : _GEN_5534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5536 = 9'h196 == _GEN_14886 ? phv_data_406 : _GEN_5535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5537 = 9'h197 == _GEN_14886 ? phv_data_407 : _GEN_5536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5538 = 9'h198 == _GEN_14886 ? phv_data_408 : _GEN_5537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5539 = 9'h199 == _GEN_14886 ? phv_data_409 : _GEN_5538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5540 = 9'h19a == _GEN_14886 ? phv_data_410 : _GEN_5539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5541 = 9'h19b == _GEN_14886 ? phv_data_411 : _GEN_5540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5542 = 9'h19c == _GEN_14886 ? phv_data_412 : _GEN_5541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5543 = 9'h19d == _GEN_14886 ? phv_data_413 : _GEN_5542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5544 = 9'h19e == _GEN_14886 ? phv_data_414 : _GEN_5543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5545 = 9'h19f == _GEN_14886 ? phv_data_415 : _GEN_5544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5546 = 9'h1a0 == _GEN_14886 ? phv_data_416 : _GEN_5545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5547 = 9'h1a1 == _GEN_14886 ? phv_data_417 : _GEN_5546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5548 = 9'h1a2 == _GEN_14886 ? phv_data_418 : _GEN_5547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5549 = 9'h1a3 == _GEN_14886 ? phv_data_419 : _GEN_5548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5550 = 9'h1a4 == _GEN_14886 ? phv_data_420 : _GEN_5549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5551 = 9'h1a5 == _GEN_14886 ? phv_data_421 : _GEN_5550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5552 = 9'h1a6 == _GEN_14886 ? phv_data_422 : _GEN_5551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5553 = 9'h1a7 == _GEN_14886 ? phv_data_423 : _GEN_5552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5554 = 9'h1a8 == _GEN_14886 ? phv_data_424 : _GEN_5553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5555 = 9'h1a9 == _GEN_14886 ? phv_data_425 : _GEN_5554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5556 = 9'h1aa == _GEN_14886 ? phv_data_426 : _GEN_5555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5557 = 9'h1ab == _GEN_14886 ? phv_data_427 : _GEN_5556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5558 = 9'h1ac == _GEN_14886 ? phv_data_428 : _GEN_5557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5559 = 9'h1ad == _GEN_14886 ? phv_data_429 : _GEN_5558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5560 = 9'h1ae == _GEN_14886 ? phv_data_430 : _GEN_5559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5561 = 9'h1af == _GEN_14886 ? phv_data_431 : _GEN_5560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5562 = 9'h1b0 == _GEN_14886 ? phv_data_432 : _GEN_5561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5563 = 9'h1b1 == _GEN_14886 ? phv_data_433 : _GEN_5562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5564 = 9'h1b2 == _GEN_14886 ? phv_data_434 : _GEN_5563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5565 = 9'h1b3 == _GEN_14886 ? phv_data_435 : _GEN_5564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5566 = 9'h1b4 == _GEN_14886 ? phv_data_436 : _GEN_5565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5567 = 9'h1b5 == _GEN_14886 ? phv_data_437 : _GEN_5566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5568 = 9'h1b6 == _GEN_14886 ? phv_data_438 : _GEN_5567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5569 = 9'h1b7 == _GEN_14886 ? phv_data_439 : _GEN_5568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5570 = 9'h1b8 == _GEN_14886 ? phv_data_440 : _GEN_5569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5571 = 9'h1b9 == _GEN_14886 ? phv_data_441 : _GEN_5570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5572 = 9'h1ba == _GEN_14886 ? phv_data_442 : _GEN_5571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5573 = 9'h1bb == _GEN_14886 ? phv_data_443 : _GEN_5572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5574 = 9'h1bc == _GEN_14886 ? phv_data_444 : _GEN_5573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5575 = 9'h1bd == _GEN_14886 ? phv_data_445 : _GEN_5574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5576 = 9'h1be == _GEN_14886 ? phv_data_446 : _GEN_5575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5577 = 9'h1bf == _GEN_14886 ? phv_data_447 : _GEN_5576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5578 = 9'h1c0 == _GEN_14886 ? phv_data_448 : _GEN_5577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5579 = 9'h1c1 == _GEN_14886 ? phv_data_449 : _GEN_5578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5580 = 9'h1c2 == _GEN_14886 ? phv_data_450 : _GEN_5579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5581 = 9'h1c3 == _GEN_14886 ? phv_data_451 : _GEN_5580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5582 = 9'h1c4 == _GEN_14886 ? phv_data_452 : _GEN_5581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5583 = 9'h1c5 == _GEN_14886 ? phv_data_453 : _GEN_5582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5584 = 9'h1c6 == _GEN_14886 ? phv_data_454 : _GEN_5583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5585 = 9'h1c7 == _GEN_14886 ? phv_data_455 : _GEN_5584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5586 = 9'h1c8 == _GEN_14886 ? phv_data_456 : _GEN_5585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5587 = 9'h1c9 == _GEN_14886 ? phv_data_457 : _GEN_5586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5588 = 9'h1ca == _GEN_14886 ? phv_data_458 : _GEN_5587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5589 = 9'h1cb == _GEN_14886 ? phv_data_459 : _GEN_5588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5590 = 9'h1cc == _GEN_14886 ? phv_data_460 : _GEN_5589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5591 = 9'h1cd == _GEN_14886 ? phv_data_461 : _GEN_5590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5592 = 9'h1ce == _GEN_14886 ? phv_data_462 : _GEN_5591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5593 = 9'h1cf == _GEN_14886 ? phv_data_463 : _GEN_5592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5594 = 9'h1d0 == _GEN_14886 ? phv_data_464 : _GEN_5593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5595 = 9'h1d1 == _GEN_14886 ? phv_data_465 : _GEN_5594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5596 = 9'h1d2 == _GEN_14886 ? phv_data_466 : _GEN_5595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5597 = 9'h1d3 == _GEN_14886 ? phv_data_467 : _GEN_5596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5598 = 9'h1d4 == _GEN_14886 ? phv_data_468 : _GEN_5597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5599 = 9'h1d5 == _GEN_14886 ? phv_data_469 : _GEN_5598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5600 = 9'h1d6 == _GEN_14886 ? phv_data_470 : _GEN_5599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5601 = 9'h1d7 == _GEN_14886 ? phv_data_471 : _GEN_5600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5602 = 9'h1d8 == _GEN_14886 ? phv_data_472 : _GEN_5601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5603 = 9'h1d9 == _GEN_14886 ? phv_data_473 : _GEN_5602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5604 = 9'h1da == _GEN_14886 ? phv_data_474 : _GEN_5603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5605 = 9'h1db == _GEN_14886 ? phv_data_475 : _GEN_5604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5606 = 9'h1dc == _GEN_14886 ? phv_data_476 : _GEN_5605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5607 = 9'h1dd == _GEN_14886 ? phv_data_477 : _GEN_5606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5608 = 9'h1de == _GEN_14886 ? phv_data_478 : _GEN_5607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5609 = 9'h1df == _GEN_14886 ? phv_data_479 : _GEN_5608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5610 = 9'h1e0 == _GEN_14886 ? phv_data_480 : _GEN_5609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5611 = 9'h1e1 == _GEN_14886 ? phv_data_481 : _GEN_5610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5612 = 9'h1e2 == _GEN_14886 ? phv_data_482 : _GEN_5611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5613 = 9'h1e3 == _GEN_14886 ? phv_data_483 : _GEN_5612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5614 = 9'h1e4 == _GEN_14886 ? phv_data_484 : _GEN_5613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5615 = 9'h1e5 == _GEN_14886 ? phv_data_485 : _GEN_5614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5616 = 9'h1e6 == _GEN_14886 ? phv_data_486 : _GEN_5615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5617 = 9'h1e7 == _GEN_14886 ? phv_data_487 : _GEN_5616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5618 = 9'h1e8 == _GEN_14886 ? phv_data_488 : _GEN_5617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5619 = 9'h1e9 == _GEN_14886 ? phv_data_489 : _GEN_5618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5620 = 9'h1ea == _GEN_14886 ? phv_data_490 : _GEN_5619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5621 = 9'h1eb == _GEN_14886 ? phv_data_491 : _GEN_5620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5622 = 9'h1ec == _GEN_14886 ? phv_data_492 : _GEN_5621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5623 = 9'h1ed == _GEN_14886 ? phv_data_493 : _GEN_5622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5624 = 9'h1ee == _GEN_14886 ? phv_data_494 : _GEN_5623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5625 = 9'h1ef == _GEN_14886 ? phv_data_495 : _GEN_5624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5626 = 9'h1f0 == _GEN_14886 ? phv_data_496 : _GEN_5625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5627 = 9'h1f1 == _GEN_14886 ? phv_data_497 : _GEN_5626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5628 = 9'h1f2 == _GEN_14886 ? phv_data_498 : _GEN_5627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5629 = 9'h1f3 == _GEN_14886 ? phv_data_499 : _GEN_5628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5630 = 9'h1f4 == _GEN_14886 ? phv_data_500 : _GEN_5629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5631 = 9'h1f5 == _GEN_14886 ? phv_data_501 : _GEN_5630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5632 = 9'h1f6 == _GEN_14886 ? phv_data_502 : _GEN_5631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5633 = 9'h1f7 == _GEN_14886 ? phv_data_503 : _GEN_5632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5634 = 9'h1f8 == _GEN_14886 ? phv_data_504 : _GEN_5633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5635 = 9'h1f9 == _GEN_14886 ? phv_data_505 : _GEN_5634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5636 = 9'h1fa == _GEN_14886 ? phv_data_506 : _GEN_5635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5637 = 9'h1fb == _GEN_14886 ? phv_data_507 : _GEN_5636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5638 = 9'h1fc == _GEN_14886 ? phv_data_508 : _GEN_5637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5639 = 9'h1fd == _GEN_14886 ? phv_data_509 : _GEN_5638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5640 = 9'h1fe == _GEN_14886 ? phv_data_510 : _GEN_5639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5641 = 9'h1ff == _GEN_14886 ? phv_data_511 : _GEN_5640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5643 = 8'h1 == _match_key_qbytes_2_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5644 = 8'h2 == _match_key_qbytes_2_T_1 ? phv_data_2 : _GEN_5643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5645 = 8'h3 == _match_key_qbytes_2_T_1 ? phv_data_3 : _GEN_5644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5646 = 8'h4 == _match_key_qbytes_2_T_1 ? phv_data_4 : _GEN_5645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5647 = 8'h5 == _match_key_qbytes_2_T_1 ? phv_data_5 : _GEN_5646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5648 = 8'h6 == _match_key_qbytes_2_T_1 ? phv_data_6 : _GEN_5647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5649 = 8'h7 == _match_key_qbytes_2_T_1 ? phv_data_7 : _GEN_5648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5650 = 8'h8 == _match_key_qbytes_2_T_1 ? phv_data_8 : _GEN_5649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5651 = 8'h9 == _match_key_qbytes_2_T_1 ? phv_data_9 : _GEN_5650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5652 = 8'ha == _match_key_qbytes_2_T_1 ? phv_data_10 : _GEN_5651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5653 = 8'hb == _match_key_qbytes_2_T_1 ? phv_data_11 : _GEN_5652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5654 = 8'hc == _match_key_qbytes_2_T_1 ? phv_data_12 : _GEN_5653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5655 = 8'hd == _match_key_qbytes_2_T_1 ? phv_data_13 : _GEN_5654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5656 = 8'he == _match_key_qbytes_2_T_1 ? phv_data_14 : _GEN_5655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5657 = 8'hf == _match_key_qbytes_2_T_1 ? phv_data_15 : _GEN_5656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5658 = 8'h10 == _match_key_qbytes_2_T_1 ? phv_data_16 : _GEN_5657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5659 = 8'h11 == _match_key_qbytes_2_T_1 ? phv_data_17 : _GEN_5658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5660 = 8'h12 == _match_key_qbytes_2_T_1 ? phv_data_18 : _GEN_5659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5661 = 8'h13 == _match_key_qbytes_2_T_1 ? phv_data_19 : _GEN_5660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5662 = 8'h14 == _match_key_qbytes_2_T_1 ? phv_data_20 : _GEN_5661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5663 = 8'h15 == _match_key_qbytes_2_T_1 ? phv_data_21 : _GEN_5662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5664 = 8'h16 == _match_key_qbytes_2_T_1 ? phv_data_22 : _GEN_5663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5665 = 8'h17 == _match_key_qbytes_2_T_1 ? phv_data_23 : _GEN_5664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5666 = 8'h18 == _match_key_qbytes_2_T_1 ? phv_data_24 : _GEN_5665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5667 = 8'h19 == _match_key_qbytes_2_T_1 ? phv_data_25 : _GEN_5666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5668 = 8'h1a == _match_key_qbytes_2_T_1 ? phv_data_26 : _GEN_5667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5669 = 8'h1b == _match_key_qbytes_2_T_1 ? phv_data_27 : _GEN_5668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5670 = 8'h1c == _match_key_qbytes_2_T_1 ? phv_data_28 : _GEN_5669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5671 = 8'h1d == _match_key_qbytes_2_T_1 ? phv_data_29 : _GEN_5670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5672 = 8'h1e == _match_key_qbytes_2_T_1 ? phv_data_30 : _GEN_5671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5673 = 8'h1f == _match_key_qbytes_2_T_1 ? phv_data_31 : _GEN_5672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5674 = 8'h20 == _match_key_qbytes_2_T_1 ? phv_data_32 : _GEN_5673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5675 = 8'h21 == _match_key_qbytes_2_T_1 ? phv_data_33 : _GEN_5674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5676 = 8'h22 == _match_key_qbytes_2_T_1 ? phv_data_34 : _GEN_5675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5677 = 8'h23 == _match_key_qbytes_2_T_1 ? phv_data_35 : _GEN_5676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5678 = 8'h24 == _match_key_qbytes_2_T_1 ? phv_data_36 : _GEN_5677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5679 = 8'h25 == _match_key_qbytes_2_T_1 ? phv_data_37 : _GEN_5678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5680 = 8'h26 == _match_key_qbytes_2_T_1 ? phv_data_38 : _GEN_5679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5681 = 8'h27 == _match_key_qbytes_2_T_1 ? phv_data_39 : _GEN_5680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5682 = 8'h28 == _match_key_qbytes_2_T_1 ? phv_data_40 : _GEN_5681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5683 = 8'h29 == _match_key_qbytes_2_T_1 ? phv_data_41 : _GEN_5682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5684 = 8'h2a == _match_key_qbytes_2_T_1 ? phv_data_42 : _GEN_5683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5685 = 8'h2b == _match_key_qbytes_2_T_1 ? phv_data_43 : _GEN_5684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5686 = 8'h2c == _match_key_qbytes_2_T_1 ? phv_data_44 : _GEN_5685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5687 = 8'h2d == _match_key_qbytes_2_T_1 ? phv_data_45 : _GEN_5686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5688 = 8'h2e == _match_key_qbytes_2_T_1 ? phv_data_46 : _GEN_5687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5689 = 8'h2f == _match_key_qbytes_2_T_1 ? phv_data_47 : _GEN_5688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5690 = 8'h30 == _match_key_qbytes_2_T_1 ? phv_data_48 : _GEN_5689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5691 = 8'h31 == _match_key_qbytes_2_T_1 ? phv_data_49 : _GEN_5690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5692 = 8'h32 == _match_key_qbytes_2_T_1 ? phv_data_50 : _GEN_5691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5693 = 8'h33 == _match_key_qbytes_2_T_1 ? phv_data_51 : _GEN_5692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5694 = 8'h34 == _match_key_qbytes_2_T_1 ? phv_data_52 : _GEN_5693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5695 = 8'h35 == _match_key_qbytes_2_T_1 ? phv_data_53 : _GEN_5694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5696 = 8'h36 == _match_key_qbytes_2_T_1 ? phv_data_54 : _GEN_5695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5697 = 8'h37 == _match_key_qbytes_2_T_1 ? phv_data_55 : _GEN_5696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5698 = 8'h38 == _match_key_qbytes_2_T_1 ? phv_data_56 : _GEN_5697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5699 = 8'h39 == _match_key_qbytes_2_T_1 ? phv_data_57 : _GEN_5698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5700 = 8'h3a == _match_key_qbytes_2_T_1 ? phv_data_58 : _GEN_5699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5701 = 8'h3b == _match_key_qbytes_2_T_1 ? phv_data_59 : _GEN_5700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5702 = 8'h3c == _match_key_qbytes_2_T_1 ? phv_data_60 : _GEN_5701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5703 = 8'h3d == _match_key_qbytes_2_T_1 ? phv_data_61 : _GEN_5702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5704 = 8'h3e == _match_key_qbytes_2_T_1 ? phv_data_62 : _GEN_5703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5705 = 8'h3f == _match_key_qbytes_2_T_1 ? phv_data_63 : _GEN_5704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5706 = 8'h40 == _match_key_qbytes_2_T_1 ? phv_data_64 : _GEN_5705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5707 = 8'h41 == _match_key_qbytes_2_T_1 ? phv_data_65 : _GEN_5706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5708 = 8'h42 == _match_key_qbytes_2_T_1 ? phv_data_66 : _GEN_5707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5709 = 8'h43 == _match_key_qbytes_2_T_1 ? phv_data_67 : _GEN_5708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5710 = 8'h44 == _match_key_qbytes_2_T_1 ? phv_data_68 : _GEN_5709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5711 = 8'h45 == _match_key_qbytes_2_T_1 ? phv_data_69 : _GEN_5710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5712 = 8'h46 == _match_key_qbytes_2_T_1 ? phv_data_70 : _GEN_5711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5713 = 8'h47 == _match_key_qbytes_2_T_1 ? phv_data_71 : _GEN_5712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5714 = 8'h48 == _match_key_qbytes_2_T_1 ? phv_data_72 : _GEN_5713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5715 = 8'h49 == _match_key_qbytes_2_T_1 ? phv_data_73 : _GEN_5714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5716 = 8'h4a == _match_key_qbytes_2_T_1 ? phv_data_74 : _GEN_5715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5717 = 8'h4b == _match_key_qbytes_2_T_1 ? phv_data_75 : _GEN_5716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5718 = 8'h4c == _match_key_qbytes_2_T_1 ? phv_data_76 : _GEN_5717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5719 = 8'h4d == _match_key_qbytes_2_T_1 ? phv_data_77 : _GEN_5718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5720 = 8'h4e == _match_key_qbytes_2_T_1 ? phv_data_78 : _GEN_5719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5721 = 8'h4f == _match_key_qbytes_2_T_1 ? phv_data_79 : _GEN_5720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5722 = 8'h50 == _match_key_qbytes_2_T_1 ? phv_data_80 : _GEN_5721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5723 = 8'h51 == _match_key_qbytes_2_T_1 ? phv_data_81 : _GEN_5722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5724 = 8'h52 == _match_key_qbytes_2_T_1 ? phv_data_82 : _GEN_5723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5725 = 8'h53 == _match_key_qbytes_2_T_1 ? phv_data_83 : _GEN_5724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5726 = 8'h54 == _match_key_qbytes_2_T_1 ? phv_data_84 : _GEN_5725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5727 = 8'h55 == _match_key_qbytes_2_T_1 ? phv_data_85 : _GEN_5726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5728 = 8'h56 == _match_key_qbytes_2_T_1 ? phv_data_86 : _GEN_5727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5729 = 8'h57 == _match_key_qbytes_2_T_1 ? phv_data_87 : _GEN_5728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5730 = 8'h58 == _match_key_qbytes_2_T_1 ? phv_data_88 : _GEN_5729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5731 = 8'h59 == _match_key_qbytes_2_T_1 ? phv_data_89 : _GEN_5730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5732 = 8'h5a == _match_key_qbytes_2_T_1 ? phv_data_90 : _GEN_5731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5733 = 8'h5b == _match_key_qbytes_2_T_1 ? phv_data_91 : _GEN_5732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5734 = 8'h5c == _match_key_qbytes_2_T_1 ? phv_data_92 : _GEN_5733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5735 = 8'h5d == _match_key_qbytes_2_T_1 ? phv_data_93 : _GEN_5734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5736 = 8'h5e == _match_key_qbytes_2_T_1 ? phv_data_94 : _GEN_5735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5737 = 8'h5f == _match_key_qbytes_2_T_1 ? phv_data_95 : _GEN_5736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5738 = 8'h60 == _match_key_qbytes_2_T_1 ? phv_data_96 : _GEN_5737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5739 = 8'h61 == _match_key_qbytes_2_T_1 ? phv_data_97 : _GEN_5738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5740 = 8'h62 == _match_key_qbytes_2_T_1 ? phv_data_98 : _GEN_5739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5741 = 8'h63 == _match_key_qbytes_2_T_1 ? phv_data_99 : _GEN_5740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5742 = 8'h64 == _match_key_qbytes_2_T_1 ? phv_data_100 : _GEN_5741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5743 = 8'h65 == _match_key_qbytes_2_T_1 ? phv_data_101 : _GEN_5742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5744 = 8'h66 == _match_key_qbytes_2_T_1 ? phv_data_102 : _GEN_5743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5745 = 8'h67 == _match_key_qbytes_2_T_1 ? phv_data_103 : _GEN_5744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5746 = 8'h68 == _match_key_qbytes_2_T_1 ? phv_data_104 : _GEN_5745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5747 = 8'h69 == _match_key_qbytes_2_T_1 ? phv_data_105 : _GEN_5746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5748 = 8'h6a == _match_key_qbytes_2_T_1 ? phv_data_106 : _GEN_5747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5749 = 8'h6b == _match_key_qbytes_2_T_1 ? phv_data_107 : _GEN_5748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5750 = 8'h6c == _match_key_qbytes_2_T_1 ? phv_data_108 : _GEN_5749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5751 = 8'h6d == _match_key_qbytes_2_T_1 ? phv_data_109 : _GEN_5750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5752 = 8'h6e == _match_key_qbytes_2_T_1 ? phv_data_110 : _GEN_5751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5753 = 8'h6f == _match_key_qbytes_2_T_1 ? phv_data_111 : _GEN_5752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5754 = 8'h70 == _match_key_qbytes_2_T_1 ? phv_data_112 : _GEN_5753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5755 = 8'h71 == _match_key_qbytes_2_T_1 ? phv_data_113 : _GEN_5754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5756 = 8'h72 == _match_key_qbytes_2_T_1 ? phv_data_114 : _GEN_5755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5757 = 8'h73 == _match_key_qbytes_2_T_1 ? phv_data_115 : _GEN_5756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5758 = 8'h74 == _match_key_qbytes_2_T_1 ? phv_data_116 : _GEN_5757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5759 = 8'h75 == _match_key_qbytes_2_T_1 ? phv_data_117 : _GEN_5758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5760 = 8'h76 == _match_key_qbytes_2_T_1 ? phv_data_118 : _GEN_5759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5761 = 8'h77 == _match_key_qbytes_2_T_1 ? phv_data_119 : _GEN_5760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5762 = 8'h78 == _match_key_qbytes_2_T_1 ? phv_data_120 : _GEN_5761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5763 = 8'h79 == _match_key_qbytes_2_T_1 ? phv_data_121 : _GEN_5762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5764 = 8'h7a == _match_key_qbytes_2_T_1 ? phv_data_122 : _GEN_5763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5765 = 8'h7b == _match_key_qbytes_2_T_1 ? phv_data_123 : _GEN_5764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5766 = 8'h7c == _match_key_qbytes_2_T_1 ? phv_data_124 : _GEN_5765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5767 = 8'h7d == _match_key_qbytes_2_T_1 ? phv_data_125 : _GEN_5766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5768 = 8'h7e == _match_key_qbytes_2_T_1 ? phv_data_126 : _GEN_5767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5769 = 8'h7f == _match_key_qbytes_2_T_1 ? phv_data_127 : _GEN_5768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5770 = 8'h80 == _match_key_qbytes_2_T_1 ? phv_data_128 : _GEN_5769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5771 = 8'h81 == _match_key_qbytes_2_T_1 ? phv_data_129 : _GEN_5770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5772 = 8'h82 == _match_key_qbytes_2_T_1 ? phv_data_130 : _GEN_5771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5773 = 8'h83 == _match_key_qbytes_2_T_1 ? phv_data_131 : _GEN_5772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5774 = 8'h84 == _match_key_qbytes_2_T_1 ? phv_data_132 : _GEN_5773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5775 = 8'h85 == _match_key_qbytes_2_T_1 ? phv_data_133 : _GEN_5774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5776 = 8'h86 == _match_key_qbytes_2_T_1 ? phv_data_134 : _GEN_5775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5777 = 8'h87 == _match_key_qbytes_2_T_1 ? phv_data_135 : _GEN_5776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5778 = 8'h88 == _match_key_qbytes_2_T_1 ? phv_data_136 : _GEN_5777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5779 = 8'h89 == _match_key_qbytes_2_T_1 ? phv_data_137 : _GEN_5778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5780 = 8'h8a == _match_key_qbytes_2_T_1 ? phv_data_138 : _GEN_5779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5781 = 8'h8b == _match_key_qbytes_2_T_1 ? phv_data_139 : _GEN_5780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5782 = 8'h8c == _match_key_qbytes_2_T_1 ? phv_data_140 : _GEN_5781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5783 = 8'h8d == _match_key_qbytes_2_T_1 ? phv_data_141 : _GEN_5782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5784 = 8'h8e == _match_key_qbytes_2_T_1 ? phv_data_142 : _GEN_5783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5785 = 8'h8f == _match_key_qbytes_2_T_1 ? phv_data_143 : _GEN_5784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5786 = 8'h90 == _match_key_qbytes_2_T_1 ? phv_data_144 : _GEN_5785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5787 = 8'h91 == _match_key_qbytes_2_T_1 ? phv_data_145 : _GEN_5786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5788 = 8'h92 == _match_key_qbytes_2_T_1 ? phv_data_146 : _GEN_5787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5789 = 8'h93 == _match_key_qbytes_2_T_1 ? phv_data_147 : _GEN_5788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5790 = 8'h94 == _match_key_qbytes_2_T_1 ? phv_data_148 : _GEN_5789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5791 = 8'h95 == _match_key_qbytes_2_T_1 ? phv_data_149 : _GEN_5790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5792 = 8'h96 == _match_key_qbytes_2_T_1 ? phv_data_150 : _GEN_5791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5793 = 8'h97 == _match_key_qbytes_2_T_1 ? phv_data_151 : _GEN_5792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5794 = 8'h98 == _match_key_qbytes_2_T_1 ? phv_data_152 : _GEN_5793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5795 = 8'h99 == _match_key_qbytes_2_T_1 ? phv_data_153 : _GEN_5794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5796 = 8'h9a == _match_key_qbytes_2_T_1 ? phv_data_154 : _GEN_5795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5797 = 8'h9b == _match_key_qbytes_2_T_1 ? phv_data_155 : _GEN_5796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5798 = 8'h9c == _match_key_qbytes_2_T_1 ? phv_data_156 : _GEN_5797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5799 = 8'h9d == _match_key_qbytes_2_T_1 ? phv_data_157 : _GEN_5798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5800 = 8'h9e == _match_key_qbytes_2_T_1 ? phv_data_158 : _GEN_5799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5801 = 8'h9f == _match_key_qbytes_2_T_1 ? phv_data_159 : _GEN_5800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5802 = 8'ha0 == _match_key_qbytes_2_T_1 ? phv_data_160 : _GEN_5801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5803 = 8'ha1 == _match_key_qbytes_2_T_1 ? phv_data_161 : _GEN_5802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5804 = 8'ha2 == _match_key_qbytes_2_T_1 ? phv_data_162 : _GEN_5803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5805 = 8'ha3 == _match_key_qbytes_2_T_1 ? phv_data_163 : _GEN_5804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5806 = 8'ha4 == _match_key_qbytes_2_T_1 ? phv_data_164 : _GEN_5805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5807 = 8'ha5 == _match_key_qbytes_2_T_1 ? phv_data_165 : _GEN_5806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5808 = 8'ha6 == _match_key_qbytes_2_T_1 ? phv_data_166 : _GEN_5807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5809 = 8'ha7 == _match_key_qbytes_2_T_1 ? phv_data_167 : _GEN_5808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5810 = 8'ha8 == _match_key_qbytes_2_T_1 ? phv_data_168 : _GEN_5809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5811 = 8'ha9 == _match_key_qbytes_2_T_1 ? phv_data_169 : _GEN_5810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5812 = 8'haa == _match_key_qbytes_2_T_1 ? phv_data_170 : _GEN_5811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5813 = 8'hab == _match_key_qbytes_2_T_1 ? phv_data_171 : _GEN_5812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5814 = 8'hac == _match_key_qbytes_2_T_1 ? phv_data_172 : _GEN_5813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5815 = 8'had == _match_key_qbytes_2_T_1 ? phv_data_173 : _GEN_5814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5816 = 8'hae == _match_key_qbytes_2_T_1 ? phv_data_174 : _GEN_5815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5817 = 8'haf == _match_key_qbytes_2_T_1 ? phv_data_175 : _GEN_5816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5818 = 8'hb0 == _match_key_qbytes_2_T_1 ? phv_data_176 : _GEN_5817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5819 = 8'hb1 == _match_key_qbytes_2_T_1 ? phv_data_177 : _GEN_5818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5820 = 8'hb2 == _match_key_qbytes_2_T_1 ? phv_data_178 : _GEN_5819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5821 = 8'hb3 == _match_key_qbytes_2_T_1 ? phv_data_179 : _GEN_5820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5822 = 8'hb4 == _match_key_qbytes_2_T_1 ? phv_data_180 : _GEN_5821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5823 = 8'hb5 == _match_key_qbytes_2_T_1 ? phv_data_181 : _GEN_5822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5824 = 8'hb6 == _match_key_qbytes_2_T_1 ? phv_data_182 : _GEN_5823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5825 = 8'hb7 == _match_key_qbytes_2_T_1 ? phv_data_183 : _GEN_5824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5826 = 8'hb8 == _match_key_qbytes_2_T_1 ? phv_data_184 : _GEN_5825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5827 = 8'hb9 == _match_key_qbytes_2_T_1 ? phv_data_185 : _GEN_5826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5828 = 8'hba == _match_key_qbytes_2_T_1 ? phv_data_186 : _GEN_5827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5829 = 8'hbb == _match_key_qbytes_2_T_1 ? phv_data_187 : _GEN_5828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5830 = 8'hbc == _match_key_qbytes_2_T_1 ? phv_data_188 : _GEN_5829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5831 = 8'hbd == _match_key_qbytes_2_T_1 ? phv_data_189 : _GEN_5830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5832 = 8'hbe == _match_key_qbytes_2_T_1 ? phv_data_190 : _GEN_5831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5833 = 8'hbf == _match_key_qbytes_2_T_1 ? phv_data_191 : _GEN_5832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5834 = 8'hc0 == _match_key_qbytes_2_T_1 ? phv_data_192 : _GEN_5833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5835 = 8'hc1 == _match_key_qbytes_2_T_1 ? phv_data_193 : _GEN_5834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5836 = 8'hc2 == _match_key_qbytes_2_T_1 ? phv_data_194 : _GEN_5835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5837 = 8'hc3 == _match_key_qbytes_2_T_1 ? phv_data_195 : _GEN_5836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5838 = 8'hc4 == _match_key_qbytes_2_T_1 ? phv_data_196 : _GEN_5837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5839 = 8'hc5 == _match_key_qbytes_2_T_1 ? phv_data_197 : _GEN_5838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5840 = 8'hc6 == _match_key_qbytes_2_T_1 ? phv_data_198 : _GEN_5839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5841 = 8'hc7 == _match_key_qbytes_2_T_1 ? phv_data_199 : _GEN_5840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5842 = 8'hc8 == _match_key_qbytes_2_T_1 ? phv_data_200 : _GEN_5841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5843 = 8'hc9 == _match_key_qbytes_2_T_1 ? phv_data_201 : _GEN_5842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5844 = 8'hca == _match_key_qbytes_2_T_1 ? phv_data_202 : _GEN_5843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5845 = 8'hcb == _match_key_qbytes_2_T_1 ? phv_data_203 : _GEN_5844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5846 = 8'hcc == _match_key_qbytes_2_T_1 ? phv_data_204 : _GEN_5845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5847 = 8'hcd == _match_key_qbytes_2_T_1 ? phv_data_205 : _GEN_5846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5848 = 8'hce == _match_key_qbytes_2_T_1 ? phv_data_206 : _GEN_5847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5849 = 8'hcf == _match_key_qbytes_2_T_1 ? phv_data_207 : _GEN_5848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5850 = 8'hd0 == _match_key_qbytes_2_T_1 ? phv_data_208 : _GEN_5849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5851 = 8'hd1 == _match_key_qbytes_2_T_1 ? phv_data_209 : _GEN_5850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5852 = 8'hd2 == _match_key_qbytes_2_T_1 ? phv_data_210 : _GEN_5851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5853 = 8'hd3 == _match_key_qbytes_2_T_1 ? phv_data_211 : _GEN_5852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5854 = 8'hd4 == _match_key_qbytes_2_T_1 ? phv_data_212 : _GEN_5853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5855 = 8'hd5 == _match_key_qbytes_2_T_1 ? phv_data_213 : _GEN_5854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5856 = 8'hd6 == _match_key_qbytes_2_T_1 ? phv_data_214 : _GEN_5855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5857 = 8'hd7 == _match_key_qbytes_2_T_1 ? phv_data_215 : _GEN_5856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5858 = 8'hd8 == _match_key_qbytes_2_T_1 ? phv_data_216 : _GEN_5857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5859 = 8'hd9 == _match_key_qbytes_2_T_1 ? phv_data_217 : _GEN_5858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5860 = 8'hda == _match_key_qbytes_2_T_1 ? phv_data_218 : _GEN_5859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5861 = 8'hdb == _match_key_qbytes_2_T_1 ? phv_data_219 : _GEN_5860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5862 = 8'hdc == _match_key_qbytes_2_T_1 ? phv_data_220 : _GEN_5861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5863 = 8'hdd == _match_key_qbytes_2_T_1 ? phv_data_221 : _GEN_5862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5864 = 8'hde == _match_key_qbytes_2_T_1 ? phv_data_222 : _GEN_5863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5865 = 8'hdf == _match_key_qbytes_2_T_1 ? phv_data_223 : _GEN_5864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5866 = 8'he0 == _match_key_qbytes_2_T_1 ? phv_data_224 : _GEN_5865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5867 = 8'he1 == _match_key_qbytes_2_T_1 ? phv_data_225 : _GEN_5866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5868 = 8'he2 == _match_key_qbytes_2_T_1 ? phv_data_226 : _GEN_5867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5869 = 8'he3 == _match_key_qbytes_2_T_1 ? phv_data_227 : _GEN_5868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5870 = 8'he4 == _match_key_qbytes_2_T_1 ? phv_data_228 : _GEN_5869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5871 = 8'he5 == _match_key_qbytes_2_T_1 ? phv_data_229 : _GEN_5870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5872 = 8'he6 == _match_key_qbytes_2_T_1 ? phv_data_230 : _GEN_5871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5873 = 8'he7 == _match_key_qbytes_2_T_1 ? phv_data_231 : _GEN_5872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5874 = 8'he8 == _match_key_qbytes_2_T_1 ? phv_data_232 : _GEN_5873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5875 = 8'he9 == _match_key_qbytes_2_T_1 ? phv_data_233 : _GEN_5874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5876 = 8'hea == _match_key_qbytes_2_T_1 ? phv_data_234 : _GEN_5875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5877 = 8'heb == _match_key_qbytes_2_T_1 ? phv_data_235 : _GEN_5876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5878 = 8'hec == _match_key_qbytes_2_T_1 ? phv_data_236 : _GEN_5877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5879 = 8'hed == _match_key_qbytes_2_T_1 ? phv_data_237 : _GEN_5878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5880 = 8'hee == _match_key_qbytes_2_T_1 ? phv_data_238 : _GEN_5879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5881 = 8'hef == _match_key_qbytes_2_T_1 ? phv_data_239 : _GEN_5880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5882 = 8'hf0 == _match_key_qbytes_2_T_1 ? phv_data_240 : _GEN_5881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5883 = 8'hf1 == _match_key_qbytes_2_T_1 ? phv_data_241 : _GEN_5882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5884 = 8'hf2 == _match_key_qbytes_2_T_1 ? phv_data_242 : _GEN_5883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5885 = 8'hf3 == _match_key_qbytes_2_T_1 ? phv_data_243 : _GEN_5884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5886 = 8'hf4 == _match_key_qbytes_2_T_1 ? phv_data_244 : _GEN_5885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5887 = 8'hf5 == _match_key_qbytes_2_T_1 ? phv_data_245 : _GEN_5886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5888 = 8'hf6 == _match_key_qbytes_2_T_1 ? phv_data_246 : _GEN_5887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5889 = 8'hf7 == _match_key_qbytes_2_T_1 ? phv_data_247 : _GEN_5888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5890 = 8'hf8 == _match_key_qbytes_2_T_1 ? phv_data_248 : _GEN_5889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5891 = 8'hf9 == _match_key_qbytes_2_T_1 ? phv_data_249 : _GEN_5890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5892 = 8'hfa == _match_key_qbytes_2_T_1 ? phv_data_250 : _GEN_5891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5893 = 8'hfb == _match_key_qbytes_2_T_1 ? phv_data_251 : _GEN_5892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5894 = 8'hfc == _match_key_qbytes_2_T_1 ? phv_data_252 : _GEN_5893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5895 = 8'hfd == _match_key_qbytes_2_T_1 ? phv_data_253 : _GEN_5894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5896 = 8'hfe == _match_key_qbytes_2_T_1 ? phv_data_254 : _GEN_5895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5897 = 8'hff == _match_key_qbytes_2_T_1 ? phv_data_255 : _GEN_5896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_15142 = {{1'd0}, _match_key_qbytes_2_T_1}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5898 = 9'h100 == _GEN_15142 ? phv_data_256 : _GEN_5897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5899 = 9'h101 == _GEN_15142 ? phv_data_257 : _GEN_5898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5900 = 9'h102 == _GEN_15142 ? phv_data_258 : _GEN_5899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5901 = 9'h103 == _GEN_15142 ? phv_data_259 : _GEN_5900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5902 = 9'h104 == _GEN_15142 ? phv_data_260 : _GEN_5901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5903 = 9'h105 == _GEN_15142 ? phv_data_261 : _GEN_5902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5904 = 9'h106 == _GEN_15142 ? phv_data_262 : _GEN_5903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5905 = 9'h107 == _GEN_15142 ? phv_data_263 : _GEN_5904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5906 = 9'h108 == _GEN_15142 ? phv_data_264 : _GEN_5905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5907 = 9'h109 == _GEN_15142 ? phv_data_265 : _GEN_5906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5908 = 9'h10a == _GEN_15142 ? phv_data_266 : _GEN_5907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5909 = 9'h10b == _GEN_15142 ? phv_data_267 : _GEN_5908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5910 = 9'h10c == _GEN_15142 ? phv_data_268 : _GEN_5909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5911 = 9'h10d == _GEN_15142 ? phv_data_269 : _GEN_5910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5912 = 9'h10e == _GEN_15142 ? phv_data_270 : _GEN_5911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5913 = 9'h10f == _GEN_15142 ? phv_data_271 : _GEN_5912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5914 = 9'h110 == _GEN_15142 ? phv_data_272 : _GEN_5913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5915 = 9'h111 == _GEN_15142 ? phv_data_273 : _GEN_5914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5916 = 9'h112 == _GEN_15142 ? phv_data_274 : _GEN_5915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5917 = 9'h113 == _GEN_15142 ? phv_data_275 : _GEN_5916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5918 = 9'h114 == _GEN_15142 ? phv_data_276 : _GEN_5917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5919 = 9'h115 == _GEN_15142 ? phv_data_277 : _GEN_5918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5920 = 9'h116 == _GEN_15142 ? phv_data_278 : _GEN_5919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5921 = 9'h117 == _GEN_15142 ? phv_data_279 : _GEN_5920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5922 = 9'h118 == _GEN_15142 ? phv_data_280 : _GEN_5921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5923 = 9'h119 == _GEN_15142 ? phv_data_281 : _GEN_5922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5924 = 9'h11a == _GEN_15142 ? phv_data_282 : _GEN_5923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5925 = 9'h11b == _GEN_15142 ? phv_data_283 : _GEN_5924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5926 = 9'h11c == _GEN_15142 ? phv_data_284 : _GEN_5925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5927 = 9'h11d == _GEN_15142 ? phv_data_285 : _GEN_5926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5928 = 9'h11e == _GEN_15142 ? phv_data_286 : _GEN_5927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5929 = 9'h11f == _GEN_15142 ? phv_data_287 : _GEN_5928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5930 = 9'h120 == _GEN_15142 ? phv_data_288 : _GEN_5929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5931 = 9'h121 == _GEN_15142 ? phv_data_289 : _GEN_5930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5932 = 9'h122 == _GEN_15142 ? phv_data_290 : _GEN_5931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5933 = 9'h123 == _GEN_15142 ? phv_data_291 : _GEN_5932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5934 = 9'h124 == _GEN_15142 ? phv_data_292 : _GEN_5933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5935 = 9'h125 == _GEN_15142 ? phv_data_293 : _GEN_5934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5936 = 9'h126 == _GEN_15142 ? phv_data_294 : _GEN_5935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5937 = 9'h127 == _GEN_15142 ? phv_data_295 : _GEN_5936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5938 = 9'h128 == _GEN_15142 ? phv_data_296 : _GEN_5937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5939 = 9'h129 == _GEN_15142 ? phv_data_297 : _GEN_5938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5940 = 9'h12a == _GEN_15142 ? phv_data_298 : _GEN_5939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5941 = 9'h12b == _GEN_15142 ? phv_data_299 : _GEN_5940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5942 = 9'h12c == _GEN_15142 ? phv_data_300 : _GEN_5941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5943 = 9'h12d == _GEN_15142 ? phv_data_301 : _GEN_5942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5944 = 9'h12e == _GEN_15142 ? phv_data_302 : _GEN_5943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5945 = 9'h12f == _GEN_15142 ? phv_data_303 : _GEN_5944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5946 = 9'h130 == _GEN_15142 ? phv_data_304 : _GEN_5945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5947 = 9'h131 == _GEN_15142 ? phv_data_305 : _GEN_5946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5948 = 9'h132 == _GEN_15142 ? phv_data_306 : _GEN_5947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5949 = 9'h133 == _GEN_15142 ? phv_data_307 : _GEN_5948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5950 = 9'h134 == _GEN_15142 ? phv_data_308 : _GEN_5949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5951 = 9'h135 == _GEN_15142 ? phv_data_309 : _GEN_5950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5952 = 9'h136 == _GEN_15142 ? phv_data_310 : _GEN_5951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5953 = 9'h137 == _GEN_15142 ? phv_data_311 : _GEN_5952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5954 = 9'h138 == _GEN_15142 ? phv_data_312 : _GEN_5953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5955 = 9'h139 == _GEN_15142 ? phv_data_313 : _GEN_5954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5956 = 9'h13a == _GEN_15142 ? phv_data_314 : _GEN_5955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5957 = 9'h13b == _GEN_15142 ? phv_data_315 : _GEN_5956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5958 = 9'h13c == _GEN_15142 ? phv_data_316 : _GEN_5957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5959 = 9'h13d == _GEN_15142 ? phv_data_317 : _GEN_5958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5960 = 9'h13e == _GEN_15142 ? phv_data_318 : _GEN_5959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5961 = 9'h13f == _GEN_15142 ? phv_data_319 : _GEN_5960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5962 = 9'h140 == _GEN_15142 ? phv_data_320 : _GEN_5961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5963 = 9'h141 == _GEN_15142 ? phv_data_321 : _GEN_5962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5964 = 9'h142 == _GEN_15142 ? phv_data_322 : _GEN_5963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5965 = 9'h143 == _GEN_15142 ? phv_data_323 : _GEN_5964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5966 = 9'h144 == _GEN_15142 ? phv_data_324 : _GEN_5965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5967 = 9'h145 == _GEN_15142 ? phv_data_325 : _GEN_5966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5968 = 9'h146 == _GEN_15142 ? phv_data_326 : _GEN_5967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5969 = 9'h147 == _GEN_15142 ? phv_data_327 : _GEN_5968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5970 = 9'h148 == _GEN_15142 ? phv_data_328 : _GEN_5969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5971 = 9'h149 == _GEN_15142 ? phv_data_329 : _GEN_5970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5972 = 9'h14a == _GEN_15142 ? phv_data_330 : _GEN_5971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5973 = 9'h14b == _GEN_15142 ? phv_data_331 : _GEN_5972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5974 = 9'h14c == _GEN_15142 ? phv_data_332 : _GEN_5973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5975 = 9'h14d == _GEN_15142 ? phv_data_333 : _GEN_5974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5976 = 9'h14e == _GEN_15142 ? phv_data_334 : _GEN_5975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5977 = 9'h14f == _GEN_15142 ? phv_data_335 : _GEN_5976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5978 = 9'h150 == _GEN_15142 ? phv_data_336 : _GEN_5977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5979 = 9'h151 == _GEN_15142 ? phv_data_337 : _GEN_5978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5980 = 9'h152 == _GEN_15142 ? phv_data_338 : _GEN_5979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5981 = 9'h153 == _GEN_15142 ? phv_data_339 : _GEN_5980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5982 = 9'h154 == _GEN_15142 ? phv_data_340 : _GEN_5981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5983 = 9'h155 == _GEN_15142 ? phv_data_341 : _GEN_5982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5984 = 9'h156 == _GEN_15142 ? phv_data_342 : _GEN_5983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5985 = 9'h157 == _GEN_15142 ? phv_data_343 : _GEN_5984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5986 = 9'h158 == _GEN_15142 ? phv_data_344 : _GEN_5985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5987 = 9'h159 == _GEN_15142 ? phv_data_345 : _GEN_5986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5988 = 9'h15a == _GEN_15142 ? phv_data_346 : _GEN_5987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5989 = 9'h15b == _GEN_15142 ? phv_data_347 : _GEN_5988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5990 = 9'h15c == _GEN_15142 ? phv_data_348 : _GEN_5989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5991 = 9'h15d == _GEN_15142 ? phv_data_349 : _GEN_5990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5992 = 9'h15e == _GEN_15142 ? phv_data_350 : _GEN_5991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5993 = 9'h15f == _GEN_15142 ? phv_data_351 : _GEN_5992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5994 = 9'h160 == _GEN_15142 ? phv_data_352 : _GEN_5993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5995 = 9'h161 == _GEN_15142 ? phv_data_353 : _GEN_5994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5996 = 9'h162 == _GEN_15142 ? phv_data_354 : _GEN_5995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5997 = 9'h163 == _GEN_15142 ? phv_data_355 : _GEN_5996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5998 = 9'h164 == _GEN_15142 ? phv_data_356 : _GEN_5997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5999 = 9'h165 == _GEN_15142 ? phv_data_357 : _GEN_5998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6000 = 9'h166 == _GEN_15142 ? phv_data_358 : _GEN_5999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6001 = 9'h167 == _GEN_15142 ? phv_data_359 : _GEN_6000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6002 = 9'h168 == _GEN_15142 ? phv_data_360 : _GEN_6001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6003 = 9'h169 == _GEN_15142 ? phv_data_361 : _GEN_6002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6004 = 9'h16a == _GEN_15142 ? phv_data_362 : _GEN_6003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6005 = 9'h16b == _GEN_15142 ? phv_data_363 : _GEN_6004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6006 = 9'h16c == _GEN_15142 ? phv_data_364 : _GEN_6005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6007 = 9'h16d == _GEN_15142 ? phv_data_365 : _GEN_6006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6008 = 9'h16e == _GEN_15142 ? phv_data_366 : _GEN_6007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6009 = 9'h16f == _GEN_15142 ? phv_data_367 : _GEN_6008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6010 = 9'h170 == _GEN_15142 ? phv_data_368 : _GEN_6009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6011 = 9'h171 == _GEN_15142 ? phv_data_369 : _GEN_6010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6012 = 9'h172 == _GEN_15142 ? phv_data_370 : _GEN_6011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6013 = 9'h173 == _GEN_15142 ? phv_data_371 : _GEN_6012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6014 = 9'h174 == _GEN_15142 ? phv_data_372 : _GEN_6013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6015 = 9'h175 == _GEN_15142 ? phv_data_373 : _GEN_6014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6016 = 9'h176 == _GEN_15142 ? phv_data_374 : _GEN_6015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6017 = 9'h177 == _GEN_15142 ? phv_data_375 : _GEN_6016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6018 = 9'h178 == _GEN_15142 ? phv_data_376 : _GEN_6017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6019 = 9'h179 == _GEN_15142 ? phv_data_377 : _GEN_6018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6020 = 9'h17a == _GEN_15142 ? phv_data_378 : _GEN_6019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6021 = 9'h17b == _GEN_15142 ? phv_data_379 : _GEN_6020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6022 = 9'h17c == _GEN_15142 ? phv_data_380 : _GEN_6021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6023 = 9'h17d == _GEN_15142 ? phv_data_381 : _GEN_6022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6024 = 9'h17e == _GEN_15142 ? phv_data_382 : _GEN_6023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6025 = 9'h17f == _GEN_15142 ? phv_data_383 : _GEN_6024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6026 = 9'h180 == _GEN_15142 ? phv_data_384 : _GEN_6025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6027 = 9'h181 == _GEN_15142 ? phv_data_385 : _GEN_6026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6028 = 9'h182 == _GEN_15142 ? phv_data_386 : _GEN_6027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6029 = 9'h183 == _GEN_15142 ? phv_data_387 : _GEN_6028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6030 = 9'h184 == _GEN_15142 ? phv_data_388 : _GEN_6029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6031 = 9'h185 == _GEN_15142 ? phv_data_389 : _GEN_6030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6032 = 9'h186 == _GEN_15142 ? phv_data_390 : _GEN_6031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6033 = 9'h187 == _GEN_15142 ? phv_data_391 : _GEN_6032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6034 = 9'h188 == _GEN_15142 ? phv_data_392 : _GEN_6033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6035 = 9'h189 == _GEN_15142 ? phv_data_393 : _GEN_6034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6036 = 9'h18a == _GEN_15142 ? phv_data_394 : _GEN_6035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6037 = 9'h18b == _GEN_15142 ? phv_data_395 : _GEN_6036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6038 = 9'h18c == _GEN_15142 ? phv_data_396 : _GEN_6037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6039 = 9'h18d == _GEN_15142 ? phv_data_397 : _GEN_6038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6040 = 9'h18e == _GEN_15142 ? phv_data_398 : _GEN_6039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6041 = 9'h18f == _GEN_15142 ? phv_data_399 : _GEN_6040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6042 = 9'h190 == _GEN_15142 ? phv_data_400 : _GEN_6041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6043 = 9'h191 == _GEN_15142 ? phv_data_401 : _GEN_6042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6044 = 9'h192 == _GEN_15142 ? phv_data_402 : _GEN_6043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6045 = 9'h193 == _GEN_15142 ? phv_data_403 : _GEN_6044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6046 = 9'h194 == _GEN_15142 ? phv_data_404 : _GEN_6045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6047 = 9'h195 == _GEN_15142 ? phv_data_405 : _GEN_6046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6048 = 9'h196 == _GEN_15142 ? phv_data_406 : _GEN_6047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6049 = 9'h197 == _GEN_15142 ? phv_data_407 : _GEN_6048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6050 = 9'h198 == _GEN_15142 ? phv_data_408 : _GEN_6049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6051 = 9'h199 == _GEN_15142 ? phv_data_409 : _GEN_6050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6052 = 9'h19a == _GEN_15142 ? phv_data_410 : _GEN_6051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6053 = 9'h19b == _GEN_15142 ? phv_data_411 : _GEN_6052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6054 = 9'h19c == _GEN_15142 ? phv_data_412 : _GEN_6053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6055 = 9'h19d == _GEN_15142 ? phv_data_413 : _GEN_6054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6056 = 9'h19e == _GEN_15142 ? phv_data_414 : _GEN_6055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6057 = 9'h19f == _GEN_15142 ? phv_data_415 : _GEN_6056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6058 = 9'h1a0 == _GEN_15142 ? phv_data_416 : _GEN_6057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6059 = 9'h1a1 == _GEN_15142 ? phv_data_417 : _GEN_6058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6060 = 9'h1a2 == _GEN_15142 ? phv_data_418 : _GEN_6059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6061 = 9'h1a3 == _GEN_15142 ? phv_data_419 : _GEN_6060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6062 = 9'h1a4 == _GEN_15142 ? phv_data_420 : _GEN_6061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6063 = 9'h1a5 == _GEN_15142 ? phv_data_421 : _GEN_6062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6064 = 9'h1a6 == _GEN_15142 ? phv_data_422 : _GEN_6063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6065 = 9'h1a7 == _GEN_15142 ? phv_data_423 : _GEN_6064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6066 = 9'h1a8 == _GEN_15142 ? phv_data_424 : _GEN_6065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6067 = 9'h1a9 == _GEN_15142 ? phv_data_425 : _GEN_6066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6068 = 9'h1aa == _GEN_15142 ? phv_data_426 : _GEN_6067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6069 = 9'h1ab == _GEN_15142 ? phv_data_427 : _GEN_6068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6070 = 9'h1ac == _GEN_15142 ? phv_data_428 : _GEN_6069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6071 = 9'h1ad == _GEN_15142 ? phv_data_429 : _GEN_6070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6072 = 9'h1ae == _GEN_15142 ? phv_data_430 : _GEN_6071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6073 = 9'h1af == _GEN_15142 ? phv_data_431 : _GEN_6072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6074 = 9'h1b0 == _GEN_15142 ? phv_data_432 : _GEN_6073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6075 = 9'h1b1 == _GEN_15142 ? phv_data_433 : _GEN_6074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6076 = 9'h1b2 == _GEN_15142 ? phv_data_434 : _GEN_6075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6077 = 9'h1b3 == _GEN_15142 ? phv_data_435 : _GEN_6076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6078 = 9'h1b4 == _GEN_15142 ? phv_data_436 : _GEN_6077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6079 = 9'h1b5 == _GEN_15142 ? phv_data_437 : _GEN_6078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6080 = 9'h1b6 == _GEN_15142 ? phv_data_438 : _GEN_6079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6081 = 9'h1b7 == _GEN_15142 ? phv_data_439 : _GEN_6080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6082 = 9'h1b8 == _GEN_15142 ? phv_data_440 : _GEN_6081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6083 = 9'h1b9 == _GEN_15142 ? phv_data_441 : _GEN_6082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6084 = 9'h1ba == _GEN_15142 ? phv_data_442 : _GEN_6083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6085 = 9'h1bb == _GEN_15142 ? phv_data_443 : _GEN_6084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6086 = 9'h1bc == _GEN_15142 ? phv_data_444 : _GEN_6085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6087 = 9'h1bd == _GEN_15142 ? phv_data_445 : _GEN_6086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6088 = 9'h1be == _GEN_15142 ? phv_data_446 : _GEN_6087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6089 = 9'h1bf == _GEN_15142 ? phv_data_447 : _GEN_6088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6090 = 9'h1c0 == _GEN_15142 ? phv_data_448 : _GEN_6089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6091 = 9'h1c1 == _GEN_15142 ? phv_data_449 : _GEN_6090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6092 = 9'h1c2 == _GEN_15142 ? phv_data_450 : _GEN_6091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6093 = 9'h1c3 == _GEN_15142 ? phv_data_451 : _GEN_6092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6094 = 9'h1c4 == _GEN_15142 ? phv_data_452 : _GEN_6093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6095 = 9'h1c5 == _GEN_15142 ? phv_data_453 : _GEN_6094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6096 = 9'h1c6 == _GEN_15142 ? phv_data_454 : _GEN_6095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6097 = 9'h1c7 == _GEN_15142 ? phv_data_455 : _GEN_6096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6098 = 9'h1c8 == _GEN_15142 ? phv_data_456 : _GEN_6097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6099 = 9'h1c9 == _GEN_15142 ? phv_data_457 : _GEN_6098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6100 = 9'h1ca == _GEN_15142 ? phv_data_458 : _GEN_6099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6101 = 9'h1cb == _GEN_15142 ? phv_data_459 : _GEN_6100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6102 = 9'h1cc == _GEN_15142 ? phv_data_460 : _GEN_6101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6103 = 9'h1cd == _GEN_15142 ? phv_data_461 : _GEN_6102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6104 = 9'h1ce == _GEN_15142 ? phv_data_462 : _GEN_6103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6105 = 9'h1cf == _GEN_15142 ? phv_data_463 : _GEN_6104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6106 = 9'h1d0 == _GEN_15142 ? phv_data_464 : _GEN_6105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6107 = 9'h1d1 == _GEN_15142 ? phv_data_465 : _GEN_6106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6108 = 9'h1d2 == _GEN_15142 ? phv_data_466 : _GEN_6107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6109 = 9'h1d3 == _GEN_15142 ? phv_data_467 : _GEN_6108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6110 = 9'h1d4 == _GEN_15142 ? phv_data_468 : _GEN_6109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6111 = 9'h1d5 == _GEN_15142 ? phv_data_469 : _GEN_6110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6112 = 9'h1d6 == _GEN_15142 ? phv_data_470 : _GEN_6111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6113 = 9'h1d7 == _GEN_15142 ? phv_data_471 : _GEN_6112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6114 = 9'h1d8 == _GEN_15142 ? phv_data_472 : _GEN_6113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6115 = 9'h1d9 == _GEN_15142 ? phv_data_473 : _GEN_6114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6116 = 9'h1da == _GEN_15142 ? phv_data_474 : _GEN_6115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6117 = 9'h1db == _GEN_15142 ? phv_data_475 : _GEN_6116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6118 = 9'h1dc == _GEN_15142 ? phv_data_476 : _GEN_6117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6119 = 9'h1dd == _GEN_15142 ? phv_data_477 : _GEN_6118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6120 = 9'h1de == _GEN_15142 ? phv_data_478 : _GEN_6119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6121 = 9'h1df == _GEN_15142 ? phv_data_479 : _GEN_6120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6122 = 9'h1e0 == _GEN_15142 ? phv_data_480 : _GEN_6121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6123 = 9'h1e1 == _GEN_15142 ? phv_data_481 : _GEN_6122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6124 = 9'h1e2 == _GEN_15142 ? phv_data_482 : _GEN_6123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6125 = 9'h1e3 == _GEN_15142 ? phv_data_483 : _GEN_6124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6126 = 9'h1e4 == _GEN_15142 ? phv_data_484 : _GEN_6125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6127 = 9'h1e5 == _GEN_15142 ? phv_data_485 : _GEN_6126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6128 = 9'h1e6 == _GEN_15142 ? phv_data_486 : _GEN_6127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6129 = 9'h1e7 == _GEN_15142 ? phv_data_487 : _GEN_6128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6130 = 9'h1e8 == _GEN_15142 ? phv_data_488 : _GEN_6129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6131 = 9'h1e9 == _GEN_15142 ? phv_data_489 : _GEN_6130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6132 = 9'h1ea == _GEN_15142 ? phv_data_490 : _GEN_6131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6133 = 9'h1eb == _GEN_15142 ? phv_data_491 : _GEN_6132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6134 = 9'h1ec == _GEN_15142 ? phv_data_492 : _GEN_6133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6135 = 9'h1ed == _GEN_15142 ? phv_data_493 : _GEN_6134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6136 = 9'h1ee == _GEN_15142 ? phv_data_494 : _GEN_6135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6137 = 9'h1ef == _GEN_15142 ? phv_data_495 : _GEN_6136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6138 = 9'h1f0 == _GEN_15142 ? phv_data_496 : _GEN_6137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6139 = 9'h1f1 == _GEN_15142 ? phv_data_497 : _GEN_6138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6140 = 9'h1f2 == _GEN_15142 ? phv_data_498 : _GEN_6139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6141 = 9'h1f3 == _GEN_15142 ? phv_data_499 : _GEN_6140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6142 = 9'h1f4 == _GEN_15142 ? phv_data_500 : _GEN_6141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6143 = 9'h1f5 == _GEN_15142 ? phv_data_501 : _GEN_6142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6144 = 9'h1f6 == _GEN_15142 ? phv_data_502 : _GEN_6143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6145 = 9'h1f7 == _GEN_15142 ? phv_data_503 : _GEN_6144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6146 = 9'h1f8 == _GEN_15142 ? phv_data_504 : _GEN_6145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6147 = 9'h1f9 == _GEN_15142 ? phv_data_505 : _GEN_6146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6148 = 9'h1fa == _GEN_15142 ? phv_data_506 : _GEN_6147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6149 = 9'h1fb == _GEN_15142 ? phv_data_507 : _GEN_6148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6150 = 9'h1fc == _GEN_15142 ? phv_data_508 : _GEN_6149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6151 = 9'h1fd == _GEN_15142 ? phv_data_509 : _GEN_6150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6152 = 9'h1fe == _GEN_15142 ? phv_data_510 : _GEN_6151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6153 = 9'h1ff == _GEN_15142 ? phv_data_511 : _GEN_6152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_2_T_3 = {_GEN_5641,_GEN_6153,_GEN_4617,_GEN_5129}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_2 = local_offset_2 < end_offset ? _match_key_qbytes_2_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_3 = 8'hc + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_3_hi = local_offset_3[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_3_T = {match_key_qbytes_3_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_3_T_1 = {match_key_qbytes_3_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_3_T_2 = {match_key_qbytes_3_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_6156 = 8'h1 == _match_key_qbytes_3_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6157 = 8'h2 == _match_key_qbytes_3_T_2 ? phv_data_2 : _GEN_6156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6158 = 8'h3 == _match_key_qbytes_3_T_2 ? phv_data_3 : _GEN_6157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6159 = 8'h4 == _match_key_qbytes_3_T_2 ? phv_data_4 : _GEN_6158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6160 = 8'h5 == _match_key_qbytes_3_T_2 ? phv_data_5 : _GEN_6159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6161 = 8'h6 == _match_key_qbytes_3_T_2 ? phv_data_6 : _GEN_6160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6162 = 8'h7 == _match_key_qbytes_3_T_2 ? phv_data_7 : _GEN_6161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6163 = 8'h8 == _match_key_qbytes_3_T_2 ? phv_data_8 : _GEN_6162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6164 = 8'h9 == _match_key_qbytes_3_T_2 ? phv_data_9 : _GEN_6163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6165 = 8'ha == _match_key_qbytes_3_T_2 ? phv_data_10 : _GEN_6164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6166 = 8'hb == _match_key_qbytes_3_T_2 ? phv_data_11 : _GEN_6165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6167 = 8'hc == _match_key_qbytes_3_T_2 ? phv_data_12 : _GEN_6166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6168 = 8'hd == _match_key_qbytes_3_T_2 ? phv_data_13 : _GEN_6167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6169 = 8'he == _match_key_qbytes_3_T_2 ? phv_data_14 : _GEN_6168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6170 = 8'hf == _match_key_qbytes_3_T_2 ? phv_data_15 : _GEN_6169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6171 = 8'h10 == _match_key_qbytes_3_T_2 ? phv_data_16 : _GEN_6170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6172 = 8'h11 == _match_key_qbytes_3_T_2 ? phv_data_17 : _GEN_6171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6173 = 8'h12 == _match_key_qbytes_3_T_2 ? phv_data_18 : _GEN_6172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6174 = 8'h13 == _match_key_qbytes_3_T_2 ? phv_data_19 : _GEN_6173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6175 = 8'h14 == _match_key_qbytes_3_T_2 ? phv_data_20 : _GEN_6174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6176 = 8'h15 == _match_key_qbytes_3_T_2 ? phv_data_21 : _GEN_6175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6177 = 8'h16 == _match_key_qbytes_3_T_2 ? phv_data_22 : _GEN_6176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6178 = 8'h17 == _match_key_qbytes_3_T_2 ? phv_data_23 : _GEN_6177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6179 = 8'h18 == _match_key_qbytes_3_T_2 ? phv_data_24 : _GEN_6178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6180 = 8'h19 == _match_key_qbytes_3_T_2 ? phv_data_25 : _GEN_6179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6181 = 8'h1a == _match_key_qbytes_3_T_2 ? phv_data_26 : _GEN_6180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6182 = 8'h1b == _match_key_qbytes_3_T_2 ? phv_data_27 : _GEN_6181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6183 = 8'h1c == _match_key_qbytes_3_T_2 ? phv_data_28 : _GEN_6182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6184 = 8'h1d == _match_key_qbytes_3_T_2 ? phv_data_29 : _GEN_6183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6185 = 8'h1e == _match_key_qbytes_3_T_2 ? phv_data_30 : _GEN_6184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6186 = 8'h1f == _match_key_qbytes_3_T_2 ? phv_data_31 : _GEN_6185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6187 = 8'h20 == _match_key_qbytes_3_T_2 ? phv_data_32 : _GEN_6186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6188 = 8'h21 == _match_key_qbytes_3_T_2 ? phv_data_33 : _GEN_6187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6189 = 8'h22 == _match_key_qbytes_3_T_2 ? phv_data_34 : _GEN_6188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6190 = 8'h23 == _match_key_qbytes_3_T_2 ? phv_data_35 : _GEN_6189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6191 = 8'h24 == _match_key_qbytes_3_T_2 ? phv_data_36 : _GEN_6190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6192 = 8'h25 == _match_key_qbytes_3_T_2 ? phv_data_37 : _GEN_6191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6193 = 8'h26 == _match_key_qbytes_3_T_2 ? phv_data_38 : _GEN_6192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6194 = 8'h27 == _match_key_qbytes_3_T_2 ? phv_data_39 : _GEN_6193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6195 = 8'h28 == _match_key_qbytes_3_T_2 ? phv_data_40 : _GEN_6194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6196 = 8'h29 == _match_key_qbytes_3_T_2 ? phv_data_41 : _GEN_6195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6197 = 8'h2a == _match_key_qbytes_3_T_2 ? phv_data_42 : _GEN_6196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6198 = 8'h2b == _match_key_qbytes_3_T_2 ? phv_data_43 : _GEN_6197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6199 = 8'h2c == _match_key_qbytes_3_T_2 ? phv_data_44 : _GEN_6198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6200 = 8'h2d == _match_key_qbytes_3_T_2 ? phv_data_45 : _GEN_6199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6201 = 8'h2e == _match_key_qbytes_3_T_2 ? phv_data_46 : _GEN_6200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6202 = 8'h2f == _match_key_qbytes_3_T_2 ? phv_data_47 : _GEN_6201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6203 = 8'h30 == _match_key_qbytes_3_T_2 ? phv_data_48 : _GEN_6202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6204 = 8'h31 == _match_key_qbytes_3_T_2 ? phv_data_49 : _GEN_6203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6205 = 8'h32 == _match_key_qbytes_3_T_2 ? phv_data_50 : _GEN_6204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6206 = 8'h33 == _match_key_qbytes_3_T_2 ? phv_data_51 : _GEN_6205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6207 = 8'h34 == _match_key_qbytes_3_T_2 ? phv_data_52 : _GEN_6206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6208 = 8'h35 == _match_key_qbytes_3_T_2 ? phv_data_53 : _GEN_6207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6209 = 8'h36 == _match_key_qbytes_3_T_2 ? phv_data_54 : _GEN_6208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6210 = 8'h37 == _match_key_qbytes_3_T_2 ? phv_data_55 : _GEN_6209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6211 = 8'h38 == _match_key_qbytes_3_T_2 ? phv_data_56 : _GEN_6210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6212 = 8'h39 == _match_key_qbytes_3_T_2 ? phv_data_57 : _GEN_6211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6213 = 8'h3a == _match_key_qbytes_3_T_2 ? phv_data_58 : _GEN_6212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6214 = 8'h3b == _match_key_qbytes_3_T_2 ? phv_data_59 : _GEN_6213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6215 = 8'h3c == _match_key_qbytes_3_T_2 ? phv_data_60 : _GEN_6214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6216 = 8'h3d == _match_key_qbytes_3_T_2 ? phv_data_61 : _GEN_6215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6217 = 8'h3e == _match_key_qbytes_3_T_2 ? phv_data_62 : _GEN_6216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6218 = 8'h3f == _match_key_qbytes_3_T_2 ? phv_data_63 : _GEN_6217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6219 = 8'h40 == _match_key_qbytes_3_T_2 ? phv_data_64 : _GEN_6218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6220 = 8'h41 == _match_key_qbytes_3_T_2 ? phv_data_65 : _GEN_6219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6221 = 8'h42 == _match_key_qbytes_3_T_2 ? phv_data_66 : _GEN_6220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6222 = 8'h43 == _match_key_qbytes_3_T_2 ? phv_data_67 : _GEN_6221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6223 = 8'h44 == _match_key_qbytes_3_T_2 ? phv_data_68 : _GEN_6222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6224 = 8'h45 == _match_key_qbytes_3_T_2 ? phv_data_69 : _GEN_6223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6225 = 8'h46 == _match_key_qbytes_3_T_2 ? phv_data_70 : _GEN_6224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6226 = 8'h47 == _match_key_qbytes_3_T_2 ? phv_data_71 : _GEN_6225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6227 = 8'h48 == _match_key_qbytes_3_T_2 ? phv_data_72 : _GEN_6226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6228 = 8'h49 == _match_key_qbytes_3_T_2 ? phv_data_73 : _GEN_6227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6229 = 8'h4a == _match_key_qbytes_3_T_2 ? phv_data_74 : _GEN_6228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6230 = 8'h4b == _match_key_qbytes_3_T_2 ? phv_data_75 : _GEN_6229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6231 = 8'h4c == _match_key_qbytes_3_T_2 ? phv_data_76 : _GEN_6230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6232 = 8'h4d == _match_key_qbytes_3_T_2 ? phv_data_77 : _GEN_6231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6233 = 8'h4e == _match_key_qbytes_3_T_2 ? phv_data_78 : _GEN_6232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6234 = 8'h4f == _match_key_qbytes_3_T_2 ? phv_data_79 : _GEN_6233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6235 = 8'h50 == _match_key_qbytes_3_T_2 ? phv_data_80 : _GEN_6234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6236 = 8'h51 == _match_key_qbytes_3_T_2 ? phv_data_81 : _GEN_6235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6237 = 8'h52 == _match_key_qbytes_3_T_2 ? phv_data_82 : _GEN_6236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6238 = 8'h53 == _match_key_qbytes_3_T_2 ? phv_data_83 : _GEN_6237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6239 = 8'h54 == _match_key_qbytes_3_T_2 ? phv_data_84 : _GEN_6238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6240 = 8'h55 == _match_key_qbytes_3_T_2 ? phv_data_85 : _GEN_6239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6241 = 8'h56 == _match_key_qbytes_3_T_2 ? phv_data_86 : _GEN_6240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6242 = 8'h57 == _match_key_qbytes_3_T_2 ? phv_data_87 : _GEN_6241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6243 = 8'h58 == _match_key_qbytes_3_T_2 ? phv_data_88 : _GEN_6242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6244 = 8'h59 == _match_key_qbytes_3_T_2 ? phv_data_89 : _GEN_6243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6245 = 8'h5a == _match_key_qbytes_3_T_2 ? phv_data_90 : _GEN_6244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6246 = 8'h5b == _match_key_qbytes_3_T_2 ? phv_data_91 : _GEN_6245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6247 = 8'h5c == _match_key_qbytes_3_T_2 ? phv_data_92 : _GEN_6246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6248 = 8'h5d == _match_key_qbytes_3_T_2 ? phv_data_93 : _GEN_6247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6249 = 8'h5e == _match_key_qbytes_3_T_2 ? phv_data_94 : _GEN_6248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6250 = 8'h5f == _match_key_qbytes_3_T_2 ? phv_data_95 : _GEN_6249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6251 = 8'h60 == _match_key_qbytes_3_T_2 ? phv_data_96 : _GEN_6250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6252 = 8'h61 == _match_key_qbytes_3_T_2 ? phv_data_97 : _GEN_6251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6253 = 8'h62 == _match_key_qbytes_3_T_2 ? phv_data_98 : _GEN_6252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6254 = 8'h63 == _match_key_qbytes_3_T_2 ? phv_data_99 : _GEN_6253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6255 = 8'h64 == _match_key_qbytes_3_T_2 ? phv_data_100 : _GEN_6254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6256 = 8'h65 == _match_key_qbytes_3_T_2 ? phv_data_101 : _GEN_6255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6257 = 8'h66 == _match_key_qbytes_3_T_2 ? phv_data_102 : _GEN_6256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6258 = 8'h67 == _match_key_qbytes_3_T_2 ? phv_data_103 : _GEN_6257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6259 = 8'h68 == _match_key_qbytes_3_T_2 ? phv_data_104 : _GEN_6258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6260 = 8'h69 == _match_key_qbytes_3_T_2 ? phv_data_105 : _GEN_6259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6261 = 8'h6a == _match_key_qbytes_3_T_2 ? phv_data_106 : _GEN_6260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6262 = 8'h6b == _match_key_qbytes_3_T_2 ? phv_data_107 : _GEN_6261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6263 = 8'h6c == _match_key_qbytes_3_T_2 ? phv_data_108 : _GEN_6262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6264 = 8'h6d == _match_key_qbytes_3_T_2 ? phv_data_109 : _GEN_6263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6265 = 8'h6e == _match_key_qbytes_3_T_2 ? phv_data_110 : _GEN_6264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6266 = 8'h6f == _match_key_qbytes_3_T_2 ? phv_data_111 : _GEN_6265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6267 = 8'h70 == _match_key_qbytes_3_T_2 ? phv_data_112 : _GEN_6266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6268 = 8'h71 == _match_key_qbytes_3_T_2 ? phv_data_113 : _GEN_6267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6269 = 8'h72 == _match_key_qbytes_3_T_2 ? phv_data_114 : _GEN_6268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6270 = 8'h73 == _match_key_qbytes_3_T_2 ? phv_data_115 : _GEN_6269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6271 = 8'h74 == _match_key_qbytes_3_T_2 ? phv_data_116 : _GEN_6270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6272 = 8'h75 == _match_key_qbytes_3_T_2 ? phv_data_117 : _GEN_6271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6273 = 8'h76 == _match_key_qbytes_3_T_2 ? phv_data_118 : _GEN_6272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6274 = 8'h77 == _match_key_qbytes_3_T_2 ? phv_data_119 : _GEN_6273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6275 = 8'h78 == _match_key_qbytes_3_T_2 ? phv_data_120 : _GEN_6274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6276 = 8'h79 == _match_key_qbytes_3_T_2 ? phv_data_121 : _GEN_6275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6277 = 8'h7a == _match_key_qbytes_3_T_2 ? phv_data_122 : _GEN_6276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6278 = 8'h7b == _match_key_qbytes_3_T_2 ? phv_data_123 : _GEN_6277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6279 = 8'h7c == _match_key_qbytes_3_T_2 ? phv_data_124 : _GEN_6278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6280 = 8'h7d == _match_key_qbytes_3_T_2 ? phv_data_125 : _GEN_6279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6281 = 8'h7e == _match_key_qbytes_3_T_2 ? phv_data_126 : _GEN_6280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6282 = 8'h7f == _match_key_qbytes_3_T_2 ? phv_data_127 : _GEN_6281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6283 = 8'h80 == _match_key_qbytes_3_T_2 ? phv_data_128 : _GEN_6282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6284 = 8'h81 == _match_key_qbytes_3_T_2 ? phv_data_129 : _GEN_6283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6285 = 8'h82 == _match_key_qbytes_3_T_2 ? phv_data_130 : _GEN_6284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6286 = 8'h83 == _match_key_qbytes_3_T_2 ? phv_data_131 : _GEN_6285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6287 = 8'h84 == _match_key_qbytes_3_T_2 ? phv_data_132 : _GEN_6286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6288 = 8'h85 == _match_key_qbytes_3_T_2 ? phv_data_133 : _GEN_6287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6289 = 8'h86 == _match_key_qbytes_3_T_2 ? phv_data_134 : _GEN_6288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6290 = 8'h87 == _match_key_qbytes_3_T_2 ? phv_data_135 : _GEN_6289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6291 = 8'h88 == _match_key_qbytes_3_T_2 ? phv_data_136 : _GEN_6290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6292 = 8'h89 == _match_key_qbytes_3_T_2 ? phv_data_137 : _GEN_6291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6293 = 8'h8a == _match_key_qbytes_3_T_2 ? phv_data_138 : _GEN_6292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6294 = 8'h8b == _match_key_qbytes_3_T_2 ? phv_data_139 : _GEN_6293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6295 = 8'h8c == _match_key_qbytes_3_T_2 ? phv_data_140 : _GEN_6294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6296 = 8'h8d == _match_key_qbytes_3_T_2 ? phv_data_141 : _GEN_6295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6297 = 8'h8e == _match_key_qbytes_3_T_2 ? phv_data_142 : _GEN_6296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6298 = 8'h8f == _match_key_qbytes_3_T_2 ? phv_data_143 : _GEN_6297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6299 = 8'h90 == _match_key_qbytes_3_T_2 ? phv_data_144 : _GEN_6298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6300 = 8'h91 == _match_key_qbytes_3_T_2 ? phv_data_145 : _GEN_6299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6301 = 8'h92 == _match_key_qbytes_3_T_2 ? phv_data_146 : _GEN_6300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6302 = 8'h93 == _match_key_qbytes_3_T_2 ? phv_data_147 : _GEN_6301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6303 = 8'h94 == _match_key_qbytes_3_T_2 ? phv_data_148 : _GEN_6302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6304 = 8'h95 == _match_key_qbytes_3_T_2 ? phv_data_149 : _GEN_6303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6305 = 8'h96 == _match_key_qbytes_3_T_2 ? phv_data_150 : _GEN_6304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6306 = 8'h97 == _match_key_qbytes_3_T_2 ? phv_data_151 : _GEN_6305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6307 = 8'h98 == _match_key_qbytes_3_T_2 ? phv_data_152 : _GEN_6306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6308 = 8'h99 == _match_key_qbytes_3_T_2 ? phv_data_153 : _GEN_6307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6309 = 8'h9a == _match_key_qbytes_3_T_2 ? phv_data_154 : _GEN_6308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6310 = 8'h9b == _match_key_qbytes_3_T_2 ? phv_data_155 : _GEN_6309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6311 = 8'h9c == _match_key_qbytes_3_T_2 ? phv_data_156 : _GEN_6310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6312 = 8'h9d == _match_key_qbytes_3_T_2 ? phv_data_157 : _GEN_6311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6313 = 8'h9e == _match_key_qbytes_3_T_2 ? phv_data_158 : _GEN_6312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6314 = 8'h9f == _match_key_qbytes_3_T_2 ? phv_data_159 : _GEN_6313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6315 = 8'ha0 == _match_key_qbytes_3_T_2 ? phv_data_160 : _GEN_6314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6316 = 8'ha1 == _match_key_qbytes_3_T_2 ? phv_data_161 : _GEN_6315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6317 = 8'ha2 == _match_key_qbytes_3_T_2 ? phv_data_162 : _GEN_6316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6318 = 8'ha3 == _match_key_qbytes_3_T_2 ? phv_data_163 : _GEN_6317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6319 = 8'ha4 == _match_key_qbytes_3_T_2 ? phv_data_164 : _GEN_6318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6320 = 8'ha5 == _match_key_qbytes_3_T_2 ? phv_data_165 : _GEN_6319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6321 = 8'ha6 == _match_key_qbytes_3_T_2 ? phv_data_166 : _GEN_6320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6322 = 8'ha7 == _match_key_qbytes_3_T_2 ? phv_data_167 : _GEN_6321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6323 = 8'ha8 == _match_key_qbytes_3_T_2 ? phv_data_168 : _GEN_6322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6324 = 8'ha9 == _match_key_qbytes_3_T_2 ? phv_data_169 : _GEN_6323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6325 = 8'haa == _match_key_qbytes_3_T_2 ? phv_data_170 : _GEN_6324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6326 = 8'hab == _match_key_qbytes_3_T_2 ? phv_data_171 : _GEN_6325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6327 = 8'hac == _match_key_qbytes_3_T_2 ? phv_data_172 : _GEN_6326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6328 = 8'had == _match_key_qbytes_3_T_2 ? phv_data_173 : _GEN_6327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6329 = 8'hae == _match_key_qbytes_3_T_2 ? phv_data_174 : _GEN_6328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6330 = 8'haf == _match_key_qbytes_3_T_2 ? phv_data_175 : _GEN_6329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6331 = 8'hb0 == _match_key_qbytes_3_T_2 ? phv_data_176 : _GEN_6330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6332 = 8'hb1 == _match_key_qbytes_3_T_2 ? phv_data_177 : _GEN_6331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6333 = 8'hb2 == _match_key_qbytes_3_T_2 ? phv_data_178 : _GEN_6332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6334 = 8'hb3 == _match_key_qbytes_3_T_2 ? phv_data_179 : _GEN_6333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6335 = 8'hb4 == _match_key_qbytes_3_T_2 ? phv_data_180 : _GEN_6334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6336 = 8'hb5 == _match_key_qbytes_3_T_2 ? phv_data_181 : _GEN_6335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6337 = 8'hb6 == _match_key_qbytes_3_T_2 ? phv_data_182 : _GEN_6336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6338 = 8'hb7 == _match_key_qbytes_3_T_2 ? phv_data_183 : _GEN_6337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6339 = 8'hb8 == _match_key_qbytes_3_T_2 ? phv_data_184 : _GEN_6338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6340 = 8'hb9 == _match_key_qbytes_3_T_2 ? phv_data_185 : _GEN_6339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6341 = 8'hba == _match_key_qbytes_3_T_2 ? phv_data_186 : _GEN_6340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6342 = 8'hbb == _match_key_qbytes_3_T_2 ? phv_data_187 : _GEN_6341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6343 = 8'hbc == _match_key_qbytes_3_T_2 ? phv_data_188 : _GEN_6342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6344 = 8'hbd == _match_key_qbytes_3_T_2 ? phv_data_189 : _GEN_6343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6345 = 8'hbe == _match_key_qbytes_3_T_2 ? phv_data_190 : _GEN_6344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6346 = 8'hbf == _match_key_qbytes_3_T_2 ? phv_data_191 : _GEN_6345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6347 = 8'hc0 == _match_key_qbytes_3_T_2 ? phv_data_192 : _GEN_6346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6348 = 8'hc1 == _match_key_qbytes_3_T_2 ? phv_data_193 : _GEN_6347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6349 = 8'hc2 == _match_key_qbytes_3_T_2 ? phv_data_194 : _GEN_6348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6350 = 8'hc3 == _match_key_qbytes_3_T_2 ? phv_data_195 : _GEN_6349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6351 = 8'hc4 == _match_key_qbytes_3_T_2 ? phv_data_196 : _GEN_6350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6352 = 8'hc5 == _match_key_qbytes_3_T_2 ? phv_data_197 : _GEN_6351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6353 = 8'hc6 == _match_key_qbytes_3_T_2 ? phv_data_198 : _GEN_6352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6354 = 8'hc7 == _match_key_qbytes_3_T_2 ? phv_data_199 : _GEN_6353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6355 = 8'hc8 == _match_key_qbytes_3_T_2 ? phv_data_200 : _GEN_6354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6356 = 8'hc9 == _match_key_qbytes_3_T_2 ? phv_data_201 : _GEN_6355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6357 = 8'hca == _match_key_qbytes_3_T_2 ? phv_data_202 : _GEN_6356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6358 = 8'hcb == _match_key_qbytes_3_T_2 ? phv_data_203 : _GEN_6357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6359 = 8'hcc == _match_key_qbytes_3_T_2 ? phv_data_204 : _GEN_6358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6360 = 8'hcd == _match_key_qbytes_3_T_2 ? phv_data_205 : _GEN_6359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6361 = 8'hce == _match_key_qbytes_3_T_2 ? phv_data_206 : _GEN_6360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6362 = 8'hcf == _match_key_qbytes_3_T_2 ? phv_data_207 : _GEN_6361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6363 = 8'hd0 == _match_key_qbytes_3_T_2 ? phv_data_208 : _GEN_6362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6364 = 8'hd1 == _match_key_qbytes_3_T_2 ? phv_data_209 : _GEN_6363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6365 = 8'hd2 == _match_key_qbytes_3_T_2 ? phv_data_210 : _GEN_6364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6366 = 8'hd3 == _match_key_qbytes_3_T_2 ? phv_data_211 : _GEN_6365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6367 = 8'hd4 == _match_key_qbytes_3_T_2 ? phv_data_212 : _GEN_6366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6368 = 8'hd5 == _match_key_qbytes_3_T_2 ? phv_data_213 : _GEN_6367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6369 = 8'hd6 == _match_key_qbytes_3_T_2 ? phv_data_214 : _GEN_6368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6370 = 8'hd7 == _match_key_qbytes_3_T_2 ? phv_data_215 : _GEN_6369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6371 = 8'hd8 == _match_key_qbytes_3_T_2 ? phv_data_216 : _GEN_6370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6372 = 8'hd9 == _match_key_qbytes_3_T_2 ? phv_data_217 : _GEN_6371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6373 = 8'hda == _match_key_qbytes_3_T_2 ? phv_data_218 : _GEN_6372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6374 = 8'hdb == _match_key_qbytes_3_T_2 ? phv_data_219 : _GEN_6373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6375 = 8'hdc == _match_key_qbytes_3_T_2 ? phv_data_220 : _GEN_6374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6376 = 8'hdd == _match_key_qbytes_3_T_2 ? phv_data_221 : _GEN_6375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6377 = 8'hde == _match_key_qbytes_3_T_2 ? phv_data_222 : _GEN_6376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6378 = 8'hdf == _match_key_qbytes_3_T_2 ? phv_data_223 : _GEN_6377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6379 = 8'he0 == _match_key_qbytes_3_T_2 ? phv_data_224 : _GEN_6378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6380 = 8'he1 == _match_key_qbytes_3_T_2 ? phv_data_225 : _GEN_6379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6381 = 8'he2 == _match_key_qbytes_3_T_2 ? phv_data_226 : _GEN_6380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6382 = 8'he3 == _match_key_qbytes_3_T_2 ? phv_data_227 : _GEN_6381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6383 = 8'he4 == _match_key_qbytes_3_T_2 ? phv_data_228 : _GEN_6382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6384 = 8'he5 == _match_key_qbytes_3_T_2 ? phv_data_229 : _GEN_6383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6385 = 8'he6 == _match_key_qbytes_3_T_2 ? phv_data_230 : _GEN_6384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6386 = 8'he7 == _match_key_qbytes_3_T_2 ? phv_data_231 : _GEN_6385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6387 = 8'he8 == _match_key_qbytes_3_T_2 ? phv_data_232 : _GEN_6386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6388 = 8'he9 == _match_key_qbytes_3_T_2 ? phv_data_233 : _GEN_6387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6389 = 8'hea == _match_key_qbytes_3_T_2 ? phv_data_234 : _GEN_6388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6390 = 8'heb == _match_key_qbytes_3_T_2 ? phv_data_235 : _GEN_6389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6391 = 8'hec == _match_key_qbytes_3_T_2 ? phv_data_236 : _GEN_6390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6392 = 8'hed == _match_key_qbytes_3_T_2 ? phv_data_237 : _GEN_6391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6393 = 8'hee == _match_key_qbytes_3_T_2 ? phv_data_238 : _GEN_6392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6394 = 8'hef == _match_key_qbytes_3_T_2 ? phv_data_239 : _GEN_6393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6395 = 8'hf0 == _match_key_qbytes_3_T_2 ? phv_data_240 : _GEN_6394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6396 = 8'hf1 == _match_key_qbytes_3_T_2 ? phv_data_241 : _GEN_6395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6397 = 8'hf2 == _match_key_qbytes_3_T_2 ? phv_data_242 : _GEN_6396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6398 = 8'hf3 == _match_key_qbytes_3_T_2 ? phv_data_243 : _GEN_6397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6399 = 8'hf4 == _match_key_qbytes_3_T_2 ? phv_data_244 : _GEN_6398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6400 = 8'hf5 == _match_key_qbytes_3_T_2 ? phv_data_245 : _GEN_6399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6401 = 8'hf6 == _match_key_qbytes_3_T_2 ? phv_data_246 : _GEN_6400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6402 = 8'hf7 == _match_key_qbytes_3_T_2 ? phv_data_247 : _GEN_6401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6403 = 8'hf8 == _match_key_qbytes_3_T_2 ? phv_data_248 : _GEN_6402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6404 = 8'hf9 == _match_key_qbytes_3_T_2 ? phv_data_249 : _GEN_6403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6405 = 8'hfa == _match_key_qbytes_3_T_2 ? phv_data_250 : _GEN_6404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6406 = 8'hfb == _match_key_qbytes_3_T_2 ? phv_data_251 : _GEN_6405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6407 = 8'hfc == _match_key_qbytes_3_T_2 ? phv_data_252 : _GEN_6406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6408 = 8'hfd == _match_key_qbytes_3_T_2 ? phv_data_253 : _GEN_6407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6409 = 8'hfe == _match_key_qbytes_3_T_2 ? phv_data_254 : _GEN_6408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6410 = 8'hff == _match_key_qbytes_3_T_2 ? phv_data_255 : _GEN_6409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_15398 = {{1'd0}, _match_key_qbytes_3_T_2}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6411 = 9'h100 == _GEN_15398 ? phv_data_256 : _GEN_6410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6412 = 9'h101 == _GEN_15398 ? phv_data_257 : _GEN_6411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6413 = 9'h102 == _GEN_15398 ? phv_data_258 : _GEN_6412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6414 = 9'h103 == _GEN_15398 ? phv_data_259 : _GEN_6413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6415 = 9'h104 == _GEN_15398 ? phv_data_260 : _GEN_6414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6416 = 9'h105 == _GEN_15398 ? phv_data_261 : _GEN_6415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6417 = 9'h106 == _GEN_15398 ? phv_data_262 : _GEN_6416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6418 = 9'h107 == _GEN_15398 ? phv_data_263 : _GEN_6417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6419 = 9'h108 == _GEN_15398 ? phv_data_264 : _GEN_6418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6420 = 9'h109 == _GEN_15398 ? phv_data_265 : _GEN_6419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6421 = 9'h10a == _GEN_15398 ? phv_data_266 : _GEN_6420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6422 = 9'h10b == _GEN_15398 ? phv_data_267 : _GEN_6421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6423 = 9'h10c == _GEN_15398 ? phv_data_268 : _GEN_6422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6424 = 9'h10d == _GEN_15398 ? phv_data_269 : _GEN_6423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6425 = 9'h10e == _GEN_15398 ? phv_data_270 : _GEN_6424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6426 = 9'h10f == _GEN_15398 ? phv_data_271 : _GEN_6425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6427 = 9'h110 == _GEN_15398 ? phv_data_272 : _GEN_6426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6428 = 9'h111 == _GEN_15398 ? phv_data_273 : _GEN_6427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6429 = 9'h112 == _GEN_15398 ? phv_data_274 : _GEN_6428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6430 = 9'h113 == _GEN_15398 ? phv_data_275 : _GEN_6429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6431 = 9'h114 == _GEN_15398 ? phv_data_276 : _GEN_6430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6432 = 9'h115 == _GEN_15398 ? phv_data_277 : _GEN_6431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6433 = 9'h116 == _GEN_15398 ? phv_data_278 : _GEN_6432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6434 = 9'h117 == _GEN_15398 ? phv_data_279 : _GEN_6433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6435 = 9'h118 == _GEN_15398 ? phv_data_280 : _GEN_6434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6436 = 9'h119 == _GEN_15398 ? phv_data_281 : _GEN_6435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6437 = 9'h11a == _GEN_15398 ? phv_data_282 : _GEN_6436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6438 = 9'h11b == _GEN_15398 ? phv_data_283 : _GEN_6437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6439 = 9'h11c == _GEN_15398 ? phv_data_284 : _GEN_6438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6440 = 9'h11d == _GEN_15398 ? phv_data_285 : _GEN_6439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6441 = 9'h11e == _GEN_15398 ? phv_data_286 : _GEN_6440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6442 = 9'h11f == _GEN_15398 ? phv_data_287 : _GEN_6441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6443 = 9'h120 == _GEN_15398 ? phv_data_288 : _GEN_6442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6444 = 9'h121 == _GEN_15398 ? phv_data_289 : _GEN_6443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6445 = 9'h122 == _GEN_15398 ? phv_data_290 : _GEN_6444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6446 = 9'h123 == _GEN_15398 ? phv_data_291 : _GEN_6445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6447 = 9'h124 == _GEN_15398 ? phv_data_292 : _GEN_6446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6448 = 9'h125 == _GEN_15398 ? phv_data_293 : _GEN_6447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6449 = 9'h126 == _GEN_15398 ? phv_data_294 : _GEN_6448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6450 = 9'h127 == _GEN_15398 ? phv_data_295 : _GEN_6449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6451 = 9'h128 == _GEN_15398 ? phv_data_296 : _GEN_6450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6452 = 9'h129 == _GEN_15398 ? phv_data_297 : _GEN_6451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6453 = 9'h12a == _GEN_15398 ? phv_data_298 : _GEN_6452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6454 = 9'h12b == _GEN_15398 ? phv_data_299 : _GEN_6453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6455 = 9'h12c == _GEN_15398 ? phv_data_300 : _GEN_6454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6456 = 9'h12d == _GEN_15398 ? phv_data_301 : _GEN_6455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6457 = 9'h12e == _GEN_15398 ? phv_data_302 : _GEN_6456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6458 = 9'h12f == _GEN_15398 ? phv_data_303 : _GEN_6457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6459 = 9'h130 == _GEN_15398 ? phv_data_304 : _GEN_6458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6460 = 9'h131 == _GEN_15398 ? phv_data_305 : _GEN_6459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6461 = 9'h132 == _GEN_15398 ? phv_data_306 : _GEN_6460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6462 = 9'h133 == _GEN_15398 ? phv_data_307 : _GEN_6461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6463 = 9'h134 == _GEN_15398 ? phv_data_308 : _GEN_6462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6464 = 9'h135 == _GEN_15398 ? phv_data_309 : _GEN_6463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6465 = 9'h136 == _GEN_15398 ? phv_data_310 : _GEN_6464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6466 = 9'h137 == _GEN_15398 ? phv_data_311 : _GEN_6465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6467 = 9'h138 == _GEN_15398 ? phv_data_312 : _GEN_6466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6468 = 9'h139 == _GEN_15398 ? phv_data_313 : _GEN_6467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6469 = 9'h13a == _GEN_15398 ? phv_data_314 : _GEN_6468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6470 = 9'h13b == _GEN_15398 ? phv_data_315 : _GEN_6469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6471 = 9'h13c == _GEN_15398 ? phv_data_316 : _GEN_6470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6472 = 9'h13d == _GEN_15398 ? phv_data_317 : _GEN_6471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6473 = 9'h13e == _GEN_15398 ? phv_data_318 : _GEN_6472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6474 = 9'h13f == _GEN_15398 ? phv_data_319 : _GEN_6473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6475 = 9'h140 == _GEN_15398 ? phv_data_320 : _GEN_6474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6476 = 9'h141 == _GEN_15398 ? phv_data_321 : _GEN_6475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6477 = 9'h142 == _GEN_15398 ? phv_data_322 : _GEN_6476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6478 = 9'h143 == _GEN_15398 ? phv_data_323 : _GEN_6477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6479 = 9'h144 == _GEN_15398 ? phv_data_324 : _GEN_6478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6480 = 9'h145 == _GEN_15398 ? phv_data_325 : _GEN_6479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6481 = 9'h146 == _GEN_15398 ? phv_data_326 : _GEN_6480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6482 = 9'h147 == _GEN_15398 ? phv_data_327 : _GEN_6481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6483 = 9'h148 == _GEN_15398 ? phv_data_328 : _GEN_6482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6484 = 9'h149 == _GEN_15398 ? phv_data_329 : _GEN_6483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6485 = 9'h14a == _GEN_15398 ? phv_data_330 : _GEN_6484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6486 = 9'h14b == _GEN_15398 ? phv_data_331 : _GEN_6485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6487 = 9'h14c == _GEN_15398 ? phv_data_332 : _GEN_6486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6488 = 9'h14d == _GEN_15398 ? phv_data_333 : _GEN_6487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6489 = 9'h14e == _GEN_15398 ? phv_data_334 : _GEN_6488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6490 = 9'h14f == _GEN_15398 ? phv_data_335 : _GEN_6489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6491 = 9'h150 == _GEN_15398 ? phv_data_336 : _GEN_6490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6492 = 9'h151 == _GEN_15398 ? phv_data_337 : _GEN_6491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6493 = 9'h152 == _GEN_15398 ? phv_data_338 : _GEN_6492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6494 = 9'h153 == _GEN_15398 ? phv_data_339 : _GEN_6493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6495 = 9'h154 == _GEN_15398 ? phv_data_340 : _GEN_6494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6496 = 9'h155 == _GEN_15398 ? phv_data_341 : _GEN_6495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6497 = 9'h156 == _GEN_15398 ? phv_data_342 : _GEN_6496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6498 = 9'h157 == _GEN_15398 ? phv_data_343 : _GEN_6497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6499 = 9'h158 == _GEN_15398 ? phv_data_344 : _GEN_6498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6500 = 9'h159 == _GEN_15398 ? phv_data_345 : _GEN_6499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6501 = 9'h15a == _GEN_15398 ? phv_data_346 : _GEN_6500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6502 = 9'h15b == _GEN_15398 ? phv_data_347 : _GEN_6501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6503 = 9'h15c == _GEN_15398 ? phv_data_348 : _GEN_6502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6504 = 9'h15d == _GEN_15398 ? phv_data_349 : _GEN_6503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6505 = 9'h15e == _GEN_15398 ? phv_data_350 : _GEN_6504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6506 = 9'h15f == _GEN_15398 ? phv_data_351 : _GEN_6505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6507 = 9'h160 == _GEN_15398 ? phv_data_352 : _GEN_6506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6508 = 9'h161 == _GEN_15398 ? phv_data_353 : _GEN_6507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6509 = 9'h162 == _GEN_15398 ? phv_data_354 : _GEN_6508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6510 = 9'h163 == _GEN_15398 ? phv_data_355 : _GEN_6509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6511 = 9'h164 == _GEN_15398 ? phv_data_356 : _GEN_6510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6512 = 9'h165 == _GEN_15398 ? phv_data_357 : _GEN_6511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6513 = 9'h166 == _GEN_15398 ? phv_data_358 : _GEN_6512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6514 = 9'h167 == _GEN_15398 ? phv_data_359 : _GEN_6513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6515 = 9'h168 == _GEN_15398 ? phv_data_360 : _GEN_6514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6516 = 9'h169 == _GEN_15398 ? phv_data_361 : _GEN_6515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6517 = 9'h16a == _GEN_15398 ? phv_data_362 : _GEN_6516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6518 = 9'h16b == _GEN_15398 ? phv_data_363 : _GEN_6517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6519 = 9'h16c == _GEN_15398 ? phv_data_364 : _GEN_6518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6520 = 9'h16d == _GEN_15398 ? phv_data_365 : _GEN_6519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6521 = 9'h16e == _GEN_15398 ? phv_data_366 : _GEN_6520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6522 = 9'h16f == _GEN_15398 ? phv_data_367 : _GEN_6521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6523 = 9'h170 == _GEN_15398 ? phv_data_368 : _GEN_6522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6524 = 9'h171 == _GEN_15398 ? phv_data_369 : _GEN_6523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6525 = 9'h172 == _GEN_15398 ? phv_data_370 : _GEN_6524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6526 = 9'h173 == _GEN_15398 ? phv_data_371 : _GEN_6525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6527 = 9'h174 == _GEN_15398 ? phv_data_372 : _GEN_6526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6528 = 9'h175 == _GEN_15398 ? phv_data_373 : _GEN_6527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6529 = 9'h176 == _GEN_15398 ? phv_data_374 : _GEN_6528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6530 = 9'h177 == _GEN_15398 ? phv_data_375 : _GEN_6529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6531 = 9'h178 == _GEN_15398 ? phv_data_376 : _GEN_6530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6532 = 9'h179 == _GEN_15398 ? phv_data_377 : _GEN_6531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6533 = 9'h17a == _GEN_15398 ? phv_data_378 : _GEN_6532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6534 = 9'h17b == _GEN_15398 ? phv_data_379 : _GEN_6533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6535 = 9'h17c == _GEN_15398 ? phv_data_380 : _GEN_6534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6536 = 9'h17d == _GEN_15398 ? phv_data_381 : _GEN_6535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6537 = 9'h17e == _GEN_15398 ? phv_data_382 : _GEN_6536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6538 = 9'h17f == _GEN_15398 ? phv_data_383 : _GEN_6537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6539 = 9'h180 == _GEN_15398 ? phv_data_384 : _GEN_6538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6540 = 9'h181 == _GEN_15398 ? phv_data_385 : _GEN_6539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6541 = 9'h182 == _GEN_15398 ? phv_data_386 : _GEN_6540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6542 = 9'h183 == _GEN_15398 ? phv_data_387 : _GEN_6541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6543 = 9'h184 == _GEN_15398 ? phv_data_388 : _GEN_6542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6544 = 9'h185 == _GEN_15398 ? phv_data_389 : _GEN_6543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6545 = 9'h186 == _GEN_15398 ? phv_data_390 : _GEN_6544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6546 = 9'h187 == _GEN_15398 ? phv_data_391 : _GEN_6545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6547 = 9'h188 == _GEN_15398 ? phv_data_392 : _GEN_6546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6548 = 9'h189 == _GEN_15398 ? phv_data_393 : _GEN_6547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6549 = 9'h18a == _GEN_15398 ? phv_data_394 : _GEN_6548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6550 = 9'h18b == _GEN_15398 ? phv_data_395 : _GEN_6549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6551 = 9'h18c == _GEN_15398 ? phv_data_396 : _GEN_6550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6552 = 9'h18d == _GEN_15398 ? phv_data_397 : _GEN_6551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6553 = 9'h18e == _GEN_15398 ? phv_data_398 : _GEN_6552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6554 = 9'h18f == _GEN_15398 ? phv_data_399 : _GEN_6553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6555 = 9'h190 == _GEN_15398 ? phv_data_400 : _GEN_6554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6556 = 9'h191 == _GEN_15398 ? phv_data_401 : _GEN_6555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6557 = 9'h192 == _GEN_15398 ? phv_data_402 : _GEN_6556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6558 = 9'h193 == _GEN_15398 ? phv_data_403 : _GEN_6557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6559 = 9'h194 == _GEN_15398 ? phv_data_404 : _GEN_6558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6560 = 9'h195 == _GEN_15398 ? phv_data_405 : _GEN_6559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6561 = 9'h196 == _GEN_15398 ? phv_data_406 : _GEN_6560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6562 = 9'h197 == _GEN_15398 ? phv_data_407 : _GEN_6561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6563 = 9'h198 == _GEN_15398 ? phv_data_408 : _GEN_6562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6564 = 9'h199 == _GEN_15398 ? phv_data_409 : _GEN_6563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6565 = 9'h19a == _GEN_15398 ? phv_data_410 : _GEN_6564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6566 = 9'h19b == _GEN_15398 ? phv_data_411 : _GEN_6565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6567 = 9'h19c == _GEN_15398 ? phv_data_412 : _GEN_6566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6568 = 9'h19d == _GEN_15398 ? phv_data_413 : _GEN_6567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6569 = 9'h19e == _GEN_15398 ? phv_data_414 : _GEN_6568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6570 = 9'h19f == _GEN_15398 ? phv_data_415 : _GEN_6569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6571 = 9'h1a0 == _GEN_15398 ? phv_data_416 : _GEN_6570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6572 = 9'h1a1 == _GEN_15398 ? phv_data_417 : _GEN_6571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6573 = 9'h1a2 == _GEN_15398 ? phv_data_418 : _GEN_6572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6574 = 9'h1a3 == _GEN_15398 ? phv_data_419 : _GEN_6573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6575 = 9'h1a4 == _GEN_15398 ? phv_data_420 : _GEN_6574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6576 = 9'h1a5 == _GEN_15398 ? phv_data_421 : _GEN_6575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6577 = 9'h1a6 == _GEN_15398 ? phv_data_422 : _GEN_6576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6578 = 9'h1a7 == _GEN_15398 ? phv_data_423 : _GEN_6577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6579 = 9'h1a8 == _GEN_15398 ? phv_data_424 : _GEN_6578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6580 = 9'h1a9 == _GEN_15398 ? phv_data_425 : _GEN_6579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6581 = 9'h1aa == _GEN_15398 ? phv_data_426 : _GEN_6580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6582 = 9'h1ab == _GEN_15398 ? phv_data_427 : _GEN_6581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6583 = 9'h1ac == _GEN_15398 ? phv_data_428 : _GEN_6582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6584 = 9'h1ad == _GEN_15398 ? phv_data_429 : _GEN_6583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6585 = 9'h1ae == _GEN_15398 ? phv_data_430 : _GEN_6584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6586 = 9'h1af == _GEN_15398 ? phv_data_431 : _GEN_6585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6587 = 9'h1b0 == _GEN_15398 ? phv_data_432 : _GEN_6586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6588 = 9'h1b1 == _GEN_15398 ? phv_data_433 : _GEN_6587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6589 = 9'h1b2 == _GEN_15398 ? phv_data_434 : _GEN_6588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6590 = 9'h1b3 == _GEN_15398 ? phv_data_435 : _GEN_6589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6591 = 9'h1b4 == _GEN_15398 ? phv_data_436 : _GEN_6590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6592 = 9'h1b5 == _GEN_15398 ? phv_data_437 : _GEN_6591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6593 = 9'h1b6 == _GEN_15398 ? phv_data_438 : _GEN_6592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6594 = 9'h1b7 == _GEN_15398 ? phv_data_439 : _GEN_6593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6595 = 9'h1b8 == _GEN_15398 ? phv_data_440 : _GEN_6594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6596 = 9'h1b9 == _GEN_15398 ? phv_data_441 : _GEN_6595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6597 = 9'h1ba == _GEN_15398 ? phv_data_442 : _GEN_6596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6598 = 9'h1bb == _GEN_15398 ? phv_data_443 : _GEN_6597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6599 = 9'h1bc == _GEN_15398 ? phv_data_444 : _GEN_6598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6600 = 9'h1bd == _GEN_15398 ? phv_data_445 : _GEN_6599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6601 = 9'h1be == _GEN_15398 ? phv_data_446 : _GEN_6600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6602 = 9'h1bf == _GEN_15398 ? phv_data_447 : _GEN_6601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6603 = 9'h1c0 == _GEN_15398 ? phv_data_448 : _GEN_6602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6604 = 9'h1c1 == _GEN_15398 ? phv_data_449 : _GEN_6603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6605 = 9'h1c2 == _GEN_15398 ? phv_data_450 : _GEN_6604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6606 = 9'h1c3 == _GEN_15398 ? phv_data_451 : _GEN_6605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6607 = 9'h1c4 == _GEN_15398 ? phv_data_452 : _GEN_6606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6608 = 9'h1c5 == _GEN_15398 ? phv_data_453 : _GEN_6607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6609 = 9'h1c6 == _GEN_15398 ? phv_data_454 : _GEN_6608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6610 = 9'h1c7 == _GEN_15398 ? phv_data_455 : _GEN_6609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6611 = 9'h1c8 == _GEN_15398 ? phv_data_456 : _GEN_6610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6612 = 9'h1c9 == _GEN_15398 ? phv_data_457 : _GEN_6611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6613 = 9'h1ca == _GEN_15398 ? phv_data_458 : _GEN_6612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6614 = 9'h1cb == _GEN_15398 ? phv_data_459 : _GEN_6613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6615 = 9'h1cc == _GEN_15398 ? phv_data_460 : _GEN_6614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6616 = 9'h1cd == _GEN_15398 ? phv_data_461 : _GEN_6615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6617 = 9'h1ce == _GEN_15398 ? phv_data_462 : _GEN_6616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6618 = 9'h1cf == _GEN_15398 ? phv_data_463 : _GEN_6617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6619 = 9'h1d0 == _GEN_15398 ? phv_data_464 : _GEN_6618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6620 = 9'h1d1 == _GEN_15398 ? phv_data_465 : _GEN_6619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6621 = 9'h1d2 == _GEN_15398 ? phv_data_466 : _GEN_6620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6622 = 9'h1d3 == _GEN_15398 ? phv_data_467 : _GEN_6621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6623 = 9'h1d4 == _GEN_15398 ? phv_data_468 : _GEN_6622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6624 = 9'h1d5 == _GEN_15398 ? phv_data_469 : _GEN_6623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6625 = 9'h1d6 == _GEN_15398 ? phv_data_470 : _GEN_6624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6626 = 9'h1d7 == _GEN_15398 ? phv_data_471 : _GEN_6625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6627 = 9'h1d8 == _GEN_15398 ? phv_data_472 : _GEN_6626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6628 = 9'h1d9 == _GEN_15398 ? phv_data_473 : _GEN_6627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6629 = 9'h1da == _GEN_15398 ? phv_data_474 : _GEN_6628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6630 = 9'h1db == _GEN_15398 ? phv_data_475 : _GEN_6629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6631 = 9'h1dc == _GEN_15398 ? phv_data_476 : _GEN_6630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6632 = 9'h1dd == _GEN_15398 ? phv_data_477 : _GEN_6631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6633 = 9'h1de == _GEN_15398 ? phv_data_478 : _GEN_6632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6634 = 9'h1df == _GEN_15398 ? phv_data_479 : _GEN_6633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6635 = 9'h1e0 == _GEN_15398 ? phv_data_480 : _GEN_6634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6636 = 9'h1e1 == _GEN_15398 ? phv_data_481 : _GEN_6635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6637 = 9'h1e2 == _GEN_15398 ? phv_data_482 : _GEN_6636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6638 = 9'h1e3 == _GEN_15398 ? phv_data_483 : _GEN_6637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6639 = 9'h1e4 == _GEN_15398 ? phv_data_484 : _GEN_6638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6640 = 9'h1e5 == _GEN_15398 ? phv_data_485 : _GEN_6639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6641 = 9'h1e6 == _GEN_15398 ? phv_data_486 : _GEN_6640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6642 = 9'h1e7 == _GEN_15398 ? phv_data_487 : _GEN_6641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6643 = 9'h1e8 == _GEN_15398 ? phv_data_488 : _GEN_6642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6644 = 9'h1e9 == _GEN_15398 ? phv_data_489 : _GEN_6643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6645 = 9'h1ea == _GEN_15398 ? phv_data_490 : _GEN_6644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6646 = 9'h1eb == _GEN_15398 ? phv_data_491 : _GEN_6645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6647 = 9'h1ec == _GEN_15398 ? phv_data_492 : _GEN_6646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6648 = 9'h1ed == _GEN_15398 ? phv_data_493 : _GEN_6647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6649 = 9'h1ee == _GEN_15398 ? phv_data_494 : _GEN_6648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6650 = 9'h1ef == _GEN_15398 ? phv_data_495 : _GEN_6649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6651 = 9'h1f0 == _GEN_15398 ? phv_data_496 : _GEN_6650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6652 = 9'h1f1 == _GEN_15398 ? phv_data_497 : _GEN_6651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6653 = 9'h1f2 == _GEN_15398 ? phv_data_498 : _GEN_6652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6654 = 9'h1f3 == _GEN_15398 ? phv_data_499 : _GEN_6653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6655 = 9'h1f4 == _GEN_15398 ? phv_data_500 : _GEN_6654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6656 = 9'h1f5 == _GEN_15398 ? phv_data_501 : _GEN_6655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6657 = 9'h1f6 == _GEN_15398 ? phv_data_502 : _GEN_6656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6658 = 9'h1f7 == _GEN_15398 ? phv_data_503 : _GEN_6657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6659 = 9'h1f8 == _GEN_15398 ? phv_data_504 : _GEN_6658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6660 = 9'h1f9 == _GEN_15398 ? phv_data_505 : _GEN_6659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6661 = 9'h1fa == _GEN_15398 ? phv_data_506 : _GEN_6660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6662 = 9'h1fb == _GEN_15398 ? phv_data_507 : _GEN_6661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6663 = 9'h1fc == _GEN_15398 ? phv_data_508 : _GEN_6662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6664 = 9'h1fd == _GEN_15398 ? phv_data_509 : _GEN_6663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6665 = 9'h1fe == _GEN_15398 ? phv_data_510 : _GEN_6664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6666 = 9'h1ff == _GEN_15398 ? phv_data_511 : _GEN_6665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6668 = 8'h1 == local_offset_3 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6669 = 8'h2 == local_offset_3 ? phv_data_2 : _GEN_6668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6670 = 8'h3 == local_offset_3 ? phv_data_3 : _GEN_6669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6671 = 8'h4 == local_offset_3 ? phv_data_4 : _GEN_6670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6672 = 8'h5 == local_offset_3 ? phv_data_5 : _GEN_6671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6673 = 8'h6 == local_offset_3 ? phv_data_6 : _GEN_6672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6674 = 8'h7 == local_offset_3 ? phv_data_7 : _GEN_6673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6675 = 8'h8 == local_offset_3 ? phv_data_8 : _GEN_6674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6676 = 8'h9 == local_offset_3 ? phv_data_9 : _GEN_6675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6677 = 8'ha == local_offset_3 ? phv_data_10 : _GEN_6676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6678 = 8'hb == local_offset_3 ? phv_data_11 : _GEN_6677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6679 = 8'hc == local_offset_3 ? phv_data_12 : _GEN_6678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6680 = 8'hd == local_offset_3 ? phv_data_13 : _GEN_6679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6681 = 8'he == local_offset_3 ? phv_data_14 : _GEN_6680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6682 = 8'hf == local_offset_3 ? phv_data_15 : _GEN_6681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6683 = 8'h10 == local_offset_3 ? phv_data_16 : _GEN_6682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6684 = 8'h11 == local_offset_3 ? phv_data_17 : _GEN_6683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6685 = 8'h12 == local_offset_3 ? phv_data_18 : _GEN_6684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6686 = 8'h13 == local_offset_3 ? phv_data_19 : _GEN_6685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6687 = 8'h14 == local_offset_3 ? phv_data_20 : _GEN_6686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6688 = 8'h15 == local_offset_3 ? phv_data_21 : _GEN_6687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6689 = 8'h16 == local_offset_3 ? phv_data_22 : _GEN_6688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6690 = 8'h17 == local_offset_3 ? phv_data_23 : _GEN_6689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6691 = 8'h18 == local_offset_3 ? phv_data_24 : _GEN_6690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6692 = 8'h19 == local_offset_3 ? phv_data_25 : _GEN_6691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6693 = 8'h1a == local_offset_3 ? phv_data_26 : _GEN_6692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6694 = 8'h1b == local_offset_3 ? phv_data_27 : _GEN_6693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6695 = 8'h1c == local_offset_3 ? phv_data_28 : _GEN_6694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6696 = 8'h1d == local_offset_3 ? phv_data_29 : _GEN_6695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6697 = 8'h1e == local_offset_3 ? phv_data_30 : _GEN_6696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6698 = 8'h1f == local_offset_3 ? phv_data_31 : _GEN_6697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6699 = 8'h20 == local_offset_3 ? phv_data_32 : _GEN_6698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6700 = 8'h21 == local_offset_3 ? phv_data_33 : _GEN_6699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6701 = 8'h22 == local_offset_3 ? phv_data_34 : _GEN_6700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6702 = 8'h23 == local_offset_3 ? phv_data_35 : _GEN_6701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6703 = 8'h24 == local_offset_3 ? phv_data_36 : _GEN_6702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6704 = 8'h25 == local_offset_3 ? phv_data_37 : _GEN_6703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6705 = 8'h26 == local_offset_3 ? phv_data_38 : _GEN_6704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6706 = 8'h27 == local_offset_3 ? phv_data_39 : _GEN_6705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6707 = 8'h28 == local_offset_3 ? phv_data_40 : _GEN_6706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6708 = 8'h29 == local_offset_3 ? phv_data_41 : _GEN_6707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6709 = 8'h2a == local_offset_3 ? phv_data_42 : _GEN_6708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6710 = 8'h2b == local_offset_3 ? phv_data_43 : _GEN_6709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6711 = 8'h2c == local_offset_3 ? phv_data_44 : _GEN_6710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6712 = 8'h2d == local_offset_3 ? phv_data_45 : _GEN_6711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6713 = 8'h2e == local_offset_3 ? phv_data_46 : _GEN_6712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6714 = 8'h2f == local_offset_3 ? phv_data_47 : _GEN_6713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6715 = 8'h30 == local_offset_3 ? phv_data_48 : _GEN_6714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6716 = 8'h31 == local_offset_3 ? phv_data_49 : _GEN_6715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6717 = 8'h32 == local_offset_3 ? phv_data_50 : _GEN_6716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6718 = 8'h33 == local_offset_3 ? phv_data_51 : _GEN_6717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6719 = 8'h34 == local_offset_3 ? phv_data_52 : _GEN_6718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6720 = 8'h35 == local_offset_3 ? phv_data_53 : _GEN_6719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6721 = 8'h36 == local_offset_3 ? phv_data_54 : _GEN_6720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6722 = 8'h37 == local_offset_3 ? phv_data_55 : _GEN_6721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6723 = 8'h38 == local_offset_3 ? phv_data_56 : _GEN_6722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6724 = 8'h39 == local_offset_3 ? phv_data_57 : _GEN_6723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6725 = 8'h3a == local_offset_3 ? phv_data_58 : _GEN_6724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6726 = 8'h3b == local_offset_3 ? phv_data_59 : _GEN_6725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6727 = 8'h3c == local_offset_3 ? phv_data_60 : _GEN_6726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6728 = 8'h3d == local_offset_3 ? phv_data_61 : _GEN_6727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6729 = 8'h3e == local_offset_3 ? phv_data_62 : _GEN_6728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6730 = 8'h3f == local_offset_3 ? phv_data_63 : _GEN_6729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6731 = 8'h40 == local_offset_3 ? phv_data_64 : _GEN_6730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6732 = 8'h41 == local_offset_3 ? phv_data_65 : _GEN_6731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6733 = 8'h42 == local_offset_3 ? phv_data_66 : _GEN_6732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6734 = 8'h43 == local_offset_3 ? phv_data_67 : _GEN_6733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6735 = 8'h44 == local_offset_3 ? phv_data_68 : _GEN_6734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6736 = 8'h45 == local_offset_3 ? phv_data_69 : _GEN_6735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6737 = 8'h46 == local_offset_3 ? phv_data_70 : _GEN_6736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6738 = 8'h47 == local_offset_3 ? phv_data_71 : _GEN_6737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6739 = 8'h48 == local_offset_3 ? phv_data_72 : _GEN_6738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6740 = 8'h49 == local_offset_3 ? phv_data_73 : _GEN_6739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6741 = 8'h4a == local_offset_3 ? phv_data_74 : _GEN_6740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6742 = 8'h4b == local_offset_3 ? phv_data_75 : _GEN_6741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6743 = 8'h4c == local_offset_3 ? phv_data_76 : _GEN_6742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6744 = 8'h4d == local_offset_3 ? phv_data_77 : _GEN_6743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6745 = 8'h4e == local_offset_3 ? phv_data_78 : _GEN_6744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6746 = 8'h4f == local_offset_3 ? phv_data_79 : _GEN_6745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6747 = 8'h50 == local_offset_3 ? phv_data_80 : _GEN_6746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6748 = 8'h51 == local_offset_3 ? phv_data_81 : _GEN_6747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6749 = 8'h52 == local_offset_3 ? phv_data_82 : _GEN_6748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6750 = 8'h53 == local_offset_3 ? phv_data_83 : _GEN_6749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6751 = 8'h54 == local_offset_3 ? phv_data_84 : _GEN_6750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6752 = 8'h55 == local_offset_3 ? phv_data_85 : _GEN_6751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6753 = 8'h56 == local_offset_3 ? phv_data_86 : _GEN_6752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6754 = 8'h57 == local_offset_3 ? phv_data_87 : _GEN_6753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6755 = 8'h58 == local_offset_3 ? phv_data_88 : _GEN_6754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6756 = 8'h59 == local_offset_3 ? phv_data_89 : _GEN_6755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6757 = 8'h5a == local_offset_3 ? phv_data_90 : _GEN_6756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6758 = 8'h5b == local_offset_3 ? phv_data_91 : _GEN_6757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6759 = 8'h5c == local_offset_3 ? phv_data_92 : _GEN_6758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6760 = 8'h5d == local_offset_3 ? phv_data_93 : _GEN_6759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6761 = 8'h5e == local_offset_3 ? phv_data_94 : _GEN_6760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6762 = 8'h5f == local_offset_3 ? phv_data_95 : _GEN_6761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6763 = 8'h60 == local_offset_3 ? phv_data_96 : _GEN_6762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6764 = 8'h61 == local_offset_3 ? phv_data_97 : _GEN_6763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6765 = 8'h62 == local_offset_3 ? phv_data_98 : _GEN_6764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6766 = 8'h63 == local_offset_3 ? phv_data_99 : _GEN_6765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6767 = 8'h64 == local_offset_3 ? phv_data_100 : _GEN_6766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6768 = 8'h65 == local_offset_3 ? phv_data_101 : _GEN_6767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6769 = 8'h66 == local_offset_3 ? phv_data_102 : _GEN_6768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6770 = 8'h67 == local_offset_3 ? phv_data_103 : _GEN_6769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6771 = 8'h68 == local_offset_3 ? phv_data_104 : _GEN_6770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6772 = 8'h69 == local_offset_3 ? phv_data_105 : _GEN_6771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6773 = 8'h6a == local_offset_3 ? phv_data_106 : _GEN_6772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6774 = 8'h6b == local_offset_3 ? phv_data_107 : _GEN_6773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6775 = 8'h6c == local_offset_3 ? phv_data_108 : _GEN_6774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6776 = 8'h6d == local_offset_3 ? phv_data_109 : _GEN_6775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6777 = 8'h6e == local_offset_3 ? phv_data_110 : _GEN_6776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6778 = 8'h6f == local_offset_3 ? phv_data_111 : _GEN_6777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6779 = 8'h70 == local_offset_3 ? phv_data_112 : _GEN_6778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6780 = 8'h71 == local_offset_3 ? phv_data_113 : _GEN_6779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6781 = 8'h72 == local_offset_3 ? phv_data_114 : _GEN_6780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6782 = 8'h73 == local_offset_3 ? phv_data_115 : _GEN_6781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6783 = 8'h74 == local_offset_3 ? phv_data_116 : _GEN_6782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6784 = 8'h75 == local_offset_3 ? phv_data_117 : _GEN_6783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6785 = 8'h76 == local_offset_3 ? phv_data_118 : _GEN_6784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6786 = 8'h77 == local_offset_3 ? phv_data_119 : _GEN_6785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6787 = 8'h78 == local_offset_3 ? phv_data_120 : _GEN_6786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6788 = 8'h79 == local_offset_3 ? phv_data_121 : _GEN_6787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6789 = 8'h7a == local_offset_3 ? phv_data_122 : _GEN_6788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6790 = 8'h7b == local_offset_3 ? phv_data_123 : _GEN_6789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6791 = 8'h7c == local_offset_3 ? phv_data_124 : _GEN_6790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6792 = 8'h7d == local_offset_3 ? phv_data_125 : _GEN_6791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6793 = 8'h7e == local_offset_3 ? phv_data_126 : _GEN_6792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6794 = 8'h7f == local_offset_3 ? phv_data_127 : _GEN_6793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6795 = 8'h80 == local_offset_3 ? phv_data_128 : _GEN_6794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6796 = 8'h81 == local_offset_3 ? phv_data_129 : _GEN_6795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6797 = 8'h82 == local_offset_3 ? phv_data_130 : _GEN_6796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6798 = 8'h83 == local_offset_3 ? phv_data_131 : _GEN_6797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6799 = 8'h84 == local_offset_3 ? phv_data_132 : _GEN_6798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6800 = 8'h85 == local_offset_3 ? phv_data_133 : _GEN_6799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6801 = 8'h86 == local_offset_3 ? phv_data_134 : _GEN_6800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6802 = 8'h87 == local_offset_3 ? phv_data_135 : _GEN_6801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6803 = 8'h88 == local_offset_3 ? phv_data_136 : _GEN_6802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6804 = 8'h89 == local_offset_3 ? phv_data_137 : _GEN_6803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6805 = 8'h8a == local_offset_3 ? phv_data_138 : _GEN_6804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6806 = 8'h8b == local_offset_3 ? phv_data_139 : _GEN_6805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6807 = 8'h8c == local_offset_3 ? phv_data_140 : _GEN_6806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6808 = 8'h8d == local_offset_3 ? phv_data_141 : _GEN_6807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6809 = 8'h8e == local_offset_3 ? phv_data_142 : _GEN_6808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6810 = 8'h8f == local_offset_3 ? phv_data_143 : _GEN_6809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6811 = 8'h90 == local_offset_3 ? phv_data_144 : _GEN_6810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6812 = 8'h91 == local_offset_3 ? phv_data_145 : _GEN_6811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6813 = 8'h92 == local_offset_3 ? phv_data_146 : _GEN_6812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6814 = 8'h93 == local_offset_3 ? phv_data_147 : _GEN_6813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6815 = 8'h94 == local_offset_3 ? phv_data_148 : _GEN_6814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6816 = 8'h95 == local_offset_3 ? phv_data_149 : _GEN_6815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6817 = 8'h96 == local_offset_3 ? phv_data_150 : _GEN_6816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6818 = 8'h97 == local_offset_3 ? phv_data_151 : _GEN_6817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6819 = 8'h98 == local_offset_3 ? phv_data_152 : _GEN_6818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6820 = 8'h99 == local_offset_3 ? phv_data_153 : _GEN_6819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6821 = 8'h9a == local_offset_3 ? phv_data_154 : _GEN_6820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6822 = 8'h9b == local_offset_3 ? phv_data_155 : _GEN_6821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6823 = 8'h9c == local_offset_3 ? phv_data_156 : _GEN_6822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6824 = 8'h9d == local_offset_3 ? phv_data_157 : _GEN_6823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6825 = 8'h9e == local_offset_3 ? phv_data_158 : _GEN_6824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6826 = 8'h9f == local_offset_3 ? phv_data_159 : _GEN_6825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6827 = 8'ha0 == local_offset_3 ? phv_data_160 : _GEN_6826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6828 = 8'ha1 == local_offset_3 ? phv_data_161 : _GEN_6827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6829 = 8'ha2 == local_offset_3 ? phv_data_162 : _GEN_6828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6830 = 8'ha3 == local_offset_3 ? phv_data_163 : _GEN_6829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6831 = 8'ha4 == local_offset_3 ? phv_data_164 : _GEN_6830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6832 = 8'ha5 == local_offset_3 ? phv_data_165 : _GEN_6831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6833 = 8'ha6 == local_offset_3 ? phv_data_166 : _GEN_6832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6834 = 8'ha7 == local_offset_3 ? phv_data_167 : _GEN_6833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6835 = 8'ha8 == local_offset_3 ? phv_data_168 : _GEN_6834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6836 = 8'ha9 == local_offset_3 ? phv_data_169 : _GEN_6835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6837 = 8'haa == local_offset_3 ? phv_data_170 : _GEN_6836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6838 = 8'hab == local_offset_3 ? phv_data_171 : _GEN_6837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6839 = 8'hac == local_offset_3 ? phv_data_172 : _GEN_6838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6840 = 8'had == local_offset_3 ? phv_data_173 : _GEN_6839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6841 = 8'hae == local_offset_3 ? phv_data_174 : _GEN_6840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6842 = 8'haf == local_offset_3 ? phv_data_175 : _GEN_6841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6843 = 8'hb0 == local_offset_3 ? phv_data_176 : _GEN_6842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6844 = 8'hb1 == local_offset_3 ? phv_data_177 : _GEN_6843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6845 = 8'hb2 == local_offset_3 ? phv_data_178 : _GEN_6844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6846 = 8'hb3 == local_offset_3 ? phv_data_179 : _GEN_6845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6847 = 8'hb4 == local_offset_3 ? phv_data_180 : _GEN_6846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6848 = 8'hb5 == local_offset_3 ? phv_data_181 : _GEN_6847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6849 = 8'hb6 == local_offset_3 ? phv_data_182 : _GEN_6848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6850 = 8'hb7 == local_offset_3 ? phv_data_183 : _GEN_6849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6851 = 8'hb8 == local_offset_3 ? phv_data_184 : _GEN_6850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6852 = 8'hb9 == local_offset_3 ? phv_data_185 : _GEN_6851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6853 = 8'hba == local_offset_3 ? phv_data_186 : _GEN_6852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6854 = 8'hbb == local_offset_3 ? phv_data_187 : _GEN_6853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6855 = 8'hbc == local_offset_3 ? phv_data_188 : _GEN_6854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6856 = 8'hbd == local_offset_3 ? phv_data_189 : _GEN_6855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6857 = 8'hbe == local_offset_3 ? phv_data_190 : _GEN_6856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6858 = 8'hbf == local_offset_3 ? phv_data_191 : _GEN_6857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6859 = 8'hc0 == local_offset_3 ? phv_data_192 : _GEN_6858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6860 = 8'hc1 == local_offset_3 ? phv_data_193 : _GEN_6859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6861 = 8'hc2 == local_offset_3 ? phv_data_194 : _GEN_6860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6862 = 8'hc3 == local_offset_3 ? phv_data_195 : _GEN_6861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6863 = 8'hc4 == local_offset_3 ? phv_data_196 : _GEN_6862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6864 = 8'hc5 == local_offset_3 ? phv_data_197 : _GEN_6863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6865 = 8'hc6 == local_offset_3 ? phv_data_198 : _GEN_6864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6866 = 8'hc7 == local_offset_3 ? phv_data_199 : _GEN_6865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6867 = 8'hc8 == local_offset_3 ? phv_data_200 : _GEN_6866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6868 = 8'hc9 == local_offset_3 ? phv_data_201 : _GEN_6867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6869 = 8'hca == local_offset_3 ? phv_data_202 : _GEN_6868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6870 = 8'hcb == local_offset_3 ? phv_data_203 : _GEN_6869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6871 = 8'hcc == local_offset_3 ? phv_data_204 : _GEN_6870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6872 = 8'hcd == local_offset_3 ? phv_data_205 : _GEN_6871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6873 = 8'hce == local_offset_3 ? phv_data_206 : _GEN_6872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6874 = 8'hcf == local_offset_3 ? phv_data_207 : _GEN_6873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6875 = 8'hd0 == local_offset_3 ? phv_data_208 : _GEN_6874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6876 = 8'hd1 == local_offset_3 ? phv_data_209 : _GEN_6875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6877 = 8'hd2 == local_offset_3 ? phv_data_210 : _GEN_6876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6878 = 8'hd3 == local_offset_3 ? phv_data_211 : _GEN_6877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6879 = 8'hd4 == local_offset_3 ? phv_data_212 : _GEN_6878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6880 = 8'hd5 == local_offset_3 ? phv_data_213 : _GEN_6879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6881 = 8'hd6 == local_offset_3 ? phv_data_214 : _GEN_6880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6882 = 8'hd7 == local_offset_3 ? phv_data_215 : _GEN_6881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6883 = 8'hd8 == local_offset_3 ? phv_data_216 : _GEN_6882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6884 = 8'hd9 == local_offset_3 ? phv_data_217 : _GEN_6883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6885 = 8'hda == local_offset_3 ? phv_data_218 : _GEN_6884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6886 = 8'hdb == local_offset_3 ? phv_data_219 : _GEN_6885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6887 = 8'hdc == local_offset_3 ? phv_data_220 : _GEN_6886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6888 = 8'hdd == local_offset_3 ? phv_data_221 : _GEN_6887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6889 = 8'hde == local_offset_3 ? phv_data_222 : _GEN_6888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6890 = 8'hdf == local_offset_3 ? phv_data_223 : _GEN_6889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6891 = 8'he0 == local_offset_3 ? phv_data_224 : _GEN_6890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6892 = 8'he1 == local_offset_3 ? phv_data_225 : _GEN_6891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6893 = 8'he2 == local_offset_3 ? phv_data_226 : _GEN_6892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6894 = 8'he3 == local_offset_3 ? phv_data_227 : _GEN_6893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6895 = 8'he4 == local_offset_3 ? phv_data_228 : _GEN_6894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6896 = 8'he5 == local_offset_3 ? phv_data_229 : _GEN_6895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6897 = 8'he6 == local_offset_3 ? phv_data_230 : _GEN_6896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6898 = 8'he7 == local_offset_3 ? phv_data_231 : _GEN_6897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6899 = 8'he8 == local_offset_3 ? phv_data_232 : _GEN_6898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6900 = 8'he9 == local_offset_3 ? phv_data_233 : _GEN_6899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6901 = 8'hea == local_offset_3 ? phv_data_234 : _GEN_6900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6902 = 8'heb == local_offset_3 ? phv_data_235 : _GEN_6901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6903 = 8'hec == local_offset_3 ? phv_data_236 : _GEN_6902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6904 = 8'hed == local_offset_3 ? phv_data_237 : _GEN_6903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6905 = 8'hee == local_offset_3 ? phv_data_238 : _GEN_6904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6906 = 8'hef == local_offset_3 ? phv_data_239 : _GEN_6905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6907 = 8'hf0 == local_offset_3 ? phv_data_240 : _GEN_6906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6908 = 8'hf1 == local_offset_3 ? phv_data_241 : _GEN_6907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6909 = 8'hf2 == local_offset_3 ? phv_data_242 : _GEN_6908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6910 = 8'hf3 == local_offset_3 ? phv_data_243 : _GEN_6909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6911 = 8'hf4 == local_offset_3 ? phv_data_244 : _GEN_6910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6912 = 8'hf5 == local_offset_3 ? phv_data_245 : _GEN_6911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6913 = 8'hf6 == local_offset_3 ? phv_data_246 : _GEN_6912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6914 = 8'hf7 == local_offset_3 ? phv_data_247 : _GEN_6913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6915 = 8'hf8 == local_offset_3 ? phv_data_248 : _GEN_6914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6916 = 8'hf9 == local_offset_3 ? phv_data_249 : _GEN_6915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6917 = 8'hfa == local_offset_3 ? phv_data_250 : _GEN_6916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6918 = 8'hfb == local_offset_3 ? phv_data_251 : _GEN_6917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6919 = 8'hfc == local_offset_3 ? phv_data_252 : _GEN_6918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6920 = 8'hfd == local_offset_3 ? phv_data_253 : _GEN_6919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6921 = 8'hfe == local_offset_3 ? phv_data_254 : _GEN_6920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6922 = 8'hff == local_offset_3 ? phv_data_255 : _GEN_6921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_15654 = {{1'd0}, local_offset_3}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6923 = 9'h100 == _GEN_15654 ? phv_data_256 : _GEN_6922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6924 = 9'h101 == _GEN_15654 ? phv_data_257 : _GEN_6923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6925 = 9'h102 == _GEN_15654 ? phv_data_258 : _GEN_6924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6926 = 9'h103 == _GEN_15654 ? phv_data_259 : _GEN_6925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6927 = 9'h104 == _GEN_15654 ? phv_data_260 : _GEN_6926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6928 = 9'h105 == _GEN_15654 ? phv_data_261 : _GEN_6927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6929 = 9'h106 == _GEN_15654 ? phv_data_262 : _GEN_6928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6930 = 9'h107 == _GEN_15654 ? phv_data_263 : _GEN_6929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6931 = 9'h108 == _GEN_15654 ? phv_data_264 : _GEN_6930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6932 = 9'h109 == _GEN_15654 ? phv_data_265 : _GEN_6931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6933 = 9'h10a == _GEN_15654 ? phv_data_266 : _GEN_6932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6934 = 9'h10b == _GEN_15654 ? phv_data_267 : _GEN_6933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6935 = 9'h10c == _GEN_15654 ? phv_data_268 : _GEN_6934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6936 = 9'h10d == _GEN_15654 ? phv_data_269 : _GEN_6935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6937 = 9'h10e == _GEN_15654 ? phv_data_270 : _GEN_6936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6938 = 9'h10f == _GEN_15654 ? phv_data_271 : _GEN_6937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6939 = 9'h110 == _GEN_15654 ? phv_data_272 : _GEN_6938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6940 = 9'h111 == _GEN_15654 ? phv_data_273 : _GEN_6939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6941 = 9'h112 == _GEN_15654 ? phv_data_274 : _GEN_6940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6942 = 9'h113 == _GEN_15654 ? phv_data_275 : _GEN_6941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6943 = 9'h114 == _GEN_15654 ? phv_data_276 : _GEN_6942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6944 = 9'h115 == _GEN_15654 ? phv_data_277 : _GEN_6943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6945 = 9'h116 == _GEN_15654 ? phv_data_278 : _GEN_6944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6946 = 9'h117 == _GEN_15654 ? phv_data_279 : _GEN_6945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6947 = 9'h118 == _GEN_15654 ? phv_data_280 : _GEN_6946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6948 = 9'h119 == _GEN_15654 ? phv_data_281 : _GEN_6947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6949 = 9'h11a == _GEN_15654 ? phv_data_282 : _GEN_6948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6950 = 9'h11b == _GEN_15654 ? phv_data_283 : _GEN_6949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6951 = 9'h11c == _GEN_15654 ? phv_data_284 : _GEN_6950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6952 = 9'h11d == _GEN_15654 ? phv_data_285 : _GEN_6951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6953 = 9'h11e == _GEN_15654 ? phv_data_286 : _GEN_6952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6954 = 9'h11f == _GEN_15654 ? phv_data_287 : _GEN_6953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6955 = 9'h120 == _GEN_15654 ? phv_data_288 : _GEN_6954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6956 = 9'h121 == _GEN_15654 ? phv_data_289 : _GEN_6955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6957 = 9'h122 == _GEN_15654 ? phv_data_290 : _GEN_6956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6958 = 9'h123 == _GEN_15654 ? phv_data_291 : _GEN_6957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6959 = 9'h124 == _GEN_15654 ? phv_data_292 : _GEN_6958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6960 = 9'h125 == _GEN_15654 ? phv_data_293 : _GEN_6959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6961 = 9'h126 == _GEN_15654 ? phv_data_294 : _GEN_6960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6962 = 9'h127 == _GEN_15654 ? phv_data_295 : _GEN_6961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6963 = 9'h128 == _GEN_15654 ? phv_data_296 : _GEN_6962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6964 = 9'h129 == _GEN_15654 ? phv_data_297 : _GEN_6963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6965 = 9'h12a == _GEN_15654 ? phv_data_298 : _GEN_6964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6966 = 9'h12b == _GEN_15654 ? phv_data_299 : _GEN_6965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6967 = 9'h12c == _GEN_15654 ? phv_data_300 : _GEN_6966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6968 = 9'h12d == _GEN_15654 ? phv_data_301 : _GEN_6967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6969 = 9'h12e == _GEN_15654 ? phv_data_302 : _GEN_6968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6970 = 9'h12f == _GEN_15654 ? phv_data_303 : _GEN_6969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6971 = 9'h130 == _GEN_15654 ? phv_data_304 : _GEN_6970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6972 = 9'h131 == _GEN_15654 ? phv_data_305 : _GEN_6971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6973 = 9'h132 == _GEN_15654 ? phv_data_306 : _GEN_6972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6974 = 9'h133 == _GEN_15654 ? phv_data_307 : _GEN_6973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6975 = 9'h134 == _GEN_15654 ? phv_data_308 : _GEN_6974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6976 = 9'h135 == _GEN_15654 ? phv_data_309 : _GEN_6975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6977 = 9'h136 == _GEN_15654 ? phv_data_310 : _GEN_6976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6978 = 9'h137 == _GEN_15654 ? phv_data_311 : _GEN_6977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6979 = 9'h138 == _GEN_15654 ? phv_data_312 : _GEN_6978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6980 = 9'h139 == _GEN_15654 ? phv_data_313 : _GEN_6979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6981 = 9'h13a == _GEN_15654 ? phv_data_314 : _GEN_6980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6982 = 9'h13b == _GEN_15654 ? phv_data_315 : _GEN_6981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6983 = 9'h13c == _GEN_15654 ? phv_data_316 : _GEN_6982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6984 = 9'h13d == _GEN_15654 ? phv_data_317 : _GEN_6983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6985 = 9'h13e == _GEN_15654 ? phv_data_318 : _GEN_6984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6986 = 9'h13f == _GEN_15654 ? phv_data_319 : _GEN_6985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6987 = 9'h140 == _GEN_15654 ? phv_data_320 : _GEN_6986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6988 = 9'h141 == _GEN_15654 ? phv_data_321 : _GEN_6987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6989 = 9'h142 == _GEN_15654 ? phv_data_322 : _GEN_6988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6990 = 9'h143 == _GEN_15654 ? phv_data_323 : _GEN_6989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6991 = 9'h144 == _GEN_15654 ? phv_data_324 : _GEN_6990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6992 = 9'h145 == _GEN_15654 ? phv_data_325 : _GEN_6991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6993 = 9'h146 == _GEN_15654 ? phv_data_326 : _GEN_6992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6994 = 9'h147 == _GEN_15654 ? phv_data_327 : _GEN_6993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6995 = 9'h148 == _GEN_15654 ? phv_data_328 : _GEN_6994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6996 = 9'h149 == _GEN_15654 ? phv_data_329 : _GEN_6995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6997 = 9'h14a == _GEN_15654 ? phv_data_330 : _GEN_6996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6998 = 9'h14b == _GEN_15654 ? phv_data_331 : _GEN_6997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6999 = 9'h14c == _GEN_15654 ? phv_data_332 : _GEN_6998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7000 = 9'h14d == _GEN_15654 ? phv_data_333 : _GEN_6999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7001 = 9'h14e == _GEN_15654 ? phv_data_334 : _GEN_7000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7002 = 9'h14f == _GEN_15654 ? phv_data_335 : _GEN_7001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7003 = 9'h150 == _GEN_15654 ? phv_data_336 : _GEN_7002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7004 = 9'h151 == _GEN_15654 ? phv_data_337 : _GEN_7003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7005 = 9'h152 == _GEN_15654 ? phv_data_338 : _GEN_7004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7006 = 9'h153 == _GEN_15654 ? phv_data_339 : _GEN_7005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7007 = 9'h154 == _GEN_15654 ? phv_data_340 : _GEN_7006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7008 = 9'h155 == _GEN_15654 ? phv_data_341 : _GEN_7007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7009 = 9'h156 == _GEN_15654 ? phv_data_342 : _GEN_7008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7010 = 9'h157 == _GEN_15654 ? phv_data_343 : _GEN_7009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7011 = 9'h158 == _GEN_15654 ? phv_data_344 : _GEN_7010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7012 = 9'h159 == _GEN_15654 ? phv_data_345 : _GEN_7011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7013 = 9'h15a == _GEN_15654 ? phv_data_346 : _GEN_7012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7014 = 9'h15b == _GEN_15654 ? phv_data_347 : _GEN_7013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7015 = 9'h15c == _GEN_15654 ? phv_data_348 : _GEN_7014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7016 = 9'h15d == _GEN_15654 ? phv_data_349 : _GEN_7015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7017 = 9'h15e == _GEN_15654 ? phv_data_350 : _GEN_7016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7018 = 9'h15f == _GEN_15654 ? phv_data_351 : _GEN_7017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7019 = 9'h160 == _GEN_15654 ? phv_data_352 : _GEN_7018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7020 = 9'h161 == _GEN_15654 ? phv_data_353 : _GEN_7019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7021 = 9'h162 == _GEN_15654 ? phv_data_354 : _GEN_7020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7022 = 9'h163 == _GEN_15654 ? phv_data_355 : _GEN_7021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7023 = 9'h164 == _GEN_15654 ? phv_data_356 : _GEN_7022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7024 = 9'h165 == _GEN_15654 ? phv_data_357 : _GEN_7023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7025 = 9'h166 == _GEN_15654 ? phv_data_358 : _GEN_7024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7026 = 9'h167 == _GEN_15654 ? phv_data_359 : _GEN_7025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7027 = 9'h168 == _GEN_15654 ? phv_data_360 : _GEN_7026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7028 = 9'h169 == _GEN_15654 ? phv_data_361 : _GEN_7027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7029 = 9'h16a == _GEN_15654 ? phv_data_362 : _GEN_7028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7030 = 9'h16b == _GEN_15654 ? phv_data_363 : _GEN_7029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7031 = 9'h16c == _GEN_15654 ? phv_data_364 : _GEN_7030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7032 = 9'h16d == _GEN_15654 ? phv_data_365 : _GEN_7031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7033 = 9'h16e == _GEN_15654 ? phv_data_366 : _GEN_7032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7034 = 9'h16f == _GEN_15654 ? phv_data_367 : _GEN_7033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7035 = 9'h170 == _GEN_15654 ? phv_data_368 : _GEN_7034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7036 = 9'h171 == _GEN_15654 ? phv_data_369 : _GEN_7035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7037 = 9'h172 == _GEN_15654 ? phv_data_370 : _GEN_7036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7038 = 9'h173 == _GEN_15654 ? phv_data_371 : _GEN_7037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7039 = 9'h174 == _GEN_15654 ? phv_data_372 : _GEN_7038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7040 = 9'h175 == _GEN_15654 ? phv_data_373 : _GEN_7039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7041 = 9'h176 == _GEN_15654 ? phv_data_374 : _GEN_7040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7042 = 9'h177 == _GEN_15654 ? phv_data_375 : _GEN_7041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7043 = 9'h178 == _GEN_15654 ? phv_data_376 : _GEN_7042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7044 = 9'h179 == _GEN_15654 ? phv_data_377 : _GEN_7043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7045 = 9'h17a == _GEN_15654 ? phv_data_378 : _GEN_7044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7046 = 9'h17b == _GEN_15654 ? phv_data_379 : _GEN_7045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7047 = 9'h17c == _GEN_15654 ? phv_data_380 : _GEN_7046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7048 = 9'h17d == _GEN_15654 ? phv_data_381 : _GEN_7047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7049 = 9'h17e == _GEN_15654 ? phv_data_382 : _GEN_7048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7050 = 9'h17f == _GEN_15654 ? phv_data_383 : _GEN_7049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7051 = 9'h180 == _GEN_15654 ? phv_data_384 : _GEN_7050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7052 = 9'h181 == _GEN_15654 ? phv_data_385 : _GEN_7051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7053 = 9'h182 == _GEN_15654 ? phv_data_386 : _GEN_7052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7054 = 9'h183 == _GEN_15654 ? phv_data_387 : _GEN_7053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7055 = 9'h184 == _GEN_15654 ? phv_data_388 : _GEN_7054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7056 = 9'h185 == _GEN_15654 ? phv_data_389 : _GEN_7055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7057 = 9'h186 == _GEN_15654 ? phv_data_390 : _GEN_7056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7058 = 9'h187 == _GEN_15654 ? phv_data_391 : _GEN_7057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7059 = 9'h188 == _GEN_15654 ? phv_data_392 : _GEN_7058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7060 = 9'h189 == _GEN_15654 ? phv_data_393 : _GEN_7059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7061 = 9'h18a == _GEN_15654 ? phv_data_394 : _GEN_7060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7062 = 9'h18b == _GEN_15654 ? phv_data_395 : _GEN_7061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7063 = 9'h18c == _GEN_15654 ? phv_data_396 : _GEN_7062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7064 = 9'h18d == _GEN_15654 ? phv_data_397 : _GEN_7063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7065 = 9'h18e == _GEN_15654 ? phv_data_398 : _GEN_7064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7066 = 9'h18f == _GEN_15654 ? phv_data_399 : _GEN_7065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7067 = 9'h190 == _GEN_15654 ? phv_data_400 : _GEN_7066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7068 = 9'h191 == _GEN_15654 ? phv_data_401 : _GEN_7067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7069 = 9'h192 == _GEN_15654 ? phv_data_402 : _GEN_7068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7070 = 9'h193 == _GEN_15654 ? phv_data_403 : _GEN_7069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7071 = 9'h194 == _GEN_15654 ? phv_data_404 : _GEN_7070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7072 = 9'h195 == _GEN_15654 ? phv_data_405 : _GEN_7071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7073 = 9'h196 == _GEN_15654 ? phv_data_406 : _GEN_7072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7074 = 9'h197 == _GEN_15654 ? phv_data_407 : _GEN_7073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7075 = 9'h198 == _GEN_15654 ? phv_data_408 : _GEN_7074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7076 = 9'h199 == _GEN_15654 ? phv_data_409 : _GEN_7075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7077 = 9'h19a == _GEN_15654 ? phv_data_410 : _GEN_7076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7078 = 9'h19b == _GEN_15654 ? phv_data_411 : _GEN_7077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7079 = 9'h19c == _GEN_15654 ? phv_data_412 : _GEN_7078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7080 = 9'h19d == _GEN_15654 ? phv_data_413 : _GEN_7079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7081 = 9'h19e == _GEN_15654 ? phv_data_414 : _GEN_7080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7082 = 9'h19f == _GEN_15654 ? phv_data_415 : _GEN_7081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7083 = 9'h1a0 == _GEN_15654 ? phv_data_416 : _GEN_7082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7084 = 9'h1a1 == _GEN_15654 ? phv_data_417 : _GEN_7083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7085 = 9'h1a2 == _GEN_15654 ? phv_data_418 : _GEN_7084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7086 = 9'h1a3 == _GEN_15654 ? phv_data_419 : _GEN_7085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7087 = 9'h1a4 == _GEN_15654 ? phv_data_420 : _GEN_7086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7088 = 9'h1a5 == _GEN_15654 ? phv_data_421 : _GEN_7087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7089 = 9'h1a6 == _GEN_15654 ? phv_data_422 : _GEN_7088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7090 = 9'h1a7 == _GEN_15654 ? phv_data_423 : _GEN_7089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7091 = 9'h1a8 == _GEN_15654 ? phv_data_424 : _GEN_7090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7092 = 9'h1a9 == _GEN_15654 ? phv_data_425 : _GEN_7091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7093 = 9'h1aa == _GEN_15654 ? phv_data_426 : _GEN_7092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7094 = 9'h1ab == _GEN_15654 ? phv_data_427 : _GEN_7093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7095 = 9'h1ac == _GEN_15654 ? phv_data_428 : _GEN_7094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7096 = 9'h1ad == _GEN_15654 ? phv_data_429 : _GEN_7095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7097 = 9'h1ae == _GEN_15654 ? phv_data_430 : _GEN_7096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7098 = 9'h1af == _GEN_15654 ? phv_data_431 : _GEN_7097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7099 = 9'h1b0 == _GEN_15654 ? phv_data_432 : _GEN_7098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7100 = 9'h1b1 == _GEN_15654 ? phv_data_433 : _GEN_7099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7101 = 9'h1b2 == _GEN_15654 ? phv_data_434 : _GEN_7100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7102 = 9'h1b3 == _GEN_15654 ? phv_data_435 : _GEN_7101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7103 = 9'h1b4 == _GEN_15654 ? phv_data_436 : _GEN_7102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7104 = 9'h1b5 == _GEN_15654 ? phv_data_437 : _GEN_7103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7105 = 9'h1b6 == _GEN_15654 ? phv_data_438 : _GEN_7104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7106 = 9'h1b7 == _GEN_15654 ? phv_data_439 : _GEN_7105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7107 = 9'h1b8 == _GEN_15654 ? phv_data_440 : _GEN_7106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7108 = 9'h1b9 == _GEN_15654 ? phv_data_441 : _GEN_7107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7109 = 9'h1ba == _GEN_15654 ? phv_data_442 : _GEN_7108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7110 = 9'h1bb == _GEN_15654 ? phv_data_443 : _GEN_7109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7111 = 9'h1bc == _GEN_15654 ? phv_data_444 : _GEN_7110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7112 = 9'h1bd == _GEN_15654 ? phv_data_445 : _GEN_7111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7113 = 9'h1be == _GEN_15654 ? phv_data_446 : _GEN_7112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7114 = 9'h1bf == _GEN_15654 ? phv_data_447 : _GEN_7113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7115 = 9'h1c0 == _GEN_15654 ? phv_data_448 : _GEN_7114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7116 = 9'h1c1 == _GEN_15654 ? phv_data_449 : _GEN_7115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7117 = 9'h1c2 == _GEN_15654 ? phv_data_450 : _GEN_7116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7118 = 9'h1c3 == _GEN_15654 ? phv_data_451 : _GEN_7117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7119 = 9'h1c4 == _GEN_15654 ? phv_data_452 : _GEN_7118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7120 = 9'h1c5 == _GEN_15654 ? phv_data_453 : _GEN_7119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7121 = 9'h1c6 == _GEN_15654 ? phv_data_454 : _GEN_7120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7122 = 9'h1c7 == _GEN_15654 ? phv_data_455 : _GEN_7121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7123 = 9'h1c8 == _GEN_15654 ? phv_data_456 : _GEN_7122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7124 = 9'h1c9 == _GEN_15654 ? phv_data_457 : _GEN_7123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7125 = 9'h1ca == _GEN_15654 ? phv_data_458 : _GEN_7124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7126 = 9'h1cb == _GEN_15654 ? phv_data_459 : _GEN_7125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7127 = 9'h1cc == _GEN_15654 ? phv_data_460 : _GEN_7126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7128 = 9'h1cd == _GEN_15654 ? phv_data_461 : _GEN_7127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7129 = 9'h1ce == _GEN_15654 ? phv_data_462 : _GEN_7128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7130 = 9'h1cf == _GEN_15654 ? phv_data_463 : _GEN_7129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7131 = 9'h1d0 == _GEN_15654 ? phv_data_464 : _GEN_7130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7132 = 9'h1d1 == _GEN_15654 ? phv_data_465 : _GEN_7131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7133 = 9'h1d2 == _GEN_15654 ? phv_data_466 : _GEN_7132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7134 = 9'h1d3 == _GEN_15654 ? phv_data_467 : _GEN_7133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7135 = 9'h1d4 == _GEN_15654 ? phv_data_468 : _GEN_7134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7136 = 9'h1d5 == _GEN_15654 ? phv_data_469 : _GEN_7135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7137 = 9'h1d6 == _GEN_15654 ? phv_data_470 : _GEN_7136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7138 = 9'h1d7 == _GEN_15654 ? phv_data_471 : _GEN_7137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7139 = 9'h1d8 == _GEN_15654 ? phv_data_472 : _GEN_7138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7140 = 9'h1d9 == _GEN_15654 ? phv_data_473 : _GEN_7139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7141 = 9'h1da == _GEN_15654 ? phv_data_474 : _GEN_7140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7142 = 9'h1db == _GEN_15654 ? phv_data_475 : _GEN_7141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7143 = 9'h1dc == _GEN_15654 ? phv_data_476 : _GEN_7142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7144 = 9'h1dd == _GEN_15654 ? phv_data_477 : _GEN_7143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7145 = 9'h1de == _GEN_15654 ? phv_data_478 : _GEN_7144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7146 = 9'h1df == _GEN_15654 ? phv_data_479 : _GEN_7145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7147 = 9'h1e0 == _GEN_15654 ? phv_data_480 : _GEN_7146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7148 = 9'h1e1 == _GEN_15654 ? phv_data_481 : _GEN_7147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7149 = 9'h1e2 == _GEN_15654 ? phv_data_482 : _GEN_7148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7150 = 9'h1e3 == _GEN_15654 ? phv_data_483 : _GEN_7149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7151 = 9'h1e4 == _GEN_15654 ? phv_data_484 : _GEN_7150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7152 = 9'h1e5 == _GEN_15654 ? phv_data_485 : _GEN_7151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7153 = 9'h1e6 == _GEN_15654 ? phv_data_486 : _GEN_7152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7154 = 9'h1e7 == _GEN_15654 ? phv_data_487 : _GEN_7153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7155 = 9'h1e8 == _GEN_15654 ? phv_data_488 : _GEN_7154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7156 = 9'h1e9 == _GEN_15654 ? phv_data_489 : _GEN_7155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7157 = 9'h1ea == _GEN_15654 ? phv_data_490 : _GEN_7156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7158 = 9'h1eb == _GEN_15654 ? phv_data_491 : _GEN_7157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7159 = 9'h1ec == _GEN_15654 ? phv_data_492 : _GEN_7158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7160 = 9'h1ed == _GEN_15654 ? phv_data_493 : _GEN_7159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7161 = 9'h1ee == _GEN_15654 ? phv_data_494 : _GEN_7160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7162 = 9'h1ef == _GEN_15654 ? phv_data_495 : _GEN_7161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7163 = 9'h1f0 == _GEN_15654 ? phv_data_496 : _GEN_7162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7164 = 9'h1f1 == _GEN_15654 ? phv_data_497 : _GEN_7163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7165 = 9'h1f2 == _GEN_15654 ? phv_data_498 : _GEN_7164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7166 = 9'h1f3 == _GEN_15654 ? phv_data_499 : _GEN_7165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7167 = 9'h1f4 == _GEN_15654 ? phv_data_500 : _GEN_7166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7168 = 9'h1f5 == _GEN_15654 ? phv_data_501 : _GEN_7167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7169 = 9'h1f6 == _GEN_15654 ? phv_data_502 : _GEN_7168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7170 = 9'h1f7 == _GEN_15654 ? phv_data_503 : _GEN_7169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7171 = 9'h1f8 == _GEN_15654 ? phv_data_504 : _GEN_7170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7172 = 9'h1f9 == _GEN_15654 ? phv_data_505 : _GEN_7171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7173 = 9'h1fa == _GEN_15654 ? phv_data_506 : _GEN_7172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7174 = 9'h1fb == _GEN_15654 ? phv_data_507 : _GEN_7173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7175 = 9'h1fc == _GEN_15654 ? phv_data_508 : _GEN_7174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7176 = 9'h1fd == _GEN_15654 ? phv_data_509 : _GEN_7175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7177 = 9'h1fe == _GEN_15654 ? phv_data_510 : _GEN_7176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7178 = 9'h1ff == _GEN_15654 ? phv_data_511 : _GEN_7177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7180 = 8'h1 == _match_key_qbytes_3_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7181 = 8'h2 == _match_key_qbytes_3_T ? phv_data_2 : _GEN_7180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7182 = 8'h3 == _match_key_qbytes_3_T ? phv_data_3 : _GEN_7181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7183 = 8'h4 == _match_key_qbytes_3_T ? phv_data_4 : _GEN_7182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7184 = 8'h5 == _match_key_qbytes_3_T ? phv_data_5 : _GEN_7183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7185 = 8'h6 == _match_key_qbytes_3_T ? phv_data_6 : _GEN_7184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7186 = 8'h7 == _match_key_qbytes_3_T ? phv_data_7 : _GEN_7185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7187 = 8'h8 == _match_key_qbytes_3_T ? phv_data_8 : _GEN_7186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7188 = 8'h9 == _match_key_qbytes_3_T ? phv_data_9 : _GEN_7187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7189 = 8'ha == _match_key_qbytes_3_T ? phv_data_10 : _GEN_7188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7190 = 8'hb == _match_key_qbytes_3_T ? phv_data_11 : _GEN_7189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7191 = 8'hc == _match_key_qbytes_3_T ? phv_data_12 : _GEN_7190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7192 = 8'hd == _match_key_qbytes_3_T ? phv_data_13 : _GEN_7191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7193 = 8'he == _match_key_qbytes_3_T ? phv_data_14 : _GEN_7192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7194 = 8'hf == _match_key_qbytes_3_T ? phv_data_15 : _GEN_7193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7195 = 8'h10 == _match_key_qbytes_3_T ? phv_data_16 : _GEN_7194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7196 = 8'h11 == _match_key_qbytes_3_T ? phv_data_17 : _GEN_7195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7197 = 8'h12 == _match_key_qbytes_3_T ? phv_data_18 : _GEN_7196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7198 = 8'h13 == _match_key_qbytes_3_T ? phv_data_19 : _GEN_7197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7199 = 8'h14 == _match_key_qbytes_3_T ? phv_data_20 : _GEN_7198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7200 = 8'h15 == _match_key_qbytes_3_T ? phv_data_21 : _GEN_7199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7201 = 8'h16 == _match_key_qbytes_3_T ? phv_data_22 : _GEN_7200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7202 = 8'h17 == _match_key_qbytes_3_T ? phv_data_23 : _GEN_7201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7203 = 8'h18 == _match_key_qbytes_3_T ? phv_data_24 : _GEN_7202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7204 = 8'h19 == _match_key_qbytes_3_T ? phv_data_25 : _GEN_7203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7205 = 8'h1a == _match_key_qbytes_3_T ? phv_data_26 : _GEN_7204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7206 = 8'h1b == _match_key_qbytes_3_T ? phv_data_27 : _GEN_7205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7207 = 8'h1c == _match_key_qbytes_3_T ? phv_data_28 : _GEN_7206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7208 = 8'h1d == _match_key_qbytes_3_T ? phv_data_29 : _GEN_7207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7209 = 8'h1e == _match_key_qbytes_3_T ? phv_data_30 : _GEN_7208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7210 = 8'h1f == _match_key_qbytes_3_T ? phv_data_31 : _GEN_7209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7211 = 8'h20 == _match_key_qbytes_3_T ? phv_data_32 : _GEN_7210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7212 = 8'h21 == _match_key_qbytes_3_T ? phv_data_33 : _GEN_7211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7213 = 8'h22 == _match_key_qbytes_3_T ? phv_data_34 : _GEN_7212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7214 = 8'h23 == _match_key_qbytes_3_T ? phv_data_35 : _GEN_7213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7215 = 8'h24 == _match_key_qbytes_3_T ? phv_data_36 : _GEN_7214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7216 = 8'h25 == _match_key_qbytes_3_T ? phv_data_37 : _GEN_7215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7217 = 8'h26 == _match_key_qbytes_3_T ? phv_data_38 : _GEN_7216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7218 = 8'h27 == _match_key_qbytes_3_T ? phv_data_39 : _GEN_7217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7219 = 8'h28 == _match_key_qbytes_3_T ? phv_data_40 : _GEN_7218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7220 = 8'h29 == _match_key_qbytes_3_T ? phv_data_41 : _GEN_7219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7221 = 8'h2a == _match_key_qbytes_3_T ? phv_data_42 : _GEN_7220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7222 = 8'h2b == _match_key_qbytes_3_T ? phv_data_43 : _GEN_7221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7223 = 8'h2c == _match_key_qbytes_3_T ? phv_data_44 : _GEN_7222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7224 = 8'h2d == _match_key_qbytes_3_T ? phv_data_45 : _GEN_7223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7225 = 8'h2e == _match_key_qbytes_3_T ? phv_data_46 : _GEN_7224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7226 = 8'h2f == _match_key_qbytes_3_T ? phv_data_47 : _GEN_7225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7227 = 8'h30 == _match_key_qbytes_3_T ? phv_data_48 : _GEN_7226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7228 = 8'h31 == _match_key_qbytes_3_T ? phv_data_49 : _GEN_7227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7229 = 8'h32 == _match_key_qbytes_3_T ? phv_data_50 : _GEN_7228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7230 = 8'h33 == _match_key_qbytes_3_T ? phv_data_51 : _GEN_7229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7231 = 8'h34 == _match_key_qbytes_3_T ? phv_data_52 : _GEN_7230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7232 = 8'h35 == _match_key_qbytes_3_T ? phv_data_53 : _GEN_7231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7233 = 8'h36 == _match_key_qbytes_3_T ? phv_data_54 : _GEN_7232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7234 = 8'h37 == _match_key_qbytes_3_T ? phv_data_55 : _GEN_7233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7235 = 8'h38 == _match_key_qbytes_3_T ? phv_data_56 : _GEN_7234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7236 = 8'h39 == _match_key_qbytes_3_T ? phv_data_57 : _GEN_7235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7237 = 8'h3a == _match_key_qbytes_3_T ? phv_data_58 : _GEN_7236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7238 = 8'h3b == _match_key_qbytes_3_T ? phv_data_59 : _GEN_7237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7239 = 8'h3c == _match_key_qbytes_3_T ? phv_data_60 : _GEN_7238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7240 = 8'h3d == _match_key_qbytes_3_T ? phv_data_61 : _GEN_7239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7241 = 8'h3e == _match_key_qbytes_3_T ? phv_data_62 : _GEN_7240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7242 = 8'h3f == _match_key_qbytes_3_T ? phv_data_63 : _GEN_7241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7243 = 8'h40 == _match_key_qbytes_3_T ? phv_data_64 : _GEN_7242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7244 = 8'h41 == _match_key_qbytes_3_T ? phv_data_65 : _GEN_7243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7245 = 8'h42 == _match_key_qbytes_3_T ? phv_data_66 : _GEN_7244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7246 = 8'h43 == _match_key_qbytes_3_T ? phv_data_67 : _GEN_7245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7247 = 8'h44 == _match_key_qbytes_3_T ? phv_data_68 : _GEN_7246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7248 = 8'h45 == _match_key_qbytes_3_T ? phv_data_69 : _GEN_7247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7249 = 8'h46 == _match_key_qbytes_3_T ? phv_data_70 : _GEN_7248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7250 = 8'h47 == _match_key_qbytes_3_T ? phv_data_71 : _GEN_7249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7251 = 8'h48 == _match_key_qbytes_3_T ? phv_data_72 : _GEN_7250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7252 = 8'h49 == _match_key_qbytes_3_T ? phv_data_73 : _GEN_7251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7253 = 8'h4a == _match_key_qbytes_3_T ? phv_data_74 : _GEN_7252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7254 = 8'h4b == _match_key_qbytes_3_T ? phv_data_75 : _GEN_7253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7255 = 8'h4c == _match_key_qbytes_3_T ? phv_data_76 : _GEN_7254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7256 = 8'h4d == _match_key_qbytes_3_T ? phv_data_77 : _GEN_7255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7257 = 8'h4e == _match_key_qbytes_3_T ? phv_data_78 : _GEN_7256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7258 = 8'h4f == _match_key_qbytes_3_T ? phv_data_79 : _GEN_7257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7259 = 8'h50 == _match_key_qbytes_3_T ? phv_data_80 : _GEN_7258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7260 = 8'h51 == _match_key_qbytes_3_T ? phv_data_81 : _GEN_7259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7261 = 8'h52 == _match_key_qbytes_3_T ? phv_data_82 : _GEN_7260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7262 = 8'h53 == _match_key_qbytes_3_T ? phv_data_83 : _GEN_7261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7263 = 8'h54 == _match_key_qbytes_3_T ? phv_data_84 : _GEN_7262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7264 = 8'h55 == _match_key_qbytes_3_T ? phv_data_85 : _GEN_7263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7265 = 8'h56 == _match_key_qbytes_3_T ? phv_data_86 : _GEN_7264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7266 = 8'h57 == _match_key_qbytes_3_T ? phv_data_87 : _GEN_7265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7267 = 8'h58 == _match_key_qbytes_3_T ? phv_data_88 : _GEN_7266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7268 = 8'h59 == _match_key_qbytes_3_T ? phv_data_89 : _GEN_7267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7269 = 8'h5a == _match_key_qbytes_3_T ? phv_data_90 : _GEN_7268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7270 = 8'h5b == _match_key_qbytes_3_T ? phv_data_91 : _GEN_7269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7271 = 8'h5c == _match_key_qbytes_3_T ? phv_data_92 : _GEN_7270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7272 = 8'h5d == _match_key_qbytes_3_T ? phv_data_93 : _GEN_7271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7273 = 8'h5e == _match_key_qbytes_3_T ? phv_data_94 : _GEN_7272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7274 = 8'h5f == _match_key_qbytes_3_T ? phv_data_95 : _GEN_7273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7275 = 8'h60 == _match_key_qbytes_3_T ? phv_data_96 : _GEN_7274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7276 = 8'h61 == _match_key_qbytes_3_T ? phv_data_97 : _GEN_7275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7277 = 8'h62 == _match_key_qbytes_3_T ? phv_data_98 : _GEN_7276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7278 = 8'h63 == _match_key_qbytes_3_T ? phv_data_99 : _GEN_7277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7279 = 8'h64 == _match_key_qbytes_3_T ? phv_data_100 : _GEN_7278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7280 = 8'h65 == _match_key_qbytes_3_T ? phv_data_101 : _GEN_7279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7281 = 8'h66 == _match_key_qbytes_3_T ? phv_data_102 : _GEN_7280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7282 = 8'h67 == _match_key_qbytes_3_T ? phv_data_103 : _GEN_7281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7283 = 8'h68 == _match_key_qbytes_3_T ? phv_data_104 : _GEN_7282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7284 = 8'h69 == _match_key_qbytes_3_T ? phv_data_105 : _GEN_7283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7285 = 8'h6a == _match_key_qbytes_3_T ? phv_data_106 : _GEN_7284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7286 = 8'h6b == _match_key_qbytes_3_T ? phv_data_107 : _GEN_7285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7287 = 8'h6c == _match_key_qbytes_3_T ? phv_data_108 : _GEN_7286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7288 = 8'h6d == _match_key_qbytes_3_T ? phv_data_109 : _GEN_7287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7289 = 8'h6e == _match_key_qbytes_3_T ? phv_data_110 : _GEN_7288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7290 = 8'h6f == _match_key_qbytes_3_T ? phv_data_111 : _GEN_7289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7291 = 8'h70 == _match_key_qbytes_3_T ? phv_data_112 : _GEN_7290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7292 = 8'h71 == _match_key_qbytes_3_T ? phv_data_113 : _GEN_7291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7293 = 8'h72 == _match_key_qbytes_3_T ? phv_data_114 : _GEN_7292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7294 = 8'h73 == _match_key_qbytes_3_T ? phv_data_115 : _GEN_7293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7295 = 8'h74 == _match_key_qbytes_3_T ? phv_data_116 : _GEN_7294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7296 = 8'h75 == _match_key_qbytes_3_T ? phv_data_117 : _GEN_7295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7297 = 8'h76 == _match_key_qbytes_3_T ? phv_data_118 : _GEN_7296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7298 = 8'h77 == _match_key_qbytes_3_T ? phv_data_119 : _GEN_7297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7299 = 8'h78 == _match_key_qbytes_3_T ? phv_data_120 : _GEN_7298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7300 = 8'h79 == _match_key_qbytes_3_T ? phv_data_121 : _GEN_7299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7301 = 8'h7a == _match_key_qbytes_3_T ? phv_data_122 : _GEN_7300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7302 = 8'h7b == _match_key_qbytes_3_T ? phv_data_123 : _GEN_7301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7303 = 8'h7c == _match_key_qbytes_3_T ? phv_data_124 : _GEN_7302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7304 = 8'h7d == _match_key_qbytes_3_T ? phv_data_125 : _GEN_7303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7305 = 8'h7e == _match_key_qbytes_3_T ? phv_data_126 : _GEN_7304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7306 = 8'h7f == _match_key_qbytes_3_T ? phv_data_127 : _GEN_7305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7307 = 8'h80 == _match_key_qbytes_3_T ? phv_data_128 : _GEN_7306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7308 = 8'h81 == _match_key_qbytes_3_T ? phv_data_129 : _GEN_7307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7309 = 8'h82 == _match_key_qbytes_3_T ? phv_data_130 : _GEN_7308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7310 = 8'h83 == _match_key_qbytes_3_T ? phv_data_131 : _GEN_7309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7311 = 8'h84 == _match_key_qbytes_3_T ? phv_data_132 : _GEN_7310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7312 = 8'h85 == _match_key_qbytes_3_T ? phv_data_133 : _GEN_7311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7313 = 8'h86 == _match_key_qbytes_3_T ? phv_data_134 : _GEN_7312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7314 = 8'h87 == _match_key_qbytes_3_T ? phv_data_135 : _GEN_7313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7315 = 8'h88 == _match_key_qbytes_3_T ? phv_data_136 : _GEN_7314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7316 = 8'h89 == _match_key_qbytes_3_T ? phv_data_137 : _GEN_7315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7317 = 8'h8a == _match_key_qbytes_3_T ? phv_data_138 : _GEN_7316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7318 = 8'h8b == _match_key_qbytes_3_T ? phv_data_139 : _GEN_7317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7319 = 8'h8c == _match_key_qbytes_3_T ? phv_data_140 : _GEN_7318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7320 = 8'h8d == _match_key_qbytes_3_T ? phv_data_141 : _GEN_7319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7321 = 8'h8e == _match_key_qbytes_3_T ? phv_data_142 : _GEN_7320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7322 = 8'h8f == _match_key_qbytes_3_T ? phv_data_143 : _GEN_7321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7323 = 8'h90 == _match_key_qbytes_3_T ? phv_data_144 : _GEN_7322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7324 = 8'h91 == _match_key_qbytes_3_T ? phv_data_145 : _GEN_7323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7325 = 8'h92 == _match_key_qbytes_3_T ? phv_data_146 : _GEN_7324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7326 = 8'h93 == _match_key_qbytes_3_T ? phv_data_147 : _GEN_7325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7327 = 8'h94 == _match_key_qbytes_3_T ? phv_data_148 : _GEN_7326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7328 = 8'h95 == _match_key_qbytes_3_T ? phv_data_149 : _GEN_7327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7329 = 8'h96 == _match_key_qbytes_3_T ? phv_data_150 : _GEN_7328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7330 = 8'h97 == _match_key_qbytes_3_T ? phv_data_151 : _GEN_7329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7331 = 8'h98 == _match_key_qbytes_3_T ? phv_data_152 : _GEN_7330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7332 = 8'h99 == _match_key_qbytes_3_T ? phv_data_153 : _GEN_7331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7333 = 8'h9a == _match_key_qbytes_3_T ? phv_data_154 : _GEN_7332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7334 = 8'h9b == _match_key_qbytes_3_T ? phv_data_155 : _GEN_7333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7335 = 8'h9c == _match_key_qbytes_3_T ? phv_data_156 : _GEN_7334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7336 = 8'h9d == _match_key_qbytes_3_T ? phv_data_157 : _GEN_7335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7337 = 8'h9e == _match_key_qbytes_3_T ? phv_data_158 : _GEN_7336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7338 = 8'h9f == _match_key_qbytes_3_T ? phv_data_159 : _GEN_7337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7339 = 8'ha0 == _match_key_qbytes_3_T ? phv_data_160 : _GEN_7338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7340 = 8'ha1 == _match_key_qbytes_3_T ? phv_data_161 : _GEN_7339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7341 = 8'ha2 == _match_key_qbytes_3_T ? phv_data_162 : _GEN_7340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7342 = 8'ha3 == _match_key_qbytes_3_T ? phv_data_163 : _GEN_7341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7343 = 8'ha4 == _match_key_qbytes_3_T ? phv_data_164 : _GEN_7342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7344 = 8'ha5 == _match_key_qbytes_3_T ? phv_data_165 : _GEN_7343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7345 = 8'ha6 == _match_key_qbytes_3_T ? phv_data_166 : _GEN_7344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7346 = 8'ha7 == _match_key_qbytes_3_T ? phv_data_167 : _GEN_7345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7347 = 8'ha8 == _match_key_qbytes_3_T ? phv_data_168 : _GEN_7346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7348 = 8'ha9 == _match_key_qbytes_3_T ? phv_data_169 : _GEN_7347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7349 = 8'haa == _match_key_qbytes_3_T ? phv_data_170 : _GEN_7348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7350 = 8'hab == _match_key_qbytes_3_T ? phv_data_171 : _GEN_7349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7351 = 8'hac == _match_key_qbytes_3_T ? phv_data_172 : _GEN_7350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7352 = 8'had == _match_key_qbytes_3_T ? phv_data_173 : _GEN_7351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7353 = 8'hae == _match_key_qbytes_3_T ? phv_data_174 : _GEN_7352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7354 = 8'haf == _match_key_qbytes_3_T ? phv_data_175 : _GEN_7353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7355 = 8'hb0 == _match_key_qbytes_3_T ? phv_data_176 : _GEN_7354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7356 = 8'hb1 == _match_key_qbytes_3_T ? phv_data_177 : _GEN_7355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7357 = 8'hb2 == _match_key_qbytes_3_T ? phv_data_178 : _GEN_7356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7358 = 8'hb3 == _match_key_qbytes_3_T ? phv_data_179 : _GEN_7357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7359 = 8'hb4 == _match_key_qbytes_3_T ? phv_data_180 : _GEN_7358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7360 = 8'hb5 == _match_key_qbytes_3_T ? phv_data_181 : _GEN_7359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7361 = 8'hb6 == _match_key_qbytes_3_T ? phv_data_182 : _GEN_7360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7362 = 8'hb7 == _match_key_qbytes_3_T ? phv_data_183 : _GEN_7361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7363 = 8'hb8 == _match_key_qbytes_3_T ? phv_data_184 : _GEN_7362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7364 = 8'hb9 == _match_key_qbytes_3_T ? phv_data_185 : _GEN_7363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7365 = 8'hba == _match_key_qbytes_3_T ? phv_data_186 : _GEN_7364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7366 = 8'hbb == _match_key_qbytes_3_T ? phv_data_187 : _GEN_7365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7367 = 8'hbc == _match_key_qbytes_3_T ? phv_data_188 : _GEN_7366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7368 = 8'hbd == _match_key_qbytes_3_T ? phv_data_189 : _GEN_7367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7369 = 8'hbe == _match_key_qbytes_3_T ? phv_data_190 : _GEN_7368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7370 = 8'hbf == _match_key_qbytes_3_T ? phv_data_191 : _GEN_7369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7371 = 8'hc0 == _match_key_qbytes_3_T ? phv_data_192 : _GEN_7370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7372 = 8'hc1 == _match_key_qbytes_3_T ? phv_data_193 : _GEN_7371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7373 = 8'hc2 == _match_key_qbytes_3_T ? phv_data_194 : _GEN_7372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7374 = 8'hc3 == _match_key_qbytes_3_T ? phv_data_195 : _GEN_7373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7375 = 8'hc4 == _match_key_qbytes_3_T ? phv_data_196 : _GEN_7374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7376 = 8'hc5 == _match_key_qbytes_3_T ? phv_data_197 : _GEN_7375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7377 = 8'hc6 == _match_key_qbytes_3_T ? phv_data_198 : _GEN_7376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7378 = 8'hc7 == _match_key_qbytes_3_T ? phv_data_199 : _GEN_7377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7379 = 8'hc8 == _match_key_qbytes_3_T ? phv_data_200 : _GEN_7378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7380 = 8'hc9 == _match_key_qbytes_3_T ? phv_data_201 : _GEN_7379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7381 = 8'hca == _match_key_qbytes_3_T ? phv_data_202 : _GEN_7380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7382 = 8'hcb == _match_key_qbytes_3_T ? phv_data_203 : _GEN_7381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7383 = 8'hcc == _match_key_qbytes_3_T ? phv_data_204 : _GEN_7382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7384 = 8'hcd == _match_key_qbytes_3_T ? phv_data_205 : _GEN_7383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7385 = 8'hce == _match_key_qbytes_3_T ? phv_data_206 : _GEN_7384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7386 = 8'hcf == _match_key_qbytes_3_T ? phv_data_207 : _GEN_7385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7387 = 8'hd0 == _match_key_qbytes_3_T ? phv_data_208 : _GEN_7386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7388 = 8'hd1 == _match_key_qbytes_3_T ? phv_data_209 : _GEN_7387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7389 = 8'hd2 == _match_key_qbytes_3_T ? phv_data_210 : _GEN_7388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7390 = 8'hd3 == _match_key_qbytes_3_T ? phv_data_211 : _GEN_7389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7391 = 8'hd4 == _match_key_qbytes_3_T ? phv_data_212 : _GEN_7390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7392 = 8'hd5 == _match_key_qbytes_3_T ? phv_data_213 : _GEN_7391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7393 = 8'hd6 == _match_key_qbytes_3_T ? phv_data_214 : _GEN_7392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7394 = 8'hd7 == _match_key_qbytes_3_T ? phv_data_215 : _GEN_7393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7395 = 8'hd8 == _match_key_qbytes_3_T ? phv_data_216 : _GEN_7394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7396 = 8'hd9 == _match_key_qbytes_3_T ? phv_data_217 : _GEN_7395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7397 = 8'hda == _match_key_qbytes_3_T ? phv_data_218 : _GEN_7396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7398 = 8'hdb == _match_key_qbytes_3_T ? phv_data_219 : _GEN_7397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7399 = 8'hdc == _match_key_qbytes_3_T ? phv_data_220 : _GEN_7398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7400 = 8'hdd == _match_key_qbytes_3_T ? phv_data_221 : _GEN_7399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7401 = 8'hde == _match_key_qbytes_3_T ? phv_data_222 : _GEN_7400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7402 = 8'hdf == _match_key_qbytes_3_T ? phv_data_223 : _GEN_7401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7403 = 8'he0 == _match_key_qbytes_3_T ? phv_data_224 : _GEN_7402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7404 = 8'he1 == _match_key_qbytes_3_T ? phv_data_225 : _GEN_7403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7405 = 8'he2 == _match_key_qbytes_3_T ? phv_data_226 : _GEN_7404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7406 = 8'he3 == _match_key_qbytes_3_T ? phv_data_227 : _GEN_7405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7407 = 8'he4 == _match_key_qbytes_3_T ? phv_data_228 : _GEN_7406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7408 = 8'he5 == _match_key_qbytes_3_T ? phv_data_229 : _GEN_7407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7409 = 8'he6 == _match_key_qbytes_3_T ? phv_data_230 : _GEN_7408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7410 = 8'he7 == _match_key_qbytes_3_T ? phv_data_231 : _GEN_7409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7411 = 8'he8 == _match_key_qbytes_3_T ? phv_data_232 : _GEN_7410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7412 = 8'he9 == _match_key_qbytes_3_T ? phv_data_233 : _GEN_7411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7413 = 8'hea == _match_key_qbytes_3_T ? phv_data_234 : _GEN_7412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7414 = 8'heb == _match_key_qbytes_3_T ? phv_data_235 : _GEN_7413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7415 = 8'hec == _match_key_qbytes_3_T ? phv_data_236 : _GEN_7414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7416 = 8'hed == _match_key_qbytes_3_T ? phv_data_237 : _GEN_7415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7417 = 8'hee == _match_key_qbytes_3_T ? phv_data_238 : _GEN_7416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7418 = 8'hef == _match_key_qbytes_3_T ? phv_data_239 : _GEN_7417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7419 = 8'hf0 == _match_key_qbytes_3_T ? phv_data_240 : _GEN_7418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7420 = 8'hf1 == _match_key_qbytes_3_T ? phv_data_241 : _GEN_7419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7421 = 8'hf2 == _match_key_qbytes_3_T ? phv_data_242 : _GEN_7420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7422 = 8'hf3 == _match_key_qbytes_3_T ? phv_data_243 : _GEN_7421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7423 = 8'hf4 == _match_key_qbytes_3_T ? phv_data_244 : _GEN_7422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7424 = 8'hf5 == _match_key_qbytes_3_T ? phv_data_245 : _GEN_7423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7425 = 8'hf6 == _match_key_qbytes_3_T ? phv_data_246 : _GEN_7424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7426 = 8'hf7 == _match_key_qbytes_3_T ? phv_data_247 : _GEN_7425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7427 = 8'hf8 == _match_key_qbytes_3_T ? phv_data_248 : _GEN_7426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7428 = 8'hf9 == _match_key_qbytes_3_T ? phv_data_249 : _GEN_7427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7429 = 8'hfa == _match_key_qbytes_3_T ? phv_data_250 : _GEN_7428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7430 = 8'hfb == _match_key_qbytes_3_T ? phv_data_251 : _GEN_7429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7431 = 8'hfc == _match_key_qbytes_3_T ? phv_data_252 : _GEN_7430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7432 = 8'hfd == _match_key_qbytes_3_T ? phv_data_253 : _GEN_7431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7433 = 8'hfe == _match_key_qbytes_3_T ? phv_data_254 : _GEN_7432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7434 = 8'hff == _match_key_qbytes_3_T ? phv_data_255 : _GEN_7433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_15910 = {{1'd0}, _match_key_qbytes_3_T}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7435 = 9'h100 == _GEN_15910 ? phv_data_256 : _GEN_7434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7436 = 9'h101 == _GEN_15910 ? phv_data_257 : _GEN_7435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7437 = 9'h102 == _GEN_15910 ? phv_data_258 : _GEN_7436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7438 = 9'h103 == _GEN_15910 ? phv_data_259 : _GEN_7437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7439 = 9'h104 == _GEN_15910 ? phv_data_260 : _GEN_7438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7440 = 9'h105 == _GEN_15910 ? phv_data_261 : _GEN_7439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7441 = 9'h106 == _GEN_15910 ? phv_data_262 : _GEN_7440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7442 = 9'h107 == _GEN_15910 ? phv_data_263 : _GEN_7441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7443 = 9'h108 == _GEN_15910 ? phv_data_264 : _GEN_7442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7444 = 9'h109 == _GEN_15910 ? phv_data_265 : _GEN_7443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7445 = 9'h10a == _GEN_15910 ? phv_data_266 : _GEN_7444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7446 = 9'h10b == _GEN_15910 ? phv_data_267 : _GEN_7445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7447 = 9'h10c == _GEN_15910 ? phv_data_268 : _GEN_7446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7448 = 9'h10d == _GEN_15910 ? phv_data_269 : _GEN_7447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7449 = 9'h10e == _GEN_15910 ? phv_data_270 : _GEN_7448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7450 = 9'h10f == _GEN_15910 ? phv_data_271 : _GEN_7449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7451 = 9'h110 == _GEN_15910 ? phv_data_272 : _GEN_7450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7452 = 9'h111 == _GEN_15910 ? phv_data_273 : _GEN_7451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7453 = 9'h112 == _GEN_15910 ? phv_data_274 : _GEN_7452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7454 = 9'h113 == _GEN_15910 ? phv_data_275 : _GEN_7453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7455 = 9'h114 == _GEN_15910 ? phv_data_276 : _GEN_7454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7456 = 9'h115 == _GEN_15910 ? phv_data_277 : _GEN_7455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7457 = 9'h116 == _GEN_15910 ? phv_data_278 : _GEN_7456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7458 = 9'h117 == _GEN_15910 ? phv_data_279 : _GEN_7457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7459 = 9'h118 == _GEN_15910 ? phv_data_280 : _GEN_7458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7460 = 9'h119 == _GEN_15910 ? phv_data_281 : _GEN_7459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7461 = 9'h11a == _GEN_15910 ? phv_data_282 : _GEN_7460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7462 = 9'h11b == _GEN_15910 ? phv_data_283 : _GEN_7461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7463 = 9'h11c == _GEN_15910 ? phv_data_284 : _GEN_7462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7464 = 9'h11d == _GEN_15910 ? phv_data_285 : _GEN_7463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7465 = 9'h11e == _GEN_15910 ? phv_data_286 : _GEN_7464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7466 = 9'h11f == _GEN_15910 ? phv_data_287 : _GEN_7465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7467 = 9'h120 == _GEN_15910 ? phv_data_288 : _GEN_7466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7468 = 9'h121 == _GEN_15910 ? phv_data_289 : _GEN_7467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7469 = 9'h122 == _GEN_15910 ? phv_data_290 : _GEN_7468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7470 = 9'h123 == _GEN_15910 ? phv_data_291 : _GEN_7469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7471 = 9'h124 == _GEN_15910 ? phv_data_292 : _GEN_7470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7472 = 9'h125 == _GEN_15910 ? phv_data_293 : _GEN_7471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7473 = 9'h126 == _GEN_15910 ? phv_data_294 : _GEN_7472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7474 = 9'h127 == _GEN_15910 ? phv_data_295 : _GEN_7473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7475 = 9'h128 == _GEN_15910 ? phv_data_296 : _GEN_7474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7476 = 9'h129 == _GEN_15910 ? phv_data_297 : _GEN_7475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7477 = 9'h12a == _GEN_15910 ? phv_data_298 : _GEN_7476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7478 = 9'h12b == _GEN_15910 ? phv_data_299 : _GEN_7477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7479 = 9'h12c == _GEN_15910 ? phv_data_300 : _GEN_7478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7480 = 9'h12d == _GEN_15910 ? phv_data_301 : _GEN_7479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7481 = 9'h12e == _GEN_15910 ? phv_data_302 : _GEN_7480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7482 = 9'h12f == _GEN_15910 ? phv_data_303 : _GEN_7481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7483 = 9'h130 == _GEN_15910 ? phv_data_304 : _GEN_7482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7484 = 9'h131 == _GEN_15910 ? phv_data_305 : _GEN_7483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7485 = 9'h132 == _GEN_15910 ? phv_data_306 : _GEN_7484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7486 = 9'h133 == _GEN_15910 ? phv_data_307 : _GEN_7485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7487 = 9'h134 == _GEN_15910 ? phv_data_308 : _GEN_7486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7488 = 9'h135 == _GEN_15910 ? phv_data_309 : _GEN_7487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7489 = 9'h136 == _GEN_15910 ? phv_data_310 : _GEN_7488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7490 = 9'h137 == _GEN_15910 ? phv_data_311 : _GEN_7489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7491 = 9'h138 == _GEN_15910 ? phv_data_312 : _GEN_7490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7492 = 9'h139 == _GEN_15910 ? phv_data_313 : _GEN_7491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7493 = 9'h13a == _GEN_15910 ? phv_data_314 : _GEN_7492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7494 = 9'h13b == _GEN_15910 ? phv_data_315 : _GEN_7493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7495 = 9'h13c == _GEN_15910 ? phv_data_316 : _GEN_7494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7496 = 9'h13d == _GEN_15910 ? phv_data_317 : _GEN_7495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7497 = 9'h13e == _GEN_15910 ? phv_data_318 : _GEN_7496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7498 = 9'h13f == _GEN_15910 ? phv_data_319 : _GEN_7497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7499 = 9'h140 == _GEN_15910 ? phv_data_320 : _GEN_7498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7500 = 9'h141 == _GEN_15910 ? phv_data_321 : _GEN_7499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7501 = 9'h142 == _GEN_15910 ? phv_data_322 : _GEN_7500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7502 = 9'h143 == _GEN_15910 ? phv_data_323 : _GEN_7501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7503 = 9'h144 == _GEN_15910 ? phv_data_324 : _GEN_7502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7504 = 9'h145 == _GEN_15910 ? phv_data_325 : _GEN_7503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7505 = 9'h146 == _GEN_15910 ? phv_data_326 : _GEN_7504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7506 = 9'h147 == _GEN_15910 ? phv_data_327 : _GEN_7505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7507 = 9'h148 == _GEN_15910 ? phv_data_328 : _GEN_7506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7508 = 9'h149 == _GEN_15910 ? phv_data_329 : _GEN_7507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7509 = 9'h14a == _GEN_15910 ? phv_data_330 : _GEN_7508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7510 = 9'h14b == _GEN_15910 ? phv_data_331 : _GEN_7509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7511 = 9'h14c == _GEN_15910 ? phv_data_332 : _GEN_7510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7512 = 9'h14d == _GEN_15910 ? phv_data_333 : _GEN_7511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7513 = 9'h14e == _GEN_15910 ? phv_data_334 : _GEN_7512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7514 = 9'h14f == _GEN_15910 ? phv_data_335 : _GEN_7513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7515 = 9'h150 == _GEN_15910 ? phv_data_336 : _GEN_7514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7516 = 9'h151 == _GEN_15910 ? phv_data_337 : _GEN_7515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7517 = 9'h152 == _GEN_15910 ? phv_data_338 : _GEN_7516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7518 = 9'h153 == _GEN_15910 ? phv_data_339 : _GEN_7517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7519 = 9'h154 == _GEN_15910 ? phv_data_340 : _GEN_7518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7520 = 9'h155 == _GEN_15910 ? phv_data_341 : _GEN_7519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7521 = 9'h156 == _GEN_15910 ? phv_data_342 : _GEN_7520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7522 = 9'h157 == _GEN_15910 ? phv_data_343 : _GEN_7521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7523 = 9'h158 == _GEN_15910 ? phv_data_344 : _GEN_7522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7524 = 9'h159 == _GEN_15910 ? phv_data_345 : _GEN_7523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7525 = 9'h15a == _GEN_15910 ? phv_data_346 : _GEN_7524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7526 = 9'h15b == _GEN_15910 ? phv_data_347 : _GEN_7525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7527 = 9'h15c == _GEN_15910 ? phv_data_348 : _GEN_7526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7528 = 9'h15d == _GEN_15910 ? phv_data_349 : _GEN_7527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7529 = 9'h15e == _GEN_15910 ? phv_data_350 : _GEN_7528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7530 = 9'h15f == _GEN_15910 ? phv_data_351 : _GEN_7529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7531 = 9'h160 == _GEN_15910 ? phv_data_352 : _GEN_7530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7532 = 9'h161 == _GEN_15910 ? phv_data_353 : _GEN_7531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7533 = 9'h162 == _GEN_15910 ? phv_data_354 : _GEN_7532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7534 = 9'h163 == _GEN_15910 ? phv_data_355 : _GEN_7533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7535 = 9'h164 == _GEN_15910 ? phv_data_356 : _GEN_7534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7536 = 9'h165 == _GEN_15910 ? phv_data_357 : _GEN_7535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7537 = 9'h166 == _GEN_15910 ? phv_data_358 : _GEN_7536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7538 = 9'h167 == _GEN_15910 ? phv_data_359 : _GEN_7537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7539 = 9'h168 == _GEN_15910 ? phv_data_360 : _GEN_7538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7540 = 9'h169 == _GEN_15910 ? phv_data_361 : _GEN_7539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7541 = 9'h16a == _GEN_15910 ? phv_data_362 : _GEN_7540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7542 = 9'h16b == _GEN_15910 ? phv_data_363 : _GEN_7541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7543 = 9'h16c == _GEN_15910 ? phv_data_364 : _GEN_7542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7544 = 9'h16d == _GEN_15910 ? phv_data_365 : _GEN_7543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7545 = 9'h16e == _GEN_15910 ? phv_data_366 : _GEN_7544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7546 = 9'h16f == _GEN_15910 ? phv_data_367 : _GEN_7545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7547 = 9'h170 == _GEN_15910 ? phv_data_368 : _GEN_7546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7548 = 9'h171 == _GEN_15910 ? phv_data_369 : _GEN_7547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7549 = 9'h172 == _GEN_15910 ? phv_data_370 : _GEN_7548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7550 = 9'h173 == _GEN_15910 ? phv_data_371 : _GEN_7549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7551 = 9'h174 == _GEN_15910 ? phv_data_372 : _GEN_7550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7552 = 9'h175 == _GEN_15910 ? phv_data_373 : _GEN_7551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7553 = 9'h176 == _GEN_15910 ? phv_data_374 : _GEN_7552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7554 = 9'h177 == _GEN_15910 ? phv_data_375 : _GEN_7553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7555 = 9'h178 == _GEN_15910 ? phv_data_376 : _GEN_7554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7556 = 9'h179 == _GEN_15910 ? phv_data_377 : _GEN_7555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7557 = 9'h17a == _GEN_15910 ? phv_data_378 : _GEN_7556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7558 = 9'h17b == _GEN_15910 ? phv_data_379 : _GEN_7557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7559 = 9'h17c == _GEN_15910 ? phv_data_380 : _GEN_7558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7560 = 9'h17d == _GEN_15910 ? phv_data_381 : _GEN_7559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7561 = 9'h17e == _GEN_15910 ? phv_data_382 : _GEN_7560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7562 = 9'h17f == _GEN_15910 ? phv_data_383 : _GEN_7561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7563 = 9'h180 == _GEN_15910 ? phv_data_384 : _GEN_7562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7564 = 9'h181 == _GEN_15910 ? phv_data_385 : _GEN_7563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7565 = 9'h182 == _GEN_15910 ? phv_data_386 : _GEN_7564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7566 = 9'h183 == _GEN_15910 ? phv_data_387 : _GEN_7565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7567 = 9'h184 == _GEN_15910 ? phv_data_388 : _GEN_7566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7568 = 9'h185 == _GEN_15910 ? phv_data_389 : _GEN_7567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7569 = 9'h186 == _GEN_15910 ? phv_data_390 : _GEN_7568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7570 = 9'h187 == _GEN_15910 ? phv_data_391 : _GEN_7569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7571 = 9'h188 == _GEN_15910 ? phv_data_392 : _GEN_7570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7572 = 9'h189 == _GEN_15910 ? phv_data_393 : _GEN_7571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7573 = 9'h18a == _GEN_15910 ? phv_data_394 : _GEN_7572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7574 = 9'h18b == _GEN_15910 ? phv_data_395 : _GEN_7573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7575 = 9'h18c == _GEN_15910 ? phv_data_396 : _GEN_7574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7576 = 9'h18d == _GEN_15910 ? phv_data_397 : _GEN_7575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7577 = 9'h18e == _GEN_15910 ? phv_data_398 : _GEN_7576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7578 = 9'h18f == _GEN_15910 ? phv_data_399 : _GEN_7577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7579 = 9'h190 == _GEN_15910 ? phv_data_400 : _GEN_7578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7580 = 9'h191 == _GEN_15910 ? phv_data_401 : _GEN_7579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7581 = 9'h192 == _GEN_15910 ? phv_data_402 : _GEN_7580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7582 = 9'h193 == _GEN_15910 ? phv_data_403 : _GEN_7581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7583 = 9'h194 == _GEN_15910 ? phv_data_404 : _GEN_7582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7584 = 9'h195 == _GEN_15910 ? phv_data_405 : _GEN_7583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7585 = 9'h196 == _GEN_15910 ? phv_data_406 : _GEN_7584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7586 = 9'h197 == _GEN_15910 ? phv_data_407 : _GEN_7585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7587 = 9'h198 == _GEN_15910 ? phv_data_408 : _GEN_7586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7588 = 9'h199 == _GEN_15910 ? phv_data_409 : _GEN_7587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7589 = 9'h19a == _GEN_15910 ? phv_data_410 : _GEN_7588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7590 = 9'h19b == _GEN_15910 ? phv_data_411 : _GEN_7589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7591 = 9'h19c == _GEN_15910 ? phv_data_412 : _GEN_7590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7592 = 9'h19d == _GEN_15910 ? phv_data_413 : _GEN_7591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7593 = 9'h19e == _GEN_15910 ? phv_data_414 : _GEN_7592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7594 = 9'h19f == _GEN_15910 ? phv_data_415 : _GEN_7593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7595 = 9'h1a0 == _GEN_15910 ? phv_data_416 : _GEN_7594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7596 = 9'h1a1 == _GEN_15910 ? phv_data_417 : _GEN_7595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7597 = 9'h1a2 == _GEN_15910 ? phv_data_418 : _GEN_7596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7598 = 9'h1a3 == _GEN_15910 ? phv_data_419 : _GEN_7597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7599 = 9'h1a4 == _GEN_15910 ? phv_data_420 : _GEN_7598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7600 = 9'h1a5 == _GEN_15910 ? phv_data_421 : _GEN_7599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7601 = 9'h1a6 == _GEN_15910 ? phv_data_422 : _GEN_7600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7602 = 9'h1a7 == _GEN_15910 ? phv_data_423 : _GEN_7601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7603 = 9'h1a8 == _GEN_15910 ? phv_data_424 : _GEN_7602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7604 = 9'h1a9 == _GEN_15910 ? phv_data_425 : _GEN_7603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7605 = 9'h1aa == _GEN_15910 ? phv_data_426 : _GEN_7604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7606 = 9'h1ab == _GEN_15910 ? phv_data_427 : _GEN_7605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7607 = 9'h1ac == _GEN_15910 ? phv_data_428 : _GEN_7606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7608 = 9'h1ad == _GEN_15910 ? phv_data_429 : _GEN_7607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7609 = 9'h1ae == _GEN_15910 ? phv_data_430 : _GEN_7608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7610 = 9'h1af == _GEN_15910 ? phv_data_431 : _GEN_7609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7611 = 9'h1b0 == _GEN_15910 ? phv_data_432 : _GEN_7610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7612 = 9'h1b1 == _GEN_15910 ? phv_data_433 : _GEN_7611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7613 = 9'h1b2 == _GEN_15910 ? phv_data_434 : _GEN_7612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7614 = 9'h1b3 == _GEN_15910 ? phv_data_435 : _GEN_7613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7615 = 9'h1b4 == _GEN_15910 ? phv_data_436 : _GEN_7614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7616 = 9'h1b5 == _GEN_15910 ? phv_data_437 : _GEN_7615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7617 = 9'h1b6 == _GEN_15910 ? phv_data_438 : _GEN_7616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7618 = 9'h1b7 == _GEN_15910 ? phv_data_439 : _GEN_7617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7619 = 9'h1b8 == _GEN_15910 ? phv_data_440 : _GEN_7618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7620 = 9'h1b9 == _GEN_15910 ? phv_data_441 : _GEN_7619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7621 = 9'h1ba == _GEN_15910 ? phv_data_442 : _GEN_7620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7622 = 9'h1bb == _GEN_15910 ? phv_data_443 : _GEN_7621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7623 = 9'h1bc == _GEN_15910 ? phv_data_444 : _GEN_7622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7624 = 9'h1bd == _GEN_15910 ? phv_data_445 : _GEN_7623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7625 = 9'h1be == _GEN_15910 ? phv_data_446 : _GEN_7624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7626 = 9'h1bf == _GEN_15910 ? phv_data_447 : _GEN_7625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7627 = 9'h1c0 == _GEN_15910 ? phv_data_448 : _GEN_7626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7628 = 9'h1c1 == _GEN_15910 ? phv_data_449 : _GEN_7627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7629 = 9'h1c2 == _GEN_15910 ? phv_data_450 : _GEN_7628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7630 = 9'h1c3 == _GEN_15910 ? phv_data_451 : _GEN_7629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7631 = 9'h1c4 == _GEN_15910 ? phv_data_452 : _GEN_7630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7632 = 9'h1c5 == _GEN_15910 ? phv_data_453 : _GEN_7631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7633 = 9'h1c6 == _GEN_15910 ? phv_data_454 : _GEN_7632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7634 = 9'h1c7 == _GEN_15910 ? phv_data_455 : _GEN_7633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7635 = 9'h1c8 == _GEN_15910 ? phv_data_456 : _GEN_7634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7636 = 9'h1c9 == _GEN_15910 ? phv_data_457 : _GEN_7635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7637 = 9'h1ca == _GEN_15910 ? phv_data_458 : _GEN_7636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7638 = 9'h1cb == _GEN_15910 ? phv_data_459 : _GEN_7637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7639 = 9'h1cc == _GEN_15910 ? phv_data_460 : _GEN_7638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7640 = 9'h1cd == _GEN_15910 ? phv_data_461 : _GEN_7639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7641 = 9'h1ce == _GEN_15910 ? phv_data_462 : _GEN_7640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7642 = 9'h1cf == _GEN_15910 ? phv_data_463 : _GEN_7641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7643 = 9'h1d0 == _GEN_15910 ? phv_data_464 : _GEN_7642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7644 = 9'h1d1 == _GEN_15910 ? phv_data_465 : _GEN_7643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7645 = 9'h1d2 == _GEN_15910 ? phv_data_466 : _GEN_7644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7646 = 9'h1d3 == _GEN_15910 ? phv_data_467 : _GEN_7645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7647 = 9'h1d4 == _GEN_15910 ? phv_data_468 : _GEN_7646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7648 = 9'h1d5 == _GEN_15910 ? phv_data_469 : _GEN_7647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7649 = 9'h1d6 == _GEN_15910 ? phv_data_470 : _GEN_7648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7650 = 9'h1d7 == _GEN_15910 ? phv_data_471 : _GEN_7649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7651 = 9'h1d8 == _GEN_15910 ? phv_data_472 : _GEN_7650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7652 = 9'h1d9 == _GEN_15910 ? phv_data_473 : _GEN_7651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7653 = 9'h1da == _GEN_15910 ? phv_data_474 : _GEN_7652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7654 = 9'h1db == _GEN_15910 ? phv_data_475 : _GEN_7653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7655 = 9'h1dc == _GEN_15910 ? phv_data_476 : _GEN_7654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7656 = 9'h1dd == _GEN_15910 ? phv_data_477 : _GEN_7655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7657 = 9'h1de == _GEN_15910 ? phv_data_478 : _GEN_7656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7658 = 9'h1df == _GEN_15910 ? phv_data_479 : _GEN_7657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7659 = 9'h1e0 == _GEN_15910 ? phv_data_480 : _GEN_7658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7660 = 9'h1e1 == _GEN_15910 ? phv_data_481 : _GEN_7659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7661 = 9'h1e2 == _GEN_15910 ? phv_data_482 : _GEN_7660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7662 = 9'h1e3 == _GEN_15910 ? phv_data_483 : _GEN_7661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7663 = 9'h1e4 == _GEN_15910 ? phv_data_484 : _GEN_7662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7664 = 9'h1e5 == _GEN_15910 ? phv_data_485 : _GEN_7663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7665 = 9'h1e6 == _GEN_15910 ? phv_data_486 : _GEN_7664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7666 = 9'h1e7 == _GEN_15910 ? phv_data_487 : _GEN_7665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7667 = 9'h1e8 == _GEN_15910 ? phv_data_488 : _GEN_7666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7668 = 9'h1e9 == _GEN_15910 ? phv_data_489 : _GEN_7667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7669 = 9'h1ea == _GEN_15910 ? phv_data_490 : _GEN_7668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7670 = 9'h1eb == _GEN_15910 ? phv_data_491 : _GEN_7669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7671 = 9'h1ec == _GEN_15910 ? phv_data_492 : _GEN_7670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7672 = 9'h1ed == _GEN_15910 ? phv_data_493 : _GEN_7671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7673 = 9'h1ee == _GEN_15910 ? phv_data_494 : _GEN_7672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7674 = 9'h1ef == _GEN_15910 ? phv_data_495 : _GEN_7673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7675 = 9'h1f0 == _GEN_15910 ? phv_data_496 : _GEN_7674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7676 = 9'h1f1 == _GEN_15910 ? phv_data_497 : _GEN_7675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7677 = 9'h1f2 == _GEN_15910 ? phv_data_498 : _GEN_7676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7678 = 9'h1f3 == _GEN_15910 ? phv_data_499 : _GEN_7677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7679 = 9'h1f4 == _GEN_15910 ? phv_data_500 : _GEN_7678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7680 = 9'h1f5 == _GEN_15910 ? phv_data_501 : _GEN_7679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7681 = 9'h1f6 == _GEN_15910 ? phv_data_502 : _GEN_7680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7682 = 9'h1f7 == _GEN_15910 ? phv_data_503 : _GEN_7681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7683 = 9'h1f8 == _GEN_15910 ? phv_data_504 : _GEN_7682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7684 = 9'h1f9 == _GEN_15910 ? phv_data_505 : _GEN_7683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7685 = 9'h1fa == _GEN_15910 ? phv_data_506 : _GEN_7684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7686 = 9'h1fb == _GEN_15910 ? phv_data_507 : _GEN_7685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7687 = 9'h1fc == _GEN_15910 ? phv_data_508 : _GEN_7686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7688 = 9'h1fd == _GEN_15910 ? phv_data_509 : _GEN_7687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7689 = 9'h1fe == _GEN_15910 ? phv_data_510 : _GEN_7688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7690 = 9'h1ff == _GEN_15910 ? phv_data_511 : _GEN_7689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7692 = 8'h1 == _match_key_qbytes_3_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7693 = 8'h2 == _match_key_qbytes_3_T_1 ? phv_data_2 : _GEN_7692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7694 = 8'h3 == _match_key_qbytes_3_T_1 ? phv_data_3 : _GEN_7693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7695 = 8'h4 == _match_key_qbytes_3_T_1 ? phv_data_4 : _GEN_7694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7696 = 8'h5 == _match_key_qbytes_3_T_1 ? phv_data_5 : _GEN_7695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7697 = 8'h6 == _match_key_qbytes_3_T_1 ? phv_data_6 : _GEN_7696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7698 = 8'h7 == _match_key_qbytes_3_T_1 ? phv_data_7 : _GEN_7697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7699 = 8'h8 == _match_key_qbytes_3_T_1 ? phv_data_8 : _GEN_7698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7700 = 8'h9 == _match_key_qbytes_3_T_1 ? phv_data_9 : _GEN_7699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7701 = 8'ha == _match_key_qbytes_3_T_1 ? phv_data_10 : _GEN_7700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7702 = 8'hb == _match_key_qbytes_3_T_1 ? phv_data_11 : _GEN_7701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7703 = 8'hc == _match_key_qbytes_3_T_1 ? phv_data_12 : _GEN_7702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7704 = 8'hd == _match_key_qbytes_3_T_1 ? phv_data_13 : _GEN_7703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7705 = 8'he == _match_key_qbytes_3_T_1 ? phv_data_14 : _GEN_7704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7706 = 8'hf == _match_key_qbytes_3_T_1 ? phv_data_15 : _GEN_7705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7707 = 8'h10 == _match_key_qbytes_3_T_1 ? phv_data_16 : _GEN_7706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7708 = 8'h11 == _match_key_qbytes_3_T_1 ? phv_data_17 : _GEN_7707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7709 = 8'h12 == _match_key_qbytes_3_T_1 ? phv_data_18 : _GEN_7708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7710 = 8'h13 == _match_key_qbytes_3_T_1 ? phv_data_19 : _GEN_7709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7711 = 8'h14 == _match_key_qbytes_3_T_1 ? phv_data_20 : _GEN_7710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7712 = 8'h15 == _match_key_qbytes_3_T_1 ? phv_data_21 : _GEN_7711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7713 = 8'h16 == _match_key_qbytes_3_T_1 ? phv_data_22 : _GEN_7712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7714 = 8'h17 == _match_key_qbytes_3_T_1 ? phv_data_23 : _GEN_7713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7715 = 8'h18 == _match_key_qbytes_3_T_1 ? phv_data_24 : _GEN_7714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7716 = 8'h19 == _match_key_qbytes_3_T_1 ? phv_data_25 : _GEN_7715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7717 = 8'h1a == _match_key_qbytes_3_T_1 ? phv_data_26 : _GEN_7716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7718 = 8'h1b == _match_key_qbytes_3_T_1 ? phv_data_27 : _GEN_7717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7719 = 8'h1c == _match_key_qbytes_3_T_1 ? phv_data_28 : _GEN_7718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7720 = 8'h1d == _match_key_qbytes_3_T_1 ? phv_data_29 : _GEN_7719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7721 = 8'h1e == _match_key_qbytes_3_T_1 ? phv_data_30 : _GEN_7720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7722 = 8'h1f == _match_key_qbytes_3_T_1 ? phv_data_31 : _GEN_7721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7723 = 8'h20 == _match_key_qbytes_3_T_1 ? phv_data_32 : _GEN_7722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7724 = 8'h21 == _match_key_qbytes_3_T_1 ? phv_data_33 : _GEN_7723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7725 = 8'h22 == _match_key_qbytes_3_T_1 ? phv_data_34 : _GEN_7724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7726 = 8'h23 == _match_key_qbytes_3_T_1 ? phv_data_35 : _GEN_7725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7727 = 8'h24 == _match_key_qbytes_3_T_1 ? phv_data_36 : _GEN_7726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7728 = 8'h25 == _match_key_qbytes_3_T_1 ? phv_data_37 : _GEN_7727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7729 = 8'h26 == _match_key_qbytes_3_T_1 ? phv_data_38 : _GEN_7728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7730 = 8'h27 == _match_key_qbytes_3_T_1 ? phv_data_39 : _GEN_7729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7731 = 8'h28 == _match_key_qbytes_3_T_1 ? phv_data_40 : _GEN_7730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7732 = 8'h29 == _match_key_qbytes_3_T_1 ? phv_data_41 : _GEN_7731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7733 = 8'h2a == _match_key_qbytes_3_T_1 ? phv_data_42 : _GEN_7732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7734 = 8'h2b == _match_key_qbytes_3_T_1 ? phv_data_43 : _GEN_7733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7735 = 8'h2c == _match_key_qbytes_3_T_1 ? phv_data_44 : _GEN_7734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7736 = 8'h2d == _match_key_qbytes_3_T_1 ? phv_data_45 : _GEN_7735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7737 = 8'h2e == _match_key_qbytes_3_T_1 ? phv_data_46 : _GEN_7736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7738 = 8'h2f == _match_key_qbytes_3_T_1 ? phv_data_47 : _GEN_7737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7739 = 8'h30 == _match_key_qbytes_3_T_1 ? phv_data_48 : _GEN_7738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7740 = 8'h31 == _match_key_qbytes_3_T_1 ? phv_data_49 : _GEN_7739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7741 = 8'h32 == _match_key_qbytes_3_T_1 ? phv_data_50 : _GEN_7740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7742 = 8'h33 == _match_key_qbytes_3_T_1 ? phv_data_51 : _GEN_7741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7743 = 8'h34 == _match_key_qbytes_3_T_1 ? phv_data_52 : _GEN_7742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7744 = 8'h35 == _match_key_qbytes_3_T_1 ? phv_data_53 : _GEN_7743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7745 = 8'h36 == _match_key_qbytes_3_T_1 ? phv_data_54 : _GEN_7744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7746 = 8'h37 == _match_key_qbytes_3_T_1 ? phv_data_55 : _GEN_7745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7747 = 8'h38 == _match_key_qbytes_3_T_1 ? phv_data_56 : _GEN_7746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7748 = 8'h39 == _match_key_qbytes_3_T_1 ? phv_data_57 : _GEN_7747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7749 = 8'h3a == _match_key_qbytes_3_T_1 ? phv_data_58 : _GEN_7748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7750 = 8'h3b == _match_key_qbytes_3_T_1 ? phv_data_59 : _GEN_7749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7751 = 8'h3c == _match_key_qbytes_3_T_1 ? phv_data_60 : _GEN_7750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7752 = 8'h3d == _match_key_qbytes_3_T_1 ? phv_data_61 : _GEN_7751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7753 = 8'h3e == _match_key_qbytes_3_T_1 ? phv_data_62 : _GEN_7752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7754 = 8'h3f == _match_key_qbytes_3_T_1 ? phv_data_63 : _GEN_7753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7755 = 8'h40 == _match_key_qbytes_3_T_1 ? phv_data_64 : _GEN_7754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7756 = 8'h41 == _match_key_qbytes_3_T_1 ? phv_data_65 : _GEN_7755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7757 = 8'h42 == _match_key_qbytes_3_T_1 ? phv_data_66 : _GEN_7756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7758 = 8'h43 == _match_key_qbytes_3_T_1 ? phv_data_67 : _GEN_7757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7759 = 8'h44 == _match_key_qbytes_3_T_1 ? phv_data_68 : _GEN_7758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7760 = 8'h45 == _match_key_qbytes_3_T_1 ? phv_data_69 : _GEN_7759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7761 = 8'h46 == _match_key_qbytes_3_T_1 ? phv_data_70 : _GEN_7760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7762 = 8'h47 == _match_key_qbytes_3_T_1 ? phv_data_71 : _GEN_7761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7763 = 8'h48 == _match_key_qbytes_3_T_1 ? phv_data_72 : _GEN_7762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7764 = 8'h49 == _match_key_qbytes_3_T_1 ? phv_data_73 : _GEN_7763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7765 = 8'h4a == _match_key_qbytes_3_T_1 ? phv_data_74 : _GEN_7764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7766 = 8'h4b == _match_key_qbytes_3_T_1 ? phv_data_75 : _GEN_7765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7767 = 8'h4c == _match_key_qbytes_3_T_1 ? phv_data_76 : _GEN_7766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7768 = 8'h4d == _match_key_qbytes_3_T_1 ? phv_data_77 : _GEN_7767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7769 = 8'h4e == _match_key_qbytes_3_T_1 ? phv_data_78 : _GEN_7768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7770 = 8'h4f == _match_key_qbytes_3_T_1 ? phv_data_79 : _GEN_7769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7771 = 8'h50 == _match_key_qbytes_3_T_1 ? phv_data_80 : _GEN_7770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7772 = 8'h51 == _match_key_qbytes_3_T_1 ? phv_data_81 : _GEN_7771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7773 = 8'h52 == _match_key_qbytes_3_T_1 ? phv_data_82 : _GEN_7772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7774 = 8'h53 == _match_key_qbytes_3_T_1 ? phv_data_83 : _GEN_7773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7775 = 8'h54 == _match_key_qbytes_3_T_1 ? phv_data_84 : _GEN_7774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7776 = 8'h55 == _match_key_qbytes_3_T_1 ? phv_data_85 : _GEN_7775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7777 = 8'h56 == _match_key_qbytes_3_T_1 ? phv_data_86 : _GEN_7776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7778 = 8'h57 == _match_key_qbytes_3_T_1 ? phv_data_87 : _GEN_7777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7779 = 8'h58 == _match_key_qbytes_3_T_1 ? phv_data_88 : _GEN_7778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7780 = 8'h59 == _match_key_qbytes_3_T_1 ? phv_data_89 : _GEN_7779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7781 = 8'h5a == _match_key_qbytes_3_T_1 ? phv_data_90 : _GEN_7780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7782 = 8'h5b == _match_key_qbytes_3_T_1 ? phv_data_91 : _GEN_7781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7783 = 8'h5c == _match_key_qbytes_3_T_1 ? phv_data_92 : _GEN_7782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7784 = 8'h5d == _match_key_qbytes_3_T_1 ? phv_data_93 : _GEN_7783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7785 = 8'h5e == _match_key_qbytes_3_T_1 ? phv_data_94 : _GEN_7784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7786 = 8'h5f == _match_key_qbytes_3_T_1 ? phv_data_95 : _GEN_7785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7787 = 8'h60 == _match_key_qbytes_3_T_1 ? phv_data_96 : _GEN_7786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7788 = 8'h61 == _match_key_qbytes_3_T_1 ? phv_data_97 : _GEN_7787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7789 = 8'h62 == _match_key_qbytes_3_T_1 ? phv_data_98 : _GEN_7788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7790 = 8'h63 == _match_key_qbytes_3_T_1 ? phv_data_99 : _GEN_7789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7791 = 8'h64 == _match_key_qbytes_3_T_1 ? phv_data_100 : _GEN_7790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7792 = 8'h65 == _match_key_qbytes_3_T_1 ? phv_data_101 : _GEN_7791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7793 = 8'h66 == _match_key_qbytes_3_T_1 ? phv_data_102 : _GEN_7792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7794 = 8'h67 == _match_key_qbytes_3_T_1 ? phv_data_103 : _GEN_7793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7795 = 8'h68 == _match_key_qbytes_3_T_1 ? phv_data_104 : _GEN_7794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7796 = 8'h69 == _match_key_qbytes_3_T_1 ? phv_data_105 : _GEN_7795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7797 = 8'h6a == _match_key_qbytes_3_T_1 ? phv_data_106 : _GEN_7796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7798 = 8'h6b == _match_key_qbytes_3_T_1 ? phv_data_107 : _GEN_7797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7799 = 8'h6c == _match_key_qbytes_3_T_1 ? phv_data_108 : _GEN_7798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7800 = 8'h6d == _match_key_qbytes_3_T_1 ? phv_data_109 : _GEN_7799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7801 = 8'h6e == _match_key_qbytes_3_T_1 ? phv_data_110 : _GEN_7800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7802 = 8'h6f == _match_key_qbytes_3_T_1 ? phv_data_111 : _GEN_7801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7803 = 8'h70 == _match_key_qbytes_3_T_1 ? phv_data_112 : _GEN_7802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7804 = 8'h71 == _match_key_qbytes_3_T_1 ? phv_data_113 : _GEN_7803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7805 = 8'h72 == _match_key_qbytes_3_T_1 ? phv_data_114 : _GEN_7804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7806 = 8'h73 == _match_key_qbytes_3_T_1 ? phv_data_115 : _GEN_7805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7807 = 8'h74 == _match_key_qbytes_3_T_1 ? phv_data_116 : _GEN_7806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7808 = 8'h75 == _match_key_qbytes_3_T_1 ? phv_data_117 : _GEN_7807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7809 = 8'h76 == _match_key_qbytes_3_T_1 ? phv_data_118 : _GEN_7808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7810 = 8'h77 == _match_key_qbytes_3_T_1 ? phv_data_119 : _GEN_7809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7811 = 8'h78 == _match_key_qbytes_3_T_1 ? phv_data_120 : _GEN_7810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7812 = 8'h79 == _match_key_qbytes_3_T_1 ? phv_data_121 : _GEN_7811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7813 = 8'h7a == _match_key_qbytes_3_T_1 ? phv_data_122 : _GEN_7812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7814 = 8'h7b == _match_key_qbytes_3_T_1 ? phv_data_123 : _GEN_7813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7815 = 8'h7c == _match_key_qbytes_3_T_1 ? phv_data_124 : _GEN_7814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7816 = 8'h7d == _match_key_qbytes_3_T_1 ? phv_data_125 : _GEN_7815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7817 = 8'h7e == _match_key_qbytes_3_T_1 ? phv_data_126 : _GEN_7816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7818 = 8'h7f == _match_key_qbytes_3_T_1 ? phv_data_127 : _GEN_7817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7819 = 8'h80 == _match_key_qbytes_3_T_1 ? phv_data_128 : _GEN_7818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7820 = 8'h81 == _match_key_qbytes_3_T_1 ? phv_data_129 : _GEN_7819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7821 = 8'h82 == _match_key_qbytes_3_T_1 ? phv_data_130 : _GEN_7820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7822 = 8'h83 == _match_key_qbytes_3_T_1 ? phv_data_131 : _GEN_7821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7823 = 8'h84 == _match_key_qbytes_3_T_1 ? phv_data_132 : _GEN_7822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7824 = 8'h85 == _match_key_qbytes_3_T_1 ? phv_data_133 : _GEN_7823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7825 = 8'h86 == _match_key_qbytes_3_T_1 ? phv_data_134 : _GEN_7824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7826 = 8'h87 == _match_key_qbytes_3_T_1 ? phv_data_135 : _GEN_7825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7827 = 8'h88 == _match_key_qbytes_3_T_1 ? phv_data_136 : _GEN_7826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7828 = 8'h89 == _match_key_qbytes_3_T_1 ? phv_data_137 : _GEN_7827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7829 = 8'h8a == _match_key_qbytes_3_T_1 ? phv_data_138 : _GEN_7828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7830 = 8'h8b == _match_key_qbytes_3_T_1 ? phv_data_139 : _GEN_7829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7831 = 8'h8c == _match_key_qbytes_3_T_1 ? phv_data_140 : _GEN_7830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7832 = 8'h8d == _match_key_qbytes_3_T_1 ? phv_data_141 : _GEN_7831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7833 = 8'h8e == _match_key_qbytes_3_T_1 ? phv_data_142 : _GEN_7832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7834 = 8'h8f == _match_key_qbytes_3_T_1 ? phv_data_143 : _GEN_7833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7835 = 8'h90 == _match_key_qbytes_3_T_1 ? phv_data_144 : _GEN_7834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7836 = 8'h91 == _match_key_qbytes_3_T_1 ? phv_data_145 : _GEN_7835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7837 = 8'h92 == _match_key_qbytes_3_T_1 ? phv_data_146 : _GEN_7836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7838 = 8'h93 == _match_key_qbytes_3_T_1 ? phv_data_147 : _GEN_7837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7839 = 8'h94 == _match_key_qbytes_3_T_1 ? phv_data_148 : _GEN_7838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7840 = 8'h95 == _match_key_qbytes_3_T_1 ? phv_data_149 : _GEN_7839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7841 = 8'h96 == _match_key_qbytes_3_T_1 ? phv_data_150 : _GEN_7840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7842 = 8'h97 == _match_key_qbytes_3_T_1 ? phv_data_151 : _GEN_7841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7843 = 8'h98 == _match_key_qbytes_3_T_1 ? phv_data_152 : _GEN_7842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7844 = 8'h99 == _match_key_qbytes_3_T_1 ? phv_data_153 : _GEN_7843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7845 = 8'h9a == _match_key_qbytes_3_T_1 ? phv_data_154 : _GEN_7844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7846 = 8'h9b == _match_key_qbytes_3_T_1 ? phv_data_155 : _GEN_7845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7847 = 8'h9c == _match_key_qbytes_3_T_1 ? phv_data_156 : _GEN_7846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7848 = 8'h9d == _match_key_qbytes_3_T_1 ? phv_data_157 : _GEN_7847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7849 = 8'h9e == _match_key_qbytes_3_T_1 ? phv_data_158 : _GEN_7848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7850 = 8'h9f == _match_key_qbytes_3_T_1 ? phv_data_159 : _GEN_7849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7851 = 8'ha0 == _match_key_qbytes_3_T_1 ? phv_data_160 : _GEN_7850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7852 = 8'ha1 == _match_key_qbytes_3_T_1 ? phv_data_161 : _GEN_7851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7853 = 8'ha2 == _match_key_qbytes_3_T_1 ? phv_data_162 : _GEN_7852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7854 = 8'ha3 == _match_key_qbytes_3_T_1 ? phv_data_163 : _GEN_7853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7855 = 8'ha4 == _match_key_qbytes_3_T_1 ? phv_data_164 : _GEN_7854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7856 = 8'ha5 == _match_key_qbytes_3_T_1 ? phv_data_165 : _GEN_7855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7857 = 8'ha6 == _match_key_qbytes_3_T_1 ? phv_data_166 : _GEN_7856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7858 = 8'ha7 == _match_key_qbytes_3_T_1 ? phv_data_167 : _GEN_7857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7859 = 8'ha8 == _match_key_qbytes_3_T_1 ? phv_data_168 : _GEN_7858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7860 = 8'ha9 == _match_key_qbytes_3_T_1 ? phv_data_169 : _GEN_7859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7861 = 8'haa == _match_key_qbytes_3_T_1 ? phv_data_170 : _GEN_7860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7862 = 8'hab == _match_key_qbytes_3_T_1 ? phv_data_171 : _GEN_7861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7863 = 8'hac == _match_key_qbytes_3_T_1 ? phv_data_172 : _GEN_7862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7864 = 8'had == _match_key_qbytes_3_T_1 ? phv_data_173 : _GEN_7863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7865 = 8'hae == _match_key_qbytes_3_T_1 ? phv_data_174 : _GEN_7864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7866 = 8'haf == _match_key_qbytes_3_T_1 ? phv_data_175 : _GEN_7865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7867 = 8'hb0 == _match_key_qbytes_3_T_1 ? phv_data_176 : _GEN_7866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7868 = 8'hb1 == _match_key_qbytes_3_T_1 ? phv_data_177 : _GEN_7867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7869 = 8'hb2 == _match_key_qbytes_3_T_1 ? phv_data_178 : _GEN_7868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7870 = 8'hb3 == _match_key_qbytes_3_T_1 ? phv_data_179 : _GEN_7869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7871 = 8'hb4 == _match_key_qbytes_3_T_1 ? phv_data_180 : _GEN_7870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7872 = 8'hb5 == _match_key_qbytes_3_T_1 ? phv_data_181 : _GEN_7871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7873 = 8'hb6 == _match_key_qbytes_3_T_1 ? phv_data_182 : _GEN_7872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7874 = 8'hb7 == _match_key_qbytes_3_T_1 ? phv_data_183 : _GEN_7873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7875 = 8'hb8 == _match_key_qbytes_3_T_1 ? phv_data_184 : _GEN_7874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7876 = 8'hb9 == _match_key_qbytes_3_T_1 ? phv_data_185 : _GEN_7875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7877 = 8'hba == _match_key_qbytes_3_T_1 ? phv_data_186 : _GEN_7876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7878 = 8'hbb == _match_key_qbytes_3_T_1 ? phv_data_187 : _GEN_7877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7879 = 8'hbc == _match_key_qbytes_3_T_1 ? phv_data_188 : _GEN_7878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7880 = 8'hbd == _match_key_qbytes_3_T_1 ? phv_data_189 : _GEN_7879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7881 = 8'hbe == _match_key_qbytes_3_T_1 ? phv_data_190 : _GEN_7880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7882 = 8'hbf == _match_key_qbytes_3_T_1 ? phv_data_191 : _GEN_7881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7883 = 8'hc0 == _match_key_qbytes_3_T_1 ? phv_data_192 : _GEN_7882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7884 = 8'hc1 == _match_key_qbytes_3_T_1 ? phv_data_193 : _GEN_7883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7885 = 8'hc2 == _match_key_qbytes_3_T_1 ? phv_data_194 : _GEN_7884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7886 = 8'hc3 == _match_key_qbytes_3_T_1 ? phv_data_195 : _GEN_7885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7887 = 8'hc4 == _match_key_qbytes_3_T_1 ? phv_data_196 : _GEN_7886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7888 = 8'hc5 == _match_key_qbytes_3_T_1 ? phv_data_197 : _GEN_7887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7889 = 8'hc6 == _match_key_qbytes_3_T_1 ? phv_data_198 : _GEN_7888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7890 = 8'hc7 == _match_key_qbytes_3_T_1 ? phv_data_199 : _GEN_7889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7891 = 8'hc8 == _match_key_qbytes_3_T_1 ? phv_data_200 : _GEN_7890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7892 = 8'hc9 == _match_key_qbytes_3_T_1 ? phv_data_201 : _GEN_7891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7893 = 8'hca == _match_key_qbytes_3_T_1 ? phv_data_202 : _GEN_7892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7894 = 8'hcb == _match_key_qbytes_3_T_1 ? phv_data_203 : _GEN_7893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7895 = 8'hcc == _match_key_qbytes_3_T_1 ? phv_data_204 : _GEN_7894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7896 = 8'hcd == _match_key_qbytes_3_T_1 ? phv_data_205 : _GEN_7895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7897 = 8'hce == _match_key_qbytes_3_T_1 ? phv_data_206 : _GEN_7896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7898 = 8'hcf == _match_key_qbytes_3_T_1 ? phv_data_207 : _GEN_7897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7899 = 8'hd0 == _match_key_qbytes_3_T_1 ? phv_data_208 : _GEN_7898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7900 = 8'hd1 == _match_key_qbytes_3_T_1 ? phv_data_209 : _GEN_7899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7901 = 8'hd2 == _match_key_qbytes_3_T_1 ? phv_data_210 : _GEN_7900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7902 = 8'hd3 == _match_key_qbytes_3_T_1 ? phv_data_211 : _GEN_7901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7903 = 8'hd4 == _match_key_qbytes_3_T_1 ? phv_data_212 : _GEN_7902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7904 = 8'hd5 == _match_key_qbytes_3_T_1 ? phv_data_213 : _GEN_7903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7905 = 8'hd6 == _match_key_qbytes_3_T_1 ? phv_data_214 : _GEN_7904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7906 = 8'hd7 == _match_key_qbytes_3_T_1 ? phv_data_215 : _GEN_7905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7907 = 8'hd8 == _match_key_qbytes_3_T_1 ? phv_data_216 : _GEN_7906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7908 = 8'hd9 == _match_key_qbytes_3_T_1 ? phv_data_217 : _GEN_7907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7909 = 8'hda == _match_key_qbytes_3_T_1 ? phv_data_218 : _GEN_7908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7910 = 8'hdb == _match_key_qbytes_3_T_1 ? phv_data_219 : _GEN_7909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7911 = 8'hdc == _match_key_qbytes_3_T_1 ? phv_data_220 : _GEN_7910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7912 = 8'hdd == _match_key_qbytes_3_T_1 ? phv_data_221 : _GEN_7911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7913 = 8'hde == _match_key_qbytes_3_T_1 ? phv_data_222 : _GEN_7912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7914 = 8'hdf == _match_key_qbytes_3_T_1 ? phv_data_223 : _GEN_7913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7915 = 8'he0 == _match_key_qbytes_3_T_1 ? phv_data_224 : _GEN_7914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7916 = 8'he1 == _match_key_qbytes_3_T_1 ? phv_data_225 : _GEN_7915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7917 = 8'he2 == _match_key_qbytes_3_T_1 ? phv_data_226 : _GEN_7916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7918 = 8'he3 == _match_key_qbytes_3_T_1 ? phv_data_227 : _GEN_7917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7919 = 8'he4 == _match_key_qbytes_3_T_1 ? phv_data_228 : _GEN_7918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7920 = 8'he5 == _match_key_qbytes_3_T_1 ? phv_data_229 : _GEN_7919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7921 = 8'he6 == _match_key_qbytes_3_T_1 ? phv_data_230 : _GEN_7920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7922 = 8'he7 == _match_key_qbytes_3_T_1 ? phv_data_231 : _GEN_7921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7923 = 8'he8 == _match_key_qbytes_3_T_1 ? phv_data_232 : _GEN_7922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7924 = 8'he9 == _match_key_qbytes_3_T_1 ? phv_data_233 : _GEN_7923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7925 = 8'hea == _match_key_qbytes_3_T_1 ? phv_data_234 : _GEN_7924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7926 = 8'heb == _match_key_qbytes_3_T_1 ? phv_data_235 : _GEN_7925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7927 = 8'hec == _match_key_qbytes_3_T_1 ? phv_data_236 : _GEN_7926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7928 = 8'hed == _match_key_qbytes_3_T_1 ? phv_data_237 : _GEN_7927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7929 = 8'hee == _match_key_qbytes_3_T_1 ? phv_data_238 : _GEN_7928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7930 = 8'hef == _match_key_qbytes_3_T_1 ? phv_data_239 : _GEN_7929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7931 = 8'hf0 == _match_key_qbytes_3_T_1 ? phv_data_240 : _GEN_7930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7932 = 8'hf1 == _match_key_qbytes_3_T_1 ? phv_data_241 : _GEN_7931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7933 = 8'hf2 == _match_key_qbytes_3_T_1 ? phv_data_242 : _GEN_7932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7934 = 8'hf3 == _match_key_qbytes_3_T_1 ? phv_data_243 : _GEN_7933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7935 = 8'hf4 == _match_key_qbytes_3_T_1 ? phv_data_244 : _GEN_7934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7936 = 8'hf5 == _match_key_qbytes_3_T_1 ? phv_data_245 : _GEN_7935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7937 = 8'hf6 == _match_key_qbytes_3_T_1 ? phv_data_246 : _GEN_7936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7938 = 8'hf7 == _match_key_qbytes_3_T_1 ? phv_data_247 : _GEN_7937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7939 = 8'hf8 == _match_key_qbytes_3_T_1 ? phv_data_248 : _GEN_7938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7940 = 8'hf9 == _match_key_qbytes_3_T_1 ? phv_data_249 : _GEN_7939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7941 = 8'hfa == _match_key_qbytes_3_T_1 ? phv_data_250 : _GEN_7940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7942 = 8'hfb == _match_key_qbytes_3_T_1 ? phv_data_251 : _GEN_7941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7943 = 8'hfc == _match_key_qbytes_3_T_1 ? phv_data_252 : _GEN_7942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7944 = 8'hfd == _match_key_qbytes_3_T_1 ? phv_data_253 : _GEN_7943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7945 = 8'hfe == _match_key_qbytes_3_T_1 ? phv_data_254 : _GEN_7944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7946 = 8'hff == _match_key_qbytes_3_T_1 ? phv_data_255 : _GEN_7945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_16166 = {{1'd0}, _match_key_qbytes_3_T_1}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7947 = 9'h100 == _GEN_16166 ? phv_data_256 : _GEN_7946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7948 = 9'h101 == _GEN_16166 ? phv_data_257 : _GEN_7947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7949 = 9'h102 == _GEN_16166 ? phv_data_258 : _GEN_7948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7950 = 9'h103 == _GEN_16166 ? phv_data_259 : _GEN_7949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7951 = 9'h104 == _GEN_16166 ? phv_data_260 : _GEN_7950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7952 = 9'h105 == _GEN_16166 ? phv_data_261 : _GEN_7951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7953 = 9'h106 == _GEN_16166 ? phv_data_262 : _GEN_7952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7954 = 9'h107 == _GEN_16166 ? phv_data_263 : _GEN_7953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7955 = 9'h108 == _GEN_16166 ? phv_data_264 : _GEN_7954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7956 = 9'h109 == _GEN_16166 ? phv_data_265 : _GEN_7955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7957 = 9'h10a == _GEN_16166 ? phv_data_266 : _GEN_7956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7958 = 9'h10b == _GEN_16166 ? phv_data_267 : _GEN_7957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7959 = 9'h10c == _GEN_16166 ? phv_data_268 : _GEN_7958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7960 = 9'h10d == _GEN_16166 ? phv_data_269 : _GEN_7959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7961 = 9'h10e == _GEN_16166 ? phv_data_270 : _GEN_7960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7962 = 9'h10f == _GEN_16166 ? phv_data_271 : _GEN_7961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7963 = 9'h110 == _GEN_16166 ? phv_data_272 : _GEN_7962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7964 = 9'h111 == _GEN_16166 ? phv_data_273 : _GEN_7963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7965 = 9'h112 == _GEN_16166 ? phv_data_274 : _GEN_7964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7966 = 9'h113 == _GEN_16166 ? phv_data_275 : _GEN_7965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7967 = 9'h114 == _GEN_16166 ? phv_data_276 : _GEN_7966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7968 = 9'h115 == _GEN_16166 ? phv_data_277 : _GEN_7967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7969 = 9'h116 == _GEN_16166 ? phv_data_278 : _GEN_7968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7970 = 9'h117 == _GEN_16166 ? phv_data_279 : _GEN_7969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7971 = 9'h118 == _GEN_16166 ? phv_data_280 : _GEN_7970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7972 = 9'h119 == _GEN_16166 ? phv_data_281 : _GEN_7971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7973 = 9'h11a == _GEN_16166 ? phv_data_282 : _GEN_7972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7974 = 9'h11b == _GEN_16166 ? phv_data_283 : _GEN_7973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7975 = 9'h11c == _GEN_16166 ? phv_data_284 : _GEN_7974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7976 = 9'h11d == _GEN_16166 ? phv_data_285 : _GEN_7975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7977 = 9'h11e == _GEN_16166 ? phv_data_286 : _GEN_7976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7978 = 9'h11f == _GEN_16166 ? phv_data_287 : _GEN_7977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7979 = 9'h120 == _GEN_16166 ? phv_data_288 : _GEN_7978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7980 = 9'h121 == _GEN_16166 ? phv_data_289 : _GEN_7979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7981 = 9'h122 == _GEN_16166 ? phv_data_290 : _GEN_7980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7982 = 9'h123 == _GEN_16166 ? phv_data_291 : _GEN_7981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7983 = 9'h124 == _GEN_16166 ? phv_data_292 : _GEN_7982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7984 = 9'h125 == _GEN_16166 ? phv_data_293 : _GEN_7983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7985 = 9'h126 == _GEN_16166 ? phv_data_294 : _GEN_7984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7986 = 9'h127 == _GEN_16166 ? phv_data_295 : _GEN_7985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7987 = 9'h128 == _GEN_16166 ? phv_data_296 : _GEN_7986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7988 = 9'h129 == _GEN_16166 ? phv_data_297 : _GEN_7987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7989 = 9'h12a == _GEN_16166 ? phv_data_298 : _GEN_7988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7990 = 9'h12b == _GEN_16166 ? phv_data_299 : _GEN_7989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7991 = 9'h12c == _GEN_16166 ? phv_data_300 : _GEN_7990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7992 = 9'h12d == _GEN_16166 ? phv_data_301 : _GEN_7991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7993 = 9'h12e == _GEN_16166 ? phv_data_302 : _GEN_7992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7994 = 9'h12f == _GEN_16166 ? phv_data_303 : _GEN_7993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7995 = 9'h130 == _GEN_16166 ? phv_data_304 : _GEN_7994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7996 = 9'h131 == _GEN_16166 ? phv_data_305 : _GEN_7995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7997 = 9'h132 == _GEN_16166 ? phv_data_306 : _GEN_7996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7998 = 9'h133 == _GEN_16166 ? phv_data_307 : _GEN_7997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7999 = 9'h134 == _GEN_16166 ? phv_data_308 : _GEN_7998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8000 = 9'h135 == _GEN_16166 ? phv_data_309 : _GEN_7999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8001 = 9'h136 == _GEN_16166 ? phv_data_310 : _GEN_8000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8002 = 9'h137 == _GEN_16166 ? phv_data_311 : _GEN_8001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8003 = 9'h138 == _GEN_16166 ? phv_data_312 : _GEN_8002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8004 = 9'h139 == _GEN_16166 ? phv_data_313 : _GEN_8003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8005 = 9'h13a == _GEN_16166 ? phv_data_314 : _GEN_8004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8006 = 9'h13b == _GEN_16166 ? phv_data_315 : _GEN_8005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8007 = 9'h13c == _GEN_16166 ? phv_data_316 : _GEN_8006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8008 = 9'h13d == _GEN_16166 ? phv_data_317 : _GEN_8007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8009 = 9'h13e == _GEN_16166 ? phv_data_318 : _GEN_8008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8010 = 9'h13f == _GEN_16166 ? phv_data_319 : _GEN_8009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8011 = 9'h140 == _GEN_16166 ? phv_data_320 : _GEN_8010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8012 = 9'h141 == _GEN_16166 ? phv_data_321 : _GEN_8011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8013 = 9'h142 == _GEN_16166 ? phv_data_322 : _GEN_8012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8014 = 9'h143 == _GEN_16166 ? phv_data_323 : _GEN_8013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8015 = 9'h144 == _GEN_16166 ? phv_data_324 : _GEN_8014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8016 = 9'h145 == _GEN_16166 ? phv_data_325 : _GEN_8015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8017 = 9'h146 == _GEN_16166 ? phv_data_326 : _GEN_8016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8018 = 9'h147 == _GEN_16166 ? phv_data_327 : _GEN_8017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8019 = 9'h148 == _GEN_16166 ? phv_data_328 : _GEN_8018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8020 = 9'h149 == _GEN_16166 ? phv_data_329 : _GEN_8019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8021 = 9'h14a == _GEN_16166 ? phv_data_330 : _GEN_8020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8022 = 9'h14b == _GEN_16166 ? phv_data_331 : _GEN_8021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8023 = 9'h14c == _GEN_16166 ? phv_data_332 : _GEN_8022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8024 = 9'h14d == _GEN_16166 ? phv_data_333 : _GEN_8023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8025 = 9'h14e == _GEN_16166 ? phv_data_334 : _GEN_8024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8026 = 9'h14f == _GEN_16166 ? phv_data_335 : _GEN_8025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8027 = 9'h150 == _GEN_16166 ? phv_data_336 : _GEN_8026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8028 = 9'h151 == _GEN_16166 ? phv_data_337 : _GEN_8027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8029 = 9'h152 == _GEN_16166 ? phv_data_338 : _GEN_8028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8030 = 9'h153 == _GEN_16166 ? phv_data_339 : _GEN_8029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8031 = 9'h154 == _GEN_16166 ? phv_data_340 : _GEN_8030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8032 = 9'h155 == _GEN_16166 ? phv_data_341 : _GEN_8031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8033 = 9'h156 == _GEN_16166 ? phv_data_342 : _GEN_8032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8034 = 9'h157 == _GEN_16166 ? phv_data_343 : _GEN_8033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8035 = 9'h158 == _GEN_16166 ? phv_data_344 : _GEN_8034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8036 = 9'h159 == _GEN_16166 ? phv_data_345 : _GEN_8035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8037 = 9'h15a == _GEN_16166 ? phv_data_346 : _GEN_8036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8038 = 9'h15b == _GEN_16166 ? phv_data_347 : _GEN_8037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8039 = 9'h15c == _GEN_16166 ? phv_data_348 : _GEN_8038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8040 = 9'h15d == _GEN_16166 ? phv_data_349 : _GEN_8039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8041 = 9'h15e == _GEN_16166 ? phv_data_350 : _GEN_8040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8042 = 9'h15f == _GEN_16166 ? phv_data_351 : _GEN_8041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8043 = 9'h160 == _GEN_16166 ? phv_data_352 : _GEN_8042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8044 = 9'h161 == _GEN_16166 ? phv_data_353 : _GEN_8043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8045 = 9'h162 == _GEN_16166 ? phv_data_354 : _GEN_8044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8046 = 9'h163 == _GEN_16166 ? phv_data_355 : _GEN_8045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8047 = 9'h164 == _GEN_16166 ? phv_data_356 : _GEN_8046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8048 = 9'h165 == _GEN_16166 ? phv_data_357 : _GEN_8047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8049 = 9'h166 == _GEN_16166 ? phv_data_358 : _GEN_8048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8050 = 9'h167 == _GEN_16166 ? phv_data_359 : _GEN_8049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8051 = 9'h168 == _GEN_16166 ? phv_data_360 : _GEN_8050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8052 = 9'h169 == _GEN_16166 ? phv_data_361 : _GEN_8051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8053 = 9'h16a == _GEN_16166 ? phv_data_362 : _GEN_8052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8054 = 9'h16b == _GEN_16166 ? phv_data_363 : _GEN_8053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8055 = 9'h16c == _GEN_16166 ? phv_data_364 : _GEN_8054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8056 = 9'h16d == _GEN_16166 ? phv_data_365 : _GEN_8055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8057 = 9'h16e == _GEN_16166 ? phv_data_366 : _GEN_8056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8058 = 9'h16f == _GEN_16166 ? phv_data_367 : _GEN_8057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8059 = 9'h170 == _GEN_16166 ? phv_data_368 : _GEN_8058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8060 = 9'h171 == _GEN_16166 ? phv_data_369 : _GEN_8059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8061 = 9'h172 == _GEN_16166 ? phv_data_370 : _GEN_8060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8062 = 9'h173 == _GEN_16166 ? phv_data_371 : _GEN_8061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8063 = 9'h174 == _GEN_16166 ? phv_data_372 : _GEN_8062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8064 = 9'h175 == _GEN_16166 ? phv_data_373 : _GEN_8063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8065 = 9'h176 == _GEN_16166 ? phv_data_374 : _GEN_8064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8066 = 9'h177 == _GEN_16166 ? phv_data_375 : _GEN_8065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8067 = 9'h178 == _GEN_16166 ? phv_data_376 : _GEN_8066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8068 = 9'h179 == _GEN_16166 ? phv_data_377 : _GEN_8067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8069 = 9'h17a == _GEN_16166 ? phv_data_378 : _GEN_8068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8070 = 9'h17b == _GEN_16166 ? phv_data_379 : _GEN_8069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8071 = 9'h17c == _GEN_16166 ? phv_data_380 : _GEN_8070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8072 = 9'h17d == _GEN_16166 ? phv_data_381 : _GEN_8071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8073 = 9'h17e == _GEN_16166 ? phv_data_382 : _GEN_8072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8074 = 9'h17f == _GEN_16166 ? phv_data_383 : _GEN_8073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8075 = 9'h180 == _GEN_16166 ? phv_data_384 : _GEN_8074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8076 = 9'h181 == _GEN_16166 ? phv_data_385 : _GEN_8075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8077 = 9'h182 == _GEN_16166 ? phv_data_386 : _GEN_8076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8078 = 9'h183 == _GEN_16166 ? phv_data_387 : _GEN_8077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8079 = 9'h184 == _GEN_16166 ? phv_data_388 : _GEN_8078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8080 = 9'h185 == _GEN_16166 ? phv_data_389 : _GEN_8079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8081 = 9'h186 == _GEN_16166 ? phv_data_390 : _GEN_8080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8082 = 9'h187 == _GEN_16166 ? phv_data_391 : _GEN_8081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8083 = 9'h188 == _GEN_16166 ? phv_data_392 : _GEN_8082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8084 = 9'h189 == _GEN_16166 ? phv_data_393 : _GEN_8083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8085 = 9'h18a == _GEN_16166 ? phv_data_394 : _GEN_8084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8086 = 9'h18b == _GEN_16166 ? phv_data_395 : _GEN_8085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8087 = 9'h18c == _GEN_16166 ? phv_data_396 : _GEN_8086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8088 = 9'h18d == _GEN_16166 ? phv_data_397 : _GEN_8087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8089 = 9'h18e == _GEN_16166 ? phv_data_398 : _GEN_8088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8090 = 9'h18f == _GEN_16166 ? phv_data_399 : _GEN_8089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8091 = 9'h190 == _GEN_16166 ? phv_data_400 : _GEN_8090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8092 = 9'h191 == _GEN_16166 ? phv_data_401 : _GEN_8091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8093 = 9'h192 == _GEN_16166 ? phv_data_402 : _GEN_8092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8094 = 9'h193 == _GEN_16166 ? phv_data_403 : _GEN_8093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8095 = 9'h194 == _GEN_16166 ? phv_data_404 : _GEN_8094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8096 = 9'h195 == _GEN_16166 ? phv_data_405 : _GEN_8095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8097 = 9'h196 == _GEN_16166 ? phv_data_406 : _GEN_8096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8098 = 9'h197 == _GEN_16166 ? phv_data_407 : _GEN_8097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8099 = 9'h198 == _GEN_16166 ? phv_data_408 : _GEN_8098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8100 = 9'h199 == _GEN_16166 ? phv_data_409 : _GEN_8099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8101 = 9'h19a == _GEN_16166 ? phv_data_410 : _GEN_8100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8102 = 9'h19b == _GEN_16166 ? phv_data_411 : _GEN_8101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8103 = 9'h19c == _GEN_16166 ? phv_data_412 : _GEN_8102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8104 = 9'h19d == _GEN_16166 ? phv_data_413 : _GEN_8103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8105 = 9'h19e == _GEN_16166 ? phv_data_414 : _GEN_8104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8106 = 9'h19f == _GEN_16166 ? phv_data_415 : _GEN_8105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8107 = 9'h1a0 == _GEN_16166 ? phv_data_416 : _GEN_8106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8108 = 9'h1a1 == _GEN_16166 ? phv_data_417 : _GEN_8107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8109 = 9'h1a2 == _GEN_16166 ? phv_data_418 : _GEN_8108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8110 = 9'h1a3 == _GEN_16166 ? phv_data_419 : _GEN_8109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8111 = 9'h1a4 == _GEN_16166 ? phv_data_420 : _GEN_8110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8112 = 9'h1a5 == _GEN_16166 ? phv_data_421 : _GEN_8111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8113 = 9'h1a6 == _GEN_16166 ? phv_data_422 : _GEN_8112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8114 = 9'h1a7 == _GEN_16166 ? phv_data_423 : _GEN_8113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8115 = 9'h1a8 == _GEN_16166 ? phv_data_424 : _GEN_8114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8116 = 9'h1a9 == _GEN_16166 ? phv_data_425 : _GEN_8115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8117 = 9'h1aa == _GEN_16166 ? phv_data_426 : _GEN_8116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8118 = 9'h1ab == _GEN_16166 ? phv_data_427 : _GEN_8117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8119 = 9'h1ac == _GEN_16166 ? phv_data_428 : _GEN_8118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8120 = 9'h1ad == _GEN_16166 ? phv_data_429 : _GEN_8119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8121 = 9'h1ae == _GEN_16166 ? phv_data_430 : _GEN_8120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8122 = 9'h1af == _GEN_16166 ? phv_data_431 : _GEN_8121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8123 = 9'h1b0 == _GEN_16166 ? phv_data_432 : _GEN_8122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8124 = 9'h1b1 == _GEN_16166 ? phv_data_433 : _GEN_8123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8125 = 9'h1b2 == _GEN_16166 ? phv_data_434 : _GEN_8124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8126 = 9'h1b3 == _GEN_16166 ? phv_data_435 : _GEN_8125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8127 = 9'h1b4 == _GEN_16166 ? phv_data_436 : _GEN_8126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8128 = 9'h1b5 == _GEN_16166 ? phv_data_437 : _GEN_8127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8129 = 9'h1b6 == _GEN_16166 ? phv_data_438 : _GEN_8128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8130 = 9'h1b7 == _GEN_16166 ? phv_data_439 : _GEN_8129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8131 = 9'h1b8 == _GEN_16166 ? phv_data_440 : _GEN_8130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8132 = 9'h1b9 == _GEN_16166 ? phv_data_441 : _GEN_8131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8133 = 9'h1ba == _GEN_16166 ? phv_data_442 : _GEN_8132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8134 = 9'h1bb == _GEN_16166 ? phv_data_443 : _GEN_8133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8135 = 9'h1bc == _GEN_16166 ? phv_data_444 : _GEN_8134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8136 = 9'h1bd == _GEN_16166 ? phv_data_445 : _GEN_8135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8137 = 9'h1be == _GEN_16166 ? phv_data_446 : _GEN_8136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8138 = 9'h1bf == _GEN_16166 ? phv_data_447 : _GEN_8137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8139 = 9'h1c0 == _GEN_16166 ? phv_data_448 : _GEN_8138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8140 = 9'h1c1 == _GEN_16166 ? phv_data_449 : _GEN_8139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8141 = 9'h1c2 == _GEN_16166 ? phv_data_450 : _GEN_8140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8142 = 9'h1c3 == _GEN_16166 ? phv_data_451 : _GEN_8141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8143 = 9'h1c4 == _GEN_16166 ? phv_data_452 : _GEN_8142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8144 = 9'h1c5 == _GEN_16166 ? phv_data_453 : _GEN_8143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8145 = 9'h1c6 == _GEN_16166 ? phv_data_454 : _GEN_8144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8146 = 9'h1c7 == _GEN_16166 ? phv_data_455 : _GEN_8145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8147 = 9'h1c8 == _GEN_16166 ? phv_data_456 : _GEN_8146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8148 = 9'h1c9 == _GEN_16166 ? phv_data_457 : _GEN_8147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8149 = 9'h1ca == _GEN_16166 ? phv_data_458 : _GEN_8148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8150 = 9'h1cb == _GEN_16166 ? phv_data_459 : _GEN_8149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8151 = 9'h1cc == _GEN_16166 ? phv_data_460 : _GEN_8150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8152 = 9'h1cd == _GEN_16166 ? phv_data_461 : _GEN_8151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8153 = 9'h1ce == _GEN_16166 ? phv_data_462 : _GEN_8152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8154 = 9'h1cf == _GEN_16166 ? phv_data_463 : _GEN_8153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8155 = 9'h1d0 == _GEN_16166 ? phv_data_464 : _GEN_8154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8156 = 9'h1d1 == _GEN_16166 ? phv_data_465 : _GEN_8155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8157 = 9'h1d2 == _GEN_16166 ? phv_data_466 : _GEN_8156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8158 = 9'h1d3 == _GEN_16166 ? phv_data_467 : _GEN_8157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8159 = 9'h1d4 == _GEN_16166 ? phv_data_468 : _GEN_8158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8160 = 9'h1d5 == _GEN_16166 ? phv_data_469 : _GEN_8159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8161 = 9'h1d6 == _GEN_16166 ? phv_data_470 : _GEN_8160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8162 = 9'h1d7 == _GEN_16166 ? phv_data_471 : _GEN_8161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8163 = 9'h1d8 == _GEN_16166 ? phv_data_472 : _GEN_8162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8164 = 9'h1d9 == _GEN_16166 ? phv_data_473 : _GEN_8163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8165 = 9'h1da == _GEN_16166 ? phv_data_474 : _GEN_8164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8166 = 9'h1db == _GEN_16166 ? phv_data_475 : _GEN_8165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8167 = 9'h1dc == _GEN_16166 ? phv_data_476 : _GEN_8166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8168 = 9'h1dd == _GEN_16166 ? phv_data_477 : _GEN_8167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8169 = 9'h1de == _GEN_16166 ? phv_data_478 : _GEN_8168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8170 = 9'h1df == _GEN_16166 ? phv_data_479 : _GEN_8169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8171 = 9'h1e0 == _GEN_16166 ? phv_data_480 : _GEN_8170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8172 = 9'h1e1 == _GEN_16166 ? phv_data_481 : _GEN_8171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8173 = 9'h1e2 == _GEN_16166 ? phv_data_482 : _GEN_8172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8174 = 9'h1e3 == _GEN_16166 ? phv_data_483 : _GEN_8173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8175 = 9'h1e4 == _GEN_16166 ? phv_data_484 : _GEN_8174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8176 = 9'h1e5 == _GEN_16166 ? phv_data_485 : _GEN_8175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8177 = 9'h1e6 == _GEN_16166 ? phv_data_486 : _GEN_8176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8178 = 9'h1e7 == _GEN_16166 ? phv_data_487 : _GEN_8177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8179 = 9'h1e8 == _GEN_16166 ? phv_data_488 : _GEN_8178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8180 = 9'h1e9 == _GEN_16166 ? phv_data_489 : _GEN_8179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8181 = 9'h1ea == _GEN_16166 ? phv_data_490 : _GEN_8180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8182 = 9'h1eb == _GEN_16166 ? phv_data_491 : _GEN_8181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8183 = 9'h1ec == _GEN_16166 ? phv_data_492 : _GEN_8182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8184 = 9'h1ed == _GEN_16166 ? phv_data_493 : _GEN_8183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8185 = 9'h1ee == _GEN_16166 ? phv_data_494 : _GEN_8184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8186 = 9'h1ef == _GEN_16166 ? phv_data_495 : _GEN_8185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8187 = 9'h1f0 == _GEN_16166 ? phv_data_496 : _GEN_8186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8188 = 9'h1f1 == _GEN_16166 ? phv_data_497 : _GEN_8187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8189 = 9'h1f2 == _GEN_16166 ? phv_data_498 : _GEN_8188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8190 = 9'h1f3 == _GEN_16166 ? phv_data_499 : _GEN_8189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8191 = 9'h1f4 == _GEN_16166 ? phv_data_500 : _GEN_8190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8192 = 9'h1f5 == _GEN_16166 ? phv_data_501 : _GEN_8191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8193 = 9'h1f6 == _GEN_16166 ? phv_data_502 : _GEN_8192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8194 = 9'h1f7 == _GEN_16166 ? phv_data_503 : _GEN_8193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8195 = 9'h1f8 == _GEN_16166 ? phv_data_504 : _GEN_8194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8196 = 9'h1f9 == _GEN_16166 ? phv_data_505 : _GEN_8195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8197 = 9'h1fa == _GEN_16166 ? phv_data_506 : _GEN_8196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8198 = 9'h1fb == _GEN_16166 ? phv_data_507 : _GEN_8197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8199 = 9'h1fc == _GEN_16166 ? phv_data_508 : _GEN_8198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8200 = 9'h1fd == _GEN_16166 ? phv_data_509 : _GEN_8199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8201 = 9'h1fe == _GEN_16166 ? phv_data_510 : _GEN_8200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8202 = 9'h1ff == _GEN_16166 ? phv_data_511 : _GEN_8201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_3_T_3 = {_GEN_7690,_GEN_8202,_GEN_6666,_GEN_7178}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_3 = local_offset_3 < end_offset ? _match_key_qbytes_3_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_4 = 8'h10 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_4_hi = local_offset_4[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_4_T = {match_key_qbytes_4_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_4_T_1 = {match_key_qbytes_4_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_4_T_2 = {match_key_qbytes_4_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_8205 = 8'h1 == _match_key_qbytes_4_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8206 = 8'h2 == _match_key_qbytes_4_T_2 ? phv_data_2 : _GEN_8205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8207 = 8'h3 == _match_key_qbytes_4_T_2 ? phv_data_3 : _GEN_8206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8208 = 8'h4 == _match_key_qbytes_4_T_2 ? phv_data_4 : _GEN_8207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8209 = 8'h5 == _match_key_qbytes_4_T_2 ? phv_data_5 : _GEN_8208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8210 = 8'h6 == _match_key_qbytes_4_T_2 ? phv_data_6 : _GEN_8209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8211 = 8'h7 == _match_key_qbytes_4_T_2 ? phv_data_7 : _GEN_8210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8212 = 8'h8 == _match_key_qbytes_4_T_2 ? phv_data_8 : _GEN_8211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8213 = 8'h9 == _match_key_qbytes_4_T_2 ? phv_data_9 : _GEN_8212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8214 = 8'ha == _match_key_qbytes_4_T_2 ? phv_data_10 : _GEN_8213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8215 = 8'hb == _match_key_qbytes_4_T_2 ? phv_data_11 : _GEN_8214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8216 = 8'hc == _match_key_qbytes_4_T_2 ? phv_data_12 : _GEN_8215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8217 = 8'hd == _match_key_qbytes_4_T_2 ? phv_data_13 : _GEN_8216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8218 = 8'he == _match_key_qbytes_4_T_2 ? phv_data_14 : _GEN_8217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8219 = 8'hf == _match_key_qbytes_4_T_2 ? phv_data_15 : _GEN_8218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8220 = 8'h10 == _match_key_qbytes_4_T_2 ? phv_data_16 : _GEN_8219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8221 = 8'h11 == _match_key_qbytes_4_T_2 ? phv_data_17 : _GEN_8220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8222 = 8'h12 == _match_key_qbytes_4_T_2 ? phv_data_18 : _GEN_8221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8223 = 8'h13 == _match_key_qbytes_4_T_2 ? phv_data_19 : _GEN_8222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8224 = 8'h14 == _match_key_qbytes_4_T_2 ? phv_data_20 : _GEN_8223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8225 = 8'h15 == _match_key_qbytes_4_T_2 ? phv_data_21 : _GEN_8224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8226 = 8'h16 == _match_key_qbytes_4_T_2 ? phv_data_22 : _GEN_8225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8227 = 8'h17 == _match_key_qbytes_4_T_2 ? phv_data_23 : _GEN_8226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8228 = 8'h18 == _match_key_qbytes_4_T_2 ? phv_data_24 : _GEN_8227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8229 = 8'h19 == _match_key_qbytes_4_T_2 ? phv_data_25 : _GEN_8228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8230 = 8'h1a == _match_key_qbytes_4_T_2 ? phv_data_26 : _GEN_8229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8231 = 8'h1b == _match_key_qbytes_4_T_2 ? phv_data_27 : _GEN_8230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8232 = 8'h1c == _match_key_qbytes_4_T_2 ? phv_data_28 : _GEN_8231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8233 = 8'h1d == _match_key_qbytes_4_T_2 ? phv_data_29 : _GEN_8232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8234 = 8'h1e == _match_key_qbytes_4_T_2 ? phv_data_30 : _GEN_8233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8235 = 8'h1f == _match_key_qbytes_4_T_2 ? phv_data_31 : _GEN_8234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8236 = 8'h20 == _match_key_qbytes_4_T_2 ? phv_data_32 : _GEN_8235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8237 = 8'h21 == _match_key_qbytes_4_T_2 ? phv_data_33 : _GEN_8236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8238 = 8'h22 == _match_key_qbytes_4_T_2 ? phv_data_34 : _GEN_8237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8239 = 8'h23 == _match_key_qbytes_4_T_2 ? phv_data_35 : _GEN_8238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8240 = 8'h24 == _match_key_qbytes_4_T_2 ? phv_data_36 : _GEN_8239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8241 = 8'h25 == _match_key_qbytes_4_T_2 ? phv_data_37 : _GEN_8240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8242 = 8'h26 == _match_key_qbytes_4_T_2 ? phv_data_38 : _GEN_8241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8243 = 8'h27 == _match_key_qbytes_4_T_2 ? phv_data_39 : _GEN_8242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8244 = 8'h28 == _match_key_qbytes_4_T_2 ? phv_data_40 : _GEN_8243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8245 = 8'h29 == _match_key_qbytes_4_T_2 ? phv_data_41 : _GEN_8244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8246 = 8'h2a == _match_key_qbytes_4_T_2 ? phv_data_42 : _GEN_8245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8247 = 8'h2b == _match_key_qbytes_4_T_2 ? phv_data_43 : _GEN_8246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8248 = 8'h2c == _match_key_qbytes_4_T_2 ? phv_data_44 : _GEN_8247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8249 = 8'h2d == _match_key_qbytes_4_T_2 ? phv_data_45 : _GEN_8248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8250 = 8'h2e == _match_key_qbytes_4_T_2 ? phv_data_46 : _GEN_8249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8251 = 8'h2f == _match_key_qbytes_4_T_2 ? phv_data_47 : _GEN_8250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8252 = 8'h30 == _match_key_qbytes_4_T_2 ? phv_data_48 : _GEN_8251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8253 = 8'h31 == _match_key_qbytes_4_T_2 ? phv_data_49 : _GEN_8252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8254 = 8'h32 == _match_key_qbytes_4_T_2 ? phv_data_50 : _GEN_8253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8255 = 8'h33 == _match_key_qbytes_4_T_2 ? phv_data_51 : _GEN_8254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8256 = 8'h34 == _match_key_qbytes_4_T_2 ? phv_data_52 : _GEN_8255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8257 = 8'h35 == _match_key_qbytes_4_T_2 ? phv_data_53 : _GEN_8256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8258 = 8'h36 == _match_key_qbytes_4_T_2 ? phv_data_54 : _GEN_8257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8259 = 8'h37 == _match_key_qbytes_4_T_2 ? phv_data_55 : _GEN_8258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8260 = 8'h38 == _match_key_qbytes_4_T_2 ? phv_data_56 : _GEN_8259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8261 = 8'h39 == _match_key_qbytes_4_T_2 ? phv_data_57 : _GEN_8260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8262 = 8'h3a == _match_key_qbytes_4_T_2 ? phv_data_58 : _GEN_8261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8263 = 8'h3b == _match_key_qbytes_4_T_2 ? phv_data_59 : _GEN_8262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8264 = 8'h3c == _match_key_qbytes_4_T_2 ? phv_data_60 : _GEN_8263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8265 = 8'h3d == _match_key_qbytes_4_T_2 ? phv_data_61 : _GEN_8264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8266 = 8'h3e == _match_key_qbytes_4_T_2 ? phv_data_62 : _GEN_8265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8267 = 8'h3f == _match_key_qbytes_4_T_2 ? phv_data_63 : _GEN_8266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8268 = 8'h40 == _match_key_qbytes_4_T_2 ? phv_data_64 : _GEN_8267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8269 = 8'h41 == _match_key_qbytes_4_T_2 ? phv_data_65 : _GEN_8268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8270 = 8'h42 == _match_key_qbytes_4_T_2 ? phv_data_66 : _GEN_8269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8271 = 8'h43 == _match_key_qbytes_4_T_2 ? phv_data_67 : _GEN_8270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8272 = 8'h44 == _match_key_qbytes_4_T_2 ? phv_data_68 : _GEN_8271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8273 = 8'h45 == _match_key_qbytes_4_T_2 ? phv_data_69 : _GEN_8272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8274 = 8'h46 == _match_key_qbytes_4_T_2 ? phv_data_70 : _GEN_8273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8275 = 8'h47 == _match_key_qbytes_4_T_2 ? phv_data_71 : _GEN_8274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8276 = 8'h48 == _match_key_qbytes_4_T_2 ? phv_data_72 : _GEN_8275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8277 = 8'h49 == _match_key_qbytes_4_T_2 ? phv_data_73 : _GEN_8276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8278 = 8'h4a == _match_key_qbytes_4_T_2 ? phv_data_74 : _GEN_8277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8279 = 8'h4b == _match_key_qbytes_4_T_2 ? phv_data_75 : _GEN_8278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8280 = 8'h4c == _match_key_qbytes_4_T_2 ? phv_data_76 : _GEN_8279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8281 = 8'h4d == _match_key_qbytes_4_T_2 ? phv_data_77 : _GEN_8280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8282 = 8'h4e == _match_key_qbytes_4_T_2 ? phv_data_78 : _GEN_8281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8283 = 8'h4f == _match_key_qbytes_4_T_2 ? phv_data_79 : _GEN_8282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8284 = 8'h50 == _match_key_qbytes_4_T_2 ? phv_data_80 : _GEN_8283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8285 = 8'h51 == _match_key_qbytes_4_T_2 ? phv_data_81 : _GEN_8284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8286 = 8'h52 == _match_key_qbytes_4_T_2 ? phv_data_82 : _GEN_8285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8287 = 8'h53 == _match_key_qbytes_4_T_2 ? phv_data_83 : _GEN_8286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8288 = 8'h54 == _match_key_qbytes_4_T_2 ? phv_data_84 : _GEN_8287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8289 = 8'h55 == _match_key_qbytes_4_T_2 ? phv_data_85 : _GEN_8288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8290 = 8'h56 == _match_key_qbytes_4_T_2 ? phv_data_86 : _GEN_8289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8291 = 8'h57 == _match_key_qbytes_4_T_2 ? phv_data_87 : _GEN_8290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8292 = 8'h58 == _match_key_qbytes_4_T_2 ? phv_data_88 : _GEN_8291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8293 = 8'h59 == _match_key_qbytes_4_T_2 ? phv_data_89 : _GEN_8292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8294 = 8'h5a == _match_key_qbytes_4_T_2 ? phv_data_90 : _GEN_8293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8295 = 8'h5b == _match_key_qbytes_4_T_2 ? phv_data_91 : _GEN_8294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8296 = 8'h5c == _match_key_qbytes_4_T_2 ? phv_data_92 : _GEN_8295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8297 = 8'h5d == _match_key_qbytes_4_T_2 ? phv_data_93 : _GEN_8296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8298 = 8'h5e == _match_key_qbytes_4_T_2 ? phv_data_94 : _GEN_8297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8299 = 8'h5f == _match_key_qbytes_4_T_2 ? phv_data_95 : _GEN_8298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8300 = 8'h60 == _match_key_qbytes_4_T_2 ? phv_data_96 : _GEN_8299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8301 = 8'h61 == _match_key_qbytes_4_T_2 ? phv_data_97 : _GEN_8300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8302 = 8'h62 == _match_key_qbytes_4_T_2 ? phv_data_98 : _GEN_8301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8303 = 8'h63 == _match_key_qbytes_4_T_2 ? phv_data_99 : _GEN_8302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8304 = 8'h64 == _match_key_qbytes_4_T_2 ? phv_data_100 : _GEN_8303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8305 = 8'h65 == _match_key_qbytes_4_T_2 ? phv_data_101 : _GEN_8304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8306 = 8'h66 == _match_key_qbytes_4_T_2 ? phv_data_102 : _GEN_8305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8307 = 8'h67 == _match_key_qbytes_4_T_2 ? phv_data_103 : _GEN_8306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8308 = 8'h68 == _match_key_qbytes_4_T_2 ? phv_data_104 : _GEN_8307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8309 = 8'h69 == _match_key_qbytes_4_T_2 ? phv_data_105 : _GEN_8308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8310 = 8'h6a == _match_key_qbytes_4_T_2 ? phv_data_106 : _GEN_8309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8311 = 8'h6b == _match_key_qbytes_4_T_2 ? phv_data_107 : _GEN_8310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8312 = 8'h6c == _match_key_qbytes_4_T_2 ? phv_data_108 : _GEN_8311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8313 = 8'h6d == _match_key_qbytes_4_T_2 ? phv_data_109 : _GEN_8312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8314 = 8'h6e == _match_key_qbytes_4_T_2 ? phv_data_110 : _GEN_8313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8315 = 8'h6f == _match_key_qbytes_4_T_2 ? phv_data_111 : _GEN_8314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8316 = 8'h70 == _match_key_qbytes_4_T_2 ? phv_data_112 : _GEN_8315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8317 = 8'h71 == _match_key_qbytes_4_T_2 ? phv_data_113 : _GEN_8316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8318 = 8'h72 == _match_key_qbytes_4_T_2 ? phv_data_114 : _GEN_8317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8319 = 8'h73 == _match_key_qbytes_4_T_2 ? phv_data_115 : _GEN_8318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8320 = 8'h74 == _match_key_qbytes_4_T_2 ? phv_data_116 : _GEN_8319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8321 = 8'h75 == _match_key_qbytes_4_T_2 ? phv_data_117 : _GEN_8320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8322 = 8'h76 == _match_key_qbytes_4_T_2 ? phv_data_118 : _GEN_8321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8323 = 8'h77 == _match_key_qbytes_4_T_2 ? phv_data_119 : _GEN_8322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8324 = 8'h78 == _match_key_qbytes_4_T_2 ? phv_data_120 : _GEN_8323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8325 = 8'h79 == _match_key_qbytes_4_T_2 ? phv_data_121 : _GEN_8324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8326 = 8'h7a == _match_key_qbytes_4_T_2 ? phv_data_122 : _GEN_8325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8327 = 8'h7b == _match_key_qbytes_4_T_2 ? phv_data_123 : _GEN_8326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8328 = 8'h7c == _match_key_qbytes_4_T_2 ? phv_data_124 : _GEN_8327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8329 = 8'h7d == _match_key_qbytes_4_T_2 ? phv_data_125 : _GEN_8328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8330 = 8'h7e == _match_key_qbytes_4_T_2 ? phv_data_126 : _GEN_8329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8331 = 8'h7f == _match_key_qbytes_4_T_2 ? phv_data_127 : _GEN_8330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8332 = 8'h80 == _match_key_qbytes_4_T_2 ? phv_data_128 : _GEN_8331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8333 = 8'h81 == _match_key_qbytes_4_T_2 ? phv_data_129 : _GEN_8332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8334 = 8'h82 == _match_key_qbytes_4_T_2 ? phv_data_130 : _GEN_8333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8335 = 8'h83 == _match_key_qbytes_4_T_2 ? phv_data_131 : _GEN_8334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8336 = 8'h84 == _match_key_qbytes_4_T_2 ? phv_data_132 : _GEN_8335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8337 = 8'h85 == _match_key_qbytes_4_T_2 ? phv_data_133 : _GEN_8336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8338 = 8'h86 == _match_key_qbytes_4_T_2 ? phv_data_134 : _GEN_8337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8339 = 8'h87 == _match_key_qbytes_4_T_2 ? phv_data_135 : _GEN_8338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8340 = 8'h88 == _match_key_qbytes_4_T_2 ? phv_data_136 : _GEN_8339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8341 = 8'h89 == _match_key_qbytes_4_T_2 ? phv_data_137 : _GEN_8340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8342 = 8'h8a == _match_key_qbytes_4_T_2 ? phv_data_138 : _GEN_8341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8343 = 8'h8b == _match_key_qbytes_4_T_2 ? phv_data_139 : _GEN_8342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8344 = 8'h8c == _match_key_qbytes_4_T_2 ? phv_data_140 : _GEN_8343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8345 = 8'h8d == _match_key_qbytes_4_T_2 ? phv_data_141 : _GEN_8344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8346 = 8'h8e == _match_key_qbytes_4_T_2 ? phv_data_142 : _GEN_8345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8347 = 8'h8f == _match_key_qbytes_4_T_2 ? phv_data_143 : _GEN_8346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8348 = 8'h90 == _match_key_qbytes_4_T_2 ? phv_data_144 : _GEN_8347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8349 = 8'h91 == _match_key_qbytes_4_T_2 ? phv_data_145 : _GEN_8348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8350 = 8'h92 == _match_key_qbytes_4_T_2 ? phv_data_146 : _GEN_8349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8351 = 8'h93 == _match_key_qbytes_4_T_2 ? phv_data_147 : _GEN_8350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8352 = 8'h94 == _match_key_qbytes_4_T_2 ? phv_data_148 : _GEN_8351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8353 = 8'h95 == _match_key_qbytes_4_T_2 ? phv_data_149 : _GEN_8352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8354 = 8'h96 == _match_key_qbytes_4_T_2 ? phv_data_150 : _GEN_8353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8355 = 8'h97 == _match_key_qbytes_4_T_2 ? phv_data_151 : _GEN_8354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8356 = 8'h98 == _match_key_qbytes_4_T_2 ? phv_data_152 : _GEN_8355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8357 = 8'h99 == _match_key_qbytes_4_T_2 ? phv_data_153 : _GEN_8356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8358 = 8'h9a == _match_key_qbytes_4_T_2 ? phv_data_154 : _GEN_8357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8359 = 8'h9b == _match_key_qbytes_4_T_2 ? phv_data_155 : _GEN_8358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8360 = 8'h9c == _match_key_qbytes_4_T_2 ? phv_data_156 : _GEN_8359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8361 = 8'h9d == _match_key_qbytes_4_T_2 ? phv_data_157 : _GEN_8360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8362 = 8'h9e == _match_key_qbytes_4_T_2 ? phv_data_158 : _GEN_8361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8363 = 8'h9f == _match_key_qbytes_4_T_2 ? phv_data_159 : _GEN_8362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8364 = 8'ha0 == _match_key_qbytes_4_T_2 ? phv_data_160 : _GEN_8363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8365 = 8'ha1 == _match_key_qbytes_4_T_2 ? phv_data_161 : _GEN_8364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8366 = 8'ha2 == _match_key_qbytes_4_T_2 ? phv_data_162 : _GEN_8365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8367 = 8'ha3 == _match_key_qbytes_4_T_2 ? phv_data_163 : _GEN_8366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8368 = 8'ha4 == _match_key_qbytes_4_T_2 ? phv_data_164 : _GEN_8367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8369 = 8'ha5 == _match_key_qbytes_4_T_2 ? phv_data_165 : _GEN_8368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8370 = 8'ha6 == _match_key_qbytes_4_T_2 ? phv_data_166 : _GEN_8369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8371 = 8'ha7 == _match_key_qbytes_4_T_2 ? phv_data_167 : _GEN_8370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8372 = 8'ha8 == _match_key_qbytes_4_T_2 ? phv_data_168 : _GEN_8371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8373 = 8'ha9 == _match_key_qbytes_4_T_2 ? phv_data_169 : _GEN_8372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8374 = 8'haa == _match_key_qbytes_4_T_2 ? phv_data_170 : _GEN_8373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8375 = 8'hab == _match_key_qbytes_4_T_2 ? phv_data_171 : _GEN_8374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8376 = 8'hac == _match_key_qbytes_4_T_2 ? phv_data_172 : _GEN_8375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8377 = 8'had == _match_key_qbytes_4_T_2 ? phv_data_173 : _GEN_8376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8378 = 8'hae == _match_key_qbytes_4_T_2 ? phv_data_174 : _GEN_8377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8379 = 8'haf == _match_key_qbytes_4_T_2 ? phv_data_175 : _GEN_8378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8380 = 8'hb0 == _match_key_qbytes_4_T_2 ? phv_data_176 : _GEN_8379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8381 = 8'hb1 == _match_key_qbytes_4_T_2 ? phv_data_177 : _GEN_8380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8382 = 8'hb2 == _match_key_qbytes_4_T_2 ? phv_data_178 : _GEN_8381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8383 = 8'hb3 == _match_key_qbytes_4_T_2 ? phv_data_179 : _GEN_8382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8384 = 8'hb4 == _match_key_qbytes_4_T_2 ? phv_data_180 : _GEN_8383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8385 = 8'hb5 == _match_key_qbytes_4_T_2 ? phv_data_181 : _GEN_8384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8386 = 8'hb6 == _match_key_qbytes_4_T_2 ? phv_data_182 : _GEN_8385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8387 = 8'hb7 == _match_key_qbytes_4_T_2 ? phv_data_183 : _GEN_8386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8388 = 8'hb8 == _match_key_qbytes_4_T_2 ? phv_data_184 : _GEN_8387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8389 = 8'hb9 == _match_key_qbytes_4_T_2 ? phv_data_185 : _GEN_8388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8390 = 8'hba == _match_key_qbytes_4_T_2 ? phv_data_186 : _GEN_8389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8391 = 8'hbb == _match_key_qbytes_4_T_2 ? phv_data_187 : _GEN_8390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8392 = 8'hbc == _match_key_qbytes_4_T_2 ? phv_data_188 : _GEN_8391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8393 = 8'hbd == _match_key_qbytes_4_T_2 ? phv_data_189 : _GEN_8392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8394 = 8'hbe == _match_key_qbytes_4_T_2 ? phv_data_190 : _GEN_8393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8395 = 8'hbf == _match_key_qbytes_4_T_2 ? phv_data_191 : _GEN_8394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8396 = 8'hc0 == _match_key_qbytes_4_T_2 ? phv_data_192 : _GEN_8395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8397 = 8'hc1 == _match_key_qbytes_4_T_2 ? phv_data_193 : _GEN_8396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8398 = 8'hc2 == _match_key_qbytes_4_T_2 ? phv_data_194 : _GEN_8397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8399 = 8'hc3 == _match_key_qbytes_4_T_2 ? phv_data_195 : _GEN_8398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8400 = 8'hc4 == _match_key_qbytes_4_T_2 ? phv_data_196 : _GEN_8399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8401 = 8'hc5 == _match_key_qbytes_4_T_2 ? phv_data_197 : _GEN_8400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8402 = 8'hc6 == _match_key_qbytes_4_T_2 ? phv_data_198 : _GEN_8401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8403 = 8'hc7 == _match_key_qbytes_4_T_2 ? phv_data_199 : _GEN_8402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8404 = 8'hc8 == _match_key_qbytes_4_T_2 ? phv_data_200 : _GEN_8403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8405 = 8'hc9 == _match_key_qbytes_4_T_2 ? phv_data_201 : _GEN_8404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8406 = 8'hca == _match_key_qbytes_4_T_2 ? phv_data_202 : _GEN_8405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8407 = 8'hcb == _match_key_qbytes_4_T_2 ? phv_data_203 : _GEN_8406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8408 = 8'hcc == _match_key_qbytes_4_T_2 ? phv_data_204 : _GEN_8407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8409 = 8'hcd == _match_key_qbytes_4_T_2 ? phv_data_205 : _GEN_8408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8410 = 8'hce == _match_key_qbytes_4_T_2 ? phv_data_206 : _GEN_8409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8411 = 8'hcf == _match_key_qbytes_4_T_2 ? phv_data_207 : _GEN_8410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8412 = 8'hd0 == _match_key_qbytes_4_T_2 ? phv_data_208 : _GEN_8411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8413 = 8'hd1 == _match_key_qbytes_4_T_2 ? phv_data_209 : _GEN_8412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8414 = 8'hd2 == _match_key_qbytes_4_T_2 ? phv_data_210 : _GEN_8413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8415 = 8'hd3 == _match_key_qbytes_4_T_2 ? phv_data_211 : _GEN_8414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8416 = 8'hd4 == _match_key_qbytes_4_T_2 ? phv_data_212 : _GEN_8415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8417 = 8'hd5 == _match_key_qbytes_4_T_2 ? phv_data_213 : _GEN_8416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8418 = 8'hd6 == _match_key_qbytes_4_T_2 ? phv_data_214 : _GEN_8417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8419 = 8'hd7 == _match_key_qbytes_4_T_2 ? phv_data_215 : _GEN_8418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8420 = 8'hd8 == _match_key_qbytes_4_T_2 ? phv_data_216 : _GEN_8419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8421 = 8'hd9 == _match_key_qbytes_4_T_2 ? phv_data_217 : _GEN_8420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8422 = 8'hda == _match_key_qbytes_4_T_2 ? phv_data_218 : _GEN_8421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8423 = 8'hdb == _match_key_qbytes_4_T_2 ? phv_data_219 : _GEN_8422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8424 = 8'hdc == _match_key_qbytes_4_T_2 ? phv_data_220 : _GEN_8423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8425 = 8'hdd == _match_key_qbytes_4_T_2 ? phv_data_221 : _GEN_8424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8426 = 8'hde == _match_key_qbytes_4_T_2 ? phv_data_222 : _GEN_8425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8427 = 8'hdf == _match_key_qbytes_4_T_2 ? phv_data_223 : _GEN_8426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8428 = 8'he0 == _match_key_qbytes_4_T_2 ? phv_data_224 : _GEN_8427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8429 = 8'he1 == _match_key_qbytes_4_T_2 ? phv_data_225 : _GEN_8428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8430 = 8'he2 == _match_key_qbytes_4_T_2 ? phv_data_226 : _GEN_8429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8431 = 8'he3 == _match_key_qbytes_4_T_2 ? phv_data_227 : _GEN_8430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8432 = 8'he4 == _match_key_qbytes_4_T_2 ? phv_data_228 : _GEN_8431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8433 = 8'he5 == _match_key_qbytes_4_T_2 ? phv_data_229 : _GEN_8432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8434 = 8'he6 == _match_key_qbytes_4_T_2 ? phv_data_230 : _GEN_8433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8435 = 8'he7 == _match_key_qbytes_4_T_2 ? phv_data_231 : _GEN_8434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8436 = 8'he8 == _match_key_qbytes_4_T_2 ? phv_data_232 : _GEN_8435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8437 = 8'he9 == _match_key_qbytes_4_T_2 ? phv_data_233 : _GEN_8436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8438 = 8'hea == _match_key_qbytes_4_T_2 ? phv_data_234 : _GEN_8437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8439 = 8'heb == _match_key_qbytes_4_T_2 ? phv_data_235 : _GEN_8438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8440 = 8'hec == _match_key_qbytes_4_T_2 ? phv_data_236 : _GEN_8439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8441 = 8'hed == _match_key_qbytes_4_T_2 ? phv_data_237 : _GEN_8440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8442 = 8'hee == _match_key_qbytes_4_T_2 ? phv_data_238 : _GEN_8441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8443 = 8'hef == _match_key_qbytes_4_T_2 ? phv_data_239 : _GEN_8442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8444 = 8'hf0 == _match_key_qbytes_4_T_2 ? phv_data_240 : _GEN_8443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8445 = 8'hf1 == _match_key_qbytes_4_T_2 ? phv_data_241 : _GEN_8444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8446 = 8'hf2 == _match_key_qbytes_4_T_2 ? phv_data_242 : _GEN_8445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8447 = 8'hf3 == _match_key_qbytes_4_T_2 ? phv_data_243 : _GEN_8446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8448 = 8'hf4 == _match_key_qbytes_4_T_2 ? phv_data_244 : _GEN_8447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8449 = 8'hf5 == _match_key_qbytes_4_T_2 ? phv_data_245 : _GEN_8448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8450 = 8'hf6 == _match_key_qbytes_4_T_2 ? phv_data_246 : _GEN_8449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8451 = 8'hf7 == _match_key_qbytes_4_T_2 ? phv_data_247 : _GEN_8450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8452 = 8'hf8 == _match_key_qbytes_4_T_2 ? phv_data_248 : _GEN_8451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8453 = 8'hf9 == _match_key_qbytes_4_T_2 ? phv_data_249 : _GEN_8452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8454 = 8'hfa == _match_key_qbytes_4_T_2 ? phv_data_250 : _GEN_8453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8455 = 8'hfb == _match_key_qbytes_4_T_2 ? phv_data_251 : _GEN_8454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8456 = 8'hfc == _match_key_qbytes_4_T_2 ? phv_data_252 : _GEN_8455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8457 = 8'hfd == _match_key_qbytes_4_T_2 ? phv_data_253 : _GEN_8456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8458 = 8'hfe == _match_key_qbytes_4_T_2 ? phv_data_254 : _GEN_8457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8459 = 8'hff == _match_key_qbytes_4_T_2 ? phv_data_255 : _GEN_8458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_16422 = {{1'd0}, _match_key_qbytes_4_T_2}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8460 = 9'h100 == _GEN_16422 ? phv_data_256 : _GEN_8459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8461 = 9'h101 == _GEN_16422 ? phv_data_257 : _GEN_8460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8462 = 9'h102 == _GEN_16422 ? phv_data_258 : _GEN_8461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8463 = 9'h103 == _GEN_16422 ? phv_data_259 : _GEN_8462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8464 = 9'h104 == _GEN_16422 ? phv_data_260 : _GEN_8463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8465 = 9'h105 == _GEN_16422 ? phv_data_261 : _GEN_8464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8466 = 9'h106 == _GEN_16422 ? phv_data_262 : _GEN_8465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8467 = 9'h107 == _GEN_16422 ? phv_data_263 : _GEN_8466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8468 = 9'h108 == _GEN_16422 ? phv_data_264 : _GEN_8467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8469 = 9'h109 == _GEN_16422 ? phv_data_265 : _GEN_8468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8470 = 9'h10a == _GEN_16422 ? phv_data_266 : _GEN_8469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8471 = 9'h10b == _GEN_16422 ? phv_data_267 : _GEN_8470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8472 = 9'h10c == _GEN_16422 ? phv_data_268 : _GEN_8471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8473 = 9'h10d == _GEN_16422 ? phv_data_269 : _GEN_8472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8474 = 9'h10e == _GEN_16422 ? phv_data_270 : _GEN_8473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8475 = 9'h10f == _GEN_16422 ? phv_data_271 : _GEN_8474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8476 = 9'h110 == _GEN_16422 ? phv_data_272 : _GEN_8475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8477 = 9'h111 == _GEN_16422 ? phv_data_273 : _GEN_8476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8478 = 9'h112 == _GEN_16422 ? phv_data_274 : _GEN_8477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8479 = 9'h113 == _GEN_16422 ? phv_data_275 : _GEN_8478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8480 = 9'h114 == _GEN_16422 ? phv_data_276 : _GEN_8479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8481 = 9'h115 == _GEN_16422 ? phv_data_277 : _GEN_8480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8482 = 9'h116 == _GEN_16422 ? phv_data_278 : _GEN_8481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8483 = 9'h117 == _GEN_16422 ? phv_data_279 : _GEN_8482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8484 = 9'h118 == _GEN_16422 ? phv_data_280 : _GEN_8483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8485 = 9'h119 == _GEN_16422 ? phv_data_281 : _GEN_8484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8486 = 9'h11a == _GEN_16422 ? phv_data_282 : _GEN_8485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8487 = 9'h11b == _GEN_16422 ? phv_data_283 : _GEN_8486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8488 = 9'h11c == _GEN_16422 ? phv_data_284 : _GEN_8487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8489 = 9'h11d == _GEN_16422 ? phv_data_285 : _GEN_8488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8490 = 9'h11e == _GEN_16422 ? phv_data_286 : _GEN_8489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8491 = 9'h11f == _GEN_16422 ? phv_data_287 : _GEN_8490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8492 = 9'h120 == _GEN_16422 ? phv_data_288 : _GEN_8491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8493 = 9'h121 == _GEN_16422 ? phv_data_289 : _GEN_8492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8494 = 9'h122 == _GEN_16422 ? phv_data_290 : _GEN_8493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8495 = 9'h123 == _GEN_16422 ? phv_data_291 : _GEN_8494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8496 = 9'h124 == _GEN_16422 ? phv_data_292 : _GEN_8495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8497 = 9'h125 == _GEN_16422 ? phv_data_293 : _GEN_8496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8498 = 9'h126 == _GEN_16422 ? phv_data_294 : _GEN_8497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8499 = 9'h127 == _GEN_16422 ? phv_data_295 : _GEN_8498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8500 = 9'h128 == _GEN_16422 ? phv_data_296 : _GEN_8499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8501 = 9'h129 == _GEN_16422 ? phv_data_297 : _GEN_8500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8502 = 9'h12a == _GEN_16422 ? phv_data_298 : _GEN_8501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8503 = 9'h12b == _GEN_16422 ? phv_data_299 : _GEN_8502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8504 = 9'h12c == _GEN_16422 ? phv_data_300 : _GEN_8503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8505 = 9'h12d == _GEN_16422 ? phv_data_301 : _GEN_8504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8506 = 9'h12e == _GEN_16422 ? phv_data_302 : _GEN_8505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8507 = 9'h12f == _GEN_16422 ? phv_data_303 : _GEN_8506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8508 = 9'h130 == _GEN_16422 ? phv_data_304 : _GEN_8507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8509 = 9'h131 == _GEN_16422 ? phv_data_305 : _GEN_8508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8510 = 9'h132 == _GEN_16422 ? phv_data_306 : _GEN_8509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8511 = 9'h133 == _GEN_16422 ? phv_data_307 : _GEN_8510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8512 = 9'h134 == _GEN_16422 ? phv_data_308 : _GEN_8511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8513 = 9'h135 == _GEN_16422 ? phv_data_309 : _GEN_8512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8514 = 9'h136 == _GEN_16422 ? phv_data_310 : _GEN_8513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8515 = 9'h137 == _GEN_16422 ? phv_data_311 : _GEN_8514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8516 = 9'h138 == _GEN_16422 ? phv_data_312 : _GEN_8515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8517 = 9'h139 == _GEN_16422 ? phv_data_313 : _GEN_8516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8518 = 9'h13a == _GEN_16422 ? phv_data_314 : _GEN_8517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8519 = 9'h13b == _GEN_16422 ? phv_data_315 : _GEN_8518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8520 = 9'h13c == _GEN_16422 ? phv_data_316 : _GEN_8519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8521 = 9'h13d == _GEN_16422 ? phv_data_317 : _GEN_8520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8522 = 9'h13e == _GEN_16422 ? phv_data_318 : _GEN_8521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8523 = 9'h13f == _GEN_16422 ? phv_data_319 : _GEN_8522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8524 = 9'h140 == _GEN_16422 ? phv_data_320 : _GEN_8523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8525 = 9'h141 == _GEN_16422 ? phv_data_321 : _GEN_8524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8526 = 9'h142 == _GEN_16422 ? phv_data_322 : _GEN_8525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8527 = 9'h143 == _GEN_16422 ? phv_data_323 : _GEN_8526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8528 = 9'h144 == _GEN_16422 ? phv_data_324 : _GEN_8527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8529 = 9'h145 == _GEN_16422 ? phv_data_325 : _GEN_8528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8530 = 9'h146 == _GEN_16422 ? phv_data_326 : _GEN_8529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8531 = 9'h147 == _GEN_16422 ? phv_data_327 : _GEN_8530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8532 = 9'h148 == _GEN_16422 ? phv_data_328 : _GEN_8531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8533 = 9'h149 == _GEN_16422 ? phv_data_329 : _GEN_8532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8534 = 9'h14a == _GEN_16422 ? phv_data_330 : _GEN_8533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8535 = 9'h14b == _GEN_16422 ? phv_data_331 : _GEN_8534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8536 = 9'h14c == _GEN_16422 ? phv_data_332 : _GEN_8535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8537 = 9'h14d == _GEN_16422 ? phv_data_333 : _GEN_8536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8538 = 9'h14e == _GEN_16422 ? phv_data_334 : _GEN_8537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8539 = 9'h14f == _GEN_16422 ? phv_data_335 : _GEN_8538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8540 = 9'h150 == _GEN_16422 ? phv_data_336 : _GEN_8539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8541 = 9'h151 == _GEN_16422 ? phv_data_337 : _GEN_8540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8542 = 9'h152 == _GEN_16422 ? phv_data_338 : _GEN_8541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8543 = 9'h153 == _GEN_16422 ? phv_data_339 : _GEN_8542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8544 = 9'h154 == _GEN_16422 ? phv_data_340 : _GEN_8543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8545 = 9'h155 == _GEN_16422 ? phv_data_341 : _GEN_8544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8546 = 9'h156 == _GEN_16422 ? phv_data_342 : _GEN_8545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8547 = 9'h157 == _GEN_16422 ? phv_data_343 : _GEN_8546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8548 = 9'h158 == _GEN_16422 ? phv_data_344 : _GEN_8547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8549 = 9'h159 == _GEN_16422 ? phv_data_345 : _GEN_8548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8550 = 9'h15a == _GEN_16422 ? phv_data_346 : _GEN_8549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8551 = 9'h15b == _GEN_16422 ? phv_data_347 : _GEN_8550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8552 = 9'h15c == _GEN_16422 ? phv_data_348 : _GEN_8551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8553 = 9'h15d == _GEN_16422 ? phv_data_349 : _GEN_8552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8554 = 9'h15e == _GEN_16422 ? phv_data_350 : _GEN_8553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8555 = 9'h15f == _GEN_16422 ? phv_data_351 : _GEN_8554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8556 = 9'h160 == _GEN_16422 ? phv_data_352 : _GEN_8555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8557 = 9'h161 == _GEN_16422 ? phv_data_353 : _GEN_8556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8558 = 9'h162 == _GEN_16422 ? phv_data_354 : _GEN_8557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8559 = 9'h163 == _GEN_16422 ? phv_data_355 : _GEN_8558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8560 = 9'h164 == _GEN_16422 ? phv_data_356 : _GEN_8559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8561 = 9'h165 == _GEN_16422 ? phv_data_357 : _GEN_8560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8562 = 9'h166 == _GEN_16422 ? phv_data_358 : _GEN_8561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8563 = 9'h167 == _GEN_16422 ? phv_data_359 : _GEN_8562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8564 = 9'h168 == _GEN_16422 ? phv_data_360 : _GEN_8563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8565 = 9'h169 == _GEN_16422 ? phv_data_361 : _GEN_8564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8566 = 9'h16a == _GEN_16422 ? phv_data_362 : _GEN_8565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8567 = 9'h16b == _GEN_16422 ? phv_data_363 : _GEN_8566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8568 = 9'h16c == _GEN_16422 ? phv_data_364 : _GEN_8567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8569 = 9'h16d == _GEN_16422 ? phv_data_365 : _GEN_8568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8570 = 9'h16e == _GEN_16422 ? phv_data_366 : _GEN_8569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8571 = 9'h16f == _GEN_16422 ? phv_data_367 : _GEN_8570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8572 = 9'h170 == _GEN_16422 ? phv_data_368 : _GEN_8571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8573 = 9'h171 == _GEN_16422 ? phv_data_369 : _GEN_8572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8574 = 9'h172 == _GEN_16422 ? phv_data_370 : _GEN_8573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8575 = 9'h173 == _GEN_16422 ? phv_data_371 : _GEN_8574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8576 = 9'h174 == _GEN_16422 ? phv_data_372 : _GEN_8575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8577 = 9'h175 == _GEN_16422 ? phv_data_373 : _GEN_8576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8578 = 9'h176 == _GEN_16422 ? phv_data_374 : _GEN_8577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8579 = 9'h177 == _GEN_16422 ? phv_data_375 : _GEN_8578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8580 = 9'h178 == _GEN_16422 ? phv_data_376 : _GEN_8579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8581 = 9'h179 == _GEN_16422 ? phv_data_377 : _GEN_8580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8582 = 9'h17a == _GEN_16422 ? phv_data_378 : _GEN_8581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8583 = 9'h17b == _GEN_16422 ? phv_data_379 : _GEN_8582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8584 = 9'h17c == _GEN_16422 ? phv_data_380 : _GEN_8583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8585 = 9'h17d == _GEN_16422 ? phv_data_381 : _GEN_8584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8586 = 9'h17e == _GEN_16422 ? phv_data_382 : _GEN_8585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8587 = 9'h17f == _GEN_16422 ? phv_data_383 : _GEN_8586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8588 = 9'h180 == _GEN_16422 ? phv_data_384 : _GEN_8587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8589 = 9'h181 == _GEN_16422 ? phv_data_385 : _GEN_8588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8590 = 9'h182 == _GEN_16422 ? phv_data_386 : _GEN_8589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8591 = 9'h183 == _GEN_16422 ? phv_data_387 : _GEN_8590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8592 = 9'h184 == _GEN_16422 ? phv_data_388 : _GEN_8591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8593 = 9'h185 == _GEN_16422 ? phv_data_389 : _GEN_8592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8594 = 9'h186 == _GEN_16422 ? phv_data_390 : _GEN_8593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8595 = 9'h187 == _GEN_16422 ? phv_data_391 : _GEN_8594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8596 = 9'h188 == _GEN_16422 ? phv_data_392 : _GEN_8595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8597 = 9'h189 == _GEN_16422 ? phv_data_393 : _GEN_8596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8598 = 9'h18a == _GEN_16422 ? phv_data_394 : _GEN_8597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8599 = 9'h18b == _GEN_16422 ? phv_data_395 : _GEN_8598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8600 = 9'h18c == _GEN_16422 ? phv_data_396 : _GEN_8599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8601 = 9'h18d == _GEN_16422 ? phv_data_397 : _GEN_8600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8602 = 9'h18e == _GEN_16422 ? phv_data_398 : _GEN_8601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8603 = 9'h18f == _GEN_16422 ? phv_data_399 : _GEN_8602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8604 = 9'h190 == _GEN_16422 ? phv_data_400 : _GEN_8603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8605 = 9'h191 == _GEN_16422 ? phv_data_401 : _GEN_8604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8606 = 9'h192 == _GEN_16422 ? phv_data_402 : _GEN_8605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8607 = 9'h193 == _GEN_16422 ? phv_data_403 : _GEN_8606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8608 = 9'h194 == _GEN_16422 ? phv_data_404 : _GEN_8607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8609 = 9'h195 == _GEN_16422 ? phv_data_405 : _GEN_8608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8610 = 9'h196 == _GEN_16422 ? phv_data_406 : _GEN_8609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8611 = 9'h197 == _GEN_16422 ? phv_data_407 : _GEN_8610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8612 = 9'h198 == _GEN_16422 ? phv_data_408 : _GEN_8611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8613 = 9'h199 == _GEN_16422 ? phv_data_409 : _GEN_8612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8614 = 9'h19a == _GEN_16422 ? phv_data_410 : _GEN_8613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8615 = 9'h19b == _GEN_16422 ? phv_data_411 : _GEN_8614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8616 = 9'h19c == _GEN_16422 ? phv_data_412 : _GEN_8615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8617 = 9'h19d == _GEN_16422 ? phv_data_413 : _GEN_8616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8618 = 9'h19e == _GEN_16422 ? phv_data_414 : _GEN_8617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8619 = 9'h19f == _GEN_16422 ? phv_data_415 : _GEN_8618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8620 = 9'h1a0 == _GEN_16422 ? phv_data_416 : _GEN_8619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8621 = 9'h1a1 == _GEN_16422 ? phv_data_417 : _GEN_8620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8622 = 9'h1a2 == _GEN_16422 ? phv_data_418 : _GEN_8621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8623 = 9'h1a3 == _GEN_16422 ? phv_data_419 : _GEN_8622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8624 = 9'h1a4 == _GEN_16422 ? phv_data_420 : _GEN_8623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8625 = 9'h1a5 == _GEN_16422 ? phv_data_421 : _GEN_8624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8626 = 9'h1a6 == _GEN_16422 ? phv_data_422 : _GEN_8625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8627 = 9'h1a7 == _GEN_16422 ? phv_data_423 : _GEN_8626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8628 = 9'h1a8 == _GEN_16422 ? phv_data_424 : _GEN_8627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8629 = 9'h1a9 == _GEN_16422 ? phv_data_425 : _GEN_8628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8630 = 9'h1aa == _GEN_16422 ? phv_data_426 : _GEN_8629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8631 = 9'h1ab == _GEN_16422 ? phv_data_427 : _GEN_8630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8632 = 9'h1ac == _GEN_16422 ? phv_data_428 : _GEN_8631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8633 = 9'h1ad == _GEN_16422 ? phv_data_429 : _GEN_8632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8634 = 9'h1ae == _GEN_16422 ? phv_data_430 : _GEN_8633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8635 = 9'h1af == _GEN_16422 ? phv_data_431 : _GEN_8634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8636 = 9'h1b0 == _GEN_16422 ? phv_data_432 : _GEN_8635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8637 = 9'h1b1 == _GEN_16422 ? phv_data_433 : _GEN_8636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8638 = 9'h1b2 == _GEN_16422 ? phv_data_434 : _GEN_8637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8639 = 9'h1b3 == _GEN_16422 ? phv_data_435 : _GEN_8638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8640 = 9'h1b4 == _GEN_16422 ? phv_data_436 : _GEN_8639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8641 = 9'h1b5 == _GEN_16422 ? phv_data_437 : _GEN_8640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8642 = 9'h1b6 == _GEN_16422 ? phv_data_438 : _GEN_8641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8643 = 9'h1b7 == _GEN_16422 ? phv_data_439 : _GEN_8642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8644 = 9'h1b8 == _GEN_16422 ? phv_data_440 : _GEN_8643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8645 = 9'h1b9 == _GEN_16422 ? phv_data_441 : _GEN_8644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8646 = 9'h1ba == _GEN_16422 ? phv_data_442 : _GEN_8645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8647 = 9'h1bb == _GEN_16422 ? phv_data_443 : _GEN_8646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8648 = 9'h1bc == _GEN_16422 ? phv_data_444 : _GEN_8647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8649 = 9'h1bd == _GEN_16422 ? phv_data_445 : _GEN_8648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8650 = 9'h1be == _GEN_16422 ? phv_data_446 : _GEN_8649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8651 = 9'h1bf == _GEN_16422 ? phv_data_447 : _GEN_8650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8652 = 9'h1c0 == _GEN_16422 ? phv_data_448 : _GEN_8651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8653 = 9'h1c1 == _GEN_16422 ? phv_data_449 : _GEN_8652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8654 = 9'h1c2 == _GEN_16422 ? phv_data_450 : _GEN_8653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8655 = 9'h1c3 == _GEN_16422 ? phv_data_451 : _GEN_8654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8656 = 9'h1c4 == _GEN_16422 ? phv_data_452 : _GEN_8655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8657 = 9'h1c5 == _GEN_16422 ? phv_data_453 : _GEN_8656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8658 = 9'h1c6 == _GEN_16422 ? phv_data_454 : _GEN_8657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8659 = 9'h1c7 == _GEN_16422 ? phv_data_455 : _GEN_8658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8660 = 9'h1c8 == _GEN_16422 ? phv_data_456 : _GEN_8659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8661 = 9'h1c9 == _GEN_16422 ? phv_data_457 : _GEN_8660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8662 = 9'h1ca == _GEN_16422 ? phv_data_458 : _GEN_8661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8663 = 9'h1cb == _GEN_16422 ? phv_data_459 : _GEN_8662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8664 = 9'h1cc == _GEN_16422 ? phv_data_460 : _GEN_8663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8665 = 9'h1cd == _GEN_16422 ? phv_data_461 : _GEN_8664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8666 = 9'h1ce == _GEN_16422 ? phv_data_462 : _GEN_8665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8667 = 9'h1cf == _GEN_16422 ? phv_data_463 : _GEN_8666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8668 = 9'h1d0 == _GEN_16422 ? phv_data_464 : _GEN_8667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8669 = 9'h1d1 == _GEN_16422 ? phv_data_465 : _GEN_8668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8670 = 9'h1d2 == _GEN_16422 ? phv_data_466 : _GEN_8669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8671 = 9'h1d3 == _GEN_16422 ? phv_data_467 : _GEN_8670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8672 = 9'h1d4 == _GEN_16422 ? phv_data_468 : _GEN_8671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8673 = 9'h1d5 == _GEN_16422 ? phv_data_469 : _GEN_8672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8674 = 9'h1d6 == _GEN_16422 ? phv_data_470 : _GEN_8673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8675 = 9'h1d7 == _GEN_16422 ? phv_data_471 : _GEN_8674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8676 = 9'h1d8 == _GEN_16422 ? phv_data_472 : _GEN_8675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8677 = 9'h1d9 == _GEN_16422 ? phv_data_473 : _GEN_8676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8678 = 9'h1da == _GEN_16422 ? phv_data_474 : _GEN_8677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8679 = 9'h1db == _GEN_16422 ? phv_data_475 : _GEN_8678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8680 = 9'h1dc == _GEN_16422 ? phv_data_476 : _GEN_8679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8681 = 9'h1dd == _GEN_16422 ? phv_data_477 : _GEN_8680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8682 = 9'h1de == _GEN_16422 ? phv_data_478 : _GEN_8681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8683 = 9'h1df == _GEN_16422 ? phv_data_479 : _GEN_8682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8684 = 9'h1e0 == _GEN_16422 ? phv_data_480 : _GEN_8683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8685 = 9'h1e1 == _GEN_16422 ? phv_data_481 : _GEN_8684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8686 = 9'h1e2 == _GEN_16422 ? phv_data_482 : _GEN_8685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8687 = 9'h1e3 == _GEN_16422 ? phv_data_483 : _GEN_8686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8688 = 9'h1e4 == _GEN_16422 ? phv_data_484 : _GEN_8687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8689 = 9'h1e5 == _GEN_16422 ? phv_data_485 : _GEN_8688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8690 = 9'h1e6 == _GEN_16422 ? phv_data_486 : _GEN_8689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8691 = 9'h1e7 == _GEN_16422 ? phv_data_487 : _GEN_8690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8692 = 9'h1e8 == _GEN_16422 ? phv_data_488 : _GEN_8691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8693 = 9'h1e9 == _GEN_16422 ? phv_data_489 : _GEN_8692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8694 = 9'h1ea == _GEN_16422 ? phv_data_490 : _GEN_8693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8695 = 9'h1eb == _GEN_16422 ? phv_data_491 : _GEN_8694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8696 = 9'h1ec == _GEN_16422 ? phv_data_492 : _GEN_8695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8697 = 9'h1ed == _GEN_16422 ? phv_data_493 : _GEN_8696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8698 = 9'h1ee == _GEN_16422 ? phv_data_494 : _GEN_8697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8699 = 9'h1ef == _GEN_16422 ? phv_data_495 : _GEN_8698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8700 = 9'h1f0 == _GEN_16422 ? phv_data_496 : _GEN_8699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8701 = 9'h1f1 == _GEN_16422 ? phv_data_497 : _GEN_8700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8702 = 9'h1f2 == _GEN_16422 ? phv_data_498 : _GEN_8701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8703 = 9'h1f3 == _GEN_16422 ? phv_data_499 : _GEN_8702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8704 = 9'h1f4 == _GEN_16422 ? phv_data_500 : _GEN_8703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8705 = 9'h1f5 == _GEN_16422 ? phv_data_501 : _GEN_8704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8706 = 9'h1f6 == _GEN_16422 ? phv_data_502 : _GEN_8705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8707 = 9'h1f7 == _GEN_16422 ? phv_data_503 : _GEN_8706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8708 = 9'h1f8 == _GEN_16422 ? phv_data_504 : _GEN_8707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8709 = 9'h1f9 == _GEN_16422 ? phv_data_505 : _GEN_8708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8710 = 9'h1fa == _GEN_16422 ? phv_data_506 : _GEN_8709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8711 = 9'h1fb == _GEN_16422 ? phv_data_507 : _GEN_8710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8712 = 9'h1fc == _GEN_16422 ? phv_data_508 : _GEN_8711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8713 = 9'h1fd == _GEN_16422 ? phv_data_509 : _GEN_8712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8714 = 9'h1fe == _GEN_16422 ? phv_data_510 : _GEN_8713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8715 = 9'h1ff == _GEN_16422 ? phv_data_511 : _GEN_8714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8717 = 8'h1 == local_offset_4 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8718 = 8'h2 == local_offset_4 ? phv_data_2 : _GEN_8717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8719 = 8'h3 == local_offset_4 ? phv_data_3 : _GEN_8718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8720 = 8'h4 == local_offset_4 ? phv_data_4 : _GEN_8719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8721 = 8'h5 == local_offset_4 ? phv_data_5 : _GEN_8720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8722 = 8'h6 == local_offset_4 ? phv_data_6 : _GEN_8721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8723 = 8'h7 == local_offset_4 ? phv_data_7 : _GEN_8722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8724 = 8'h8 == local_offset_4 ? phv_data_8 : _GEN_8723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8725 = 8'h9 == local_offset_4 ? phv_data_9 : _GEN_8724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8726 = 8'ha == local_offset_4 ? phv_data_10 : _GEN_8725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8727 = 8'hb == local_offset_4 ? phv_data_11 : _GEN_8726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8728 = 8'hc == local_offset_4 ? phv_data_12 : _GEN_8727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8729 = 8'hd == local_offset_4 ? phv_data_13 : _GEN_8728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8730 = 8'he == local_offset_4 ? phv_data_14 : _GEN_8729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8731 = 8'hf == local_offset_4 ? phv_data_15 : _GEN_8730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8732 = 8'h10 == local_offset_4 ? phv_data_16 : _GEN_8731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8733 = 8'h11 == local_offset_4 ? phv_data_17 : _GEN_8732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8734 = 8'h12 == local_offset_4 ? phv_data_18 : _GEN_8733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8735 = 8'h13 == local_offset_4 ? phv_data_19 : _GEN_8734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8736 = 8'h14 == local_offset_4 ? phv_data_20 : _GEN_8735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8737 = 8'h15 == local_offset_4 ? phv_data_21 : _GEN_8736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8738 = 8'h16 == local_offset_4 ? phv_data_22 : _GEN_8737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8739 = 8'h17 == local_offset_4 ? phv_data_23 : _GEN_8738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8740 = 8'h18 == local_offset_4 ? phv_data_24 : _GEN_8739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8741 = 8'h19 == local_offset_4 ? phv_data_25 : _GEN_8740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8742 = 8'h1a == local_offset_4 ? phv_data_26 : _GEN_8741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8743 = 8'h1b == local_offset_4 ? phv_data_27 : _GEN_8742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8744 = 8'h1c == local_offset_4 ? phv_data_28 : _GEN_8743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8745 = 8'h1d == local_offset_4 ? phv_data_29 : _GEN_8744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8746 = 8'h1e == local_offset_4 ? phv_data_30 : _GEN_8745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8747 = 8'h1f == local_offset_4 ? phv_data_31 : _GEN_8746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8748 = 8'h20 == local_offset_4 ? phv_data_32 : _GEN_8747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8749 = 8'h21 == local_offset_4 ? phv_data_33 : _GEN_8748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8750 = 8'h22 == local_offset_4 ? phv_data_34 : _GEN_8749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8751 = 8'h23 == local_offset_4 ? phv_data_35 : _GEN_8750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8752 = 8'h24 == local_offset_4 ? phv_data_36 : _GEN_8751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8753 = 8'h25 == local_offset_4 ? phv_data_37 : _GEN_8752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8754 = 8'h26 == local_offset_4 ? phv_data_38 : _GEN_8753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8755 = 8'h27 == local_offset_4 ? phv_data_39 : _GEN_8754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8756 = 8'h28 == local_offset_4 ? phv_data_40 : _GEN_8755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8757 = 8'h29 == local_offset_4 ? phv_data_41 : _GEN_8756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8758 = 8'h2a == local_offset_4 ? phv_data_42 : _GEN_8757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8759 = 8'h2b == local_offset_4 ? phv_data_43 : _GEN_8758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8760 = 8'h2c == local_offset_4 ? phv_data_44 : _GEN_8759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8761 = 8'h2d == local_offset_4 ? phv_data_45 : _GEN_8760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8762 = 8'h2e == local_offset_4 ? phv_data_46 : _GEN_8761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8763 = 8'h2f == local_offset_4 ? phv_data_47 : _GEN_8762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8764 = 8'h30 == local_offset_4 ? phv_data_48 : _GEN_8763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8765 = 8'h31 == local_offset_4 ? phv_data_49 : _GEN_8764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8766 = 8'h32 == local_offset_4 ? phv_data_50 : _GEN_8765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8767 = 8'h33 == local_offset_4 ? phv_data_51 : _GEN_8766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8768 = 8'h34 == local_offset_4 ? phv_data_52 : _GEN_8767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8769 = 8'h35 == local_offset_4 ? phv_data_53 : _GEN_8768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8770 = 8'h36 == local_offset_4 ? phv_data_54 : _GEN_8769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8771 = 8'h37 == local_offset_4 ? phv_data_55 : _GEN_8770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8772 = 8'h38 == local_offset_4 ? phv_data_56 : _GEN_8771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8773 = 8'h39 == local_offset_4 ? phv_data_57 : _GEN_8772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8774 = 8'h3a == local_offset_4 ? phv_data_58 : _GEN_8773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8775 = 8'h3b == local_offset_4 ? phv_data_59 : _GEN_8774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8776 = 8'h3c == local_offset_4 ? phv_data_60 : _GEN_8775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8777 = 8'h3d == local_offset_4 ? phv_data_61 : _GEN_8776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8778 = 8'h3e == local_offset_4 ? phv_data_62 : _GEN_8777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8779 = 8'h3f == local_offset_4 ? phv_data_63 : _GEN_8778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8780 = 8'h40 == local_offset_4 ? phv_data_64 : _GEN_8779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8781 = 8'h41 == local_offset_4 ? phv_data_65 : _GEN_8780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8782 = 8'h42 == local_offset_4 ? phv_data_66 : _GEN_8781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8783 = 8'h43 == local_offset_4 ? phv_data_67 : _GEN_8782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8784 = 8'h44 == local_offset_4 ? phv_data_68 : _GEN_8783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8785 = 8'h45 == local_offset_4 ? phv_data_69 : _GEN_8784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8786 = 8'h46 == local_offset_4 ? phv_data_70 : _GEN_8785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8787 = 8'h47 == local_offset_4 ? phv_data_71 : _GEN_8786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8788 = 8'h48 == local_offset_4 ? phv_data_72 : _GEN_8787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8789 = 8'h49 == local_offset_4 ? phv_data_73 : _GEN_8788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8790 = 8'h4a == local_offset_4 ? phv_data_74 : _GEN_8789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8791 = 8'h4b == local_offset_4 ? phv_data_75 : _GEN_8790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8792 = 8'h4c == local_offset_4 ? phv_data_76 : _GEN_8791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8793 = 8'h4d == local_offset_4 ? phv_data_77 : _GEN_8792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8794 = 8'h4e == local_offset_4 ? phv_data_78 : _GEN_8793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8795 = 8'h4f == local_offset_4 ? phv_data_79 : _GEN_8794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8796 = 8'h50 == local_offset_4 ? phv_data_80 : _GEN_8795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8797 = 8'h51 == local_offset_4 ? phv_data_81 : _GEN_8796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8798 = 8'h52 == local_offset_4 ? phv_data_82 : _GEN_8797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8799 = 8'h53 == local_offset_4 ? phv_data_83 : _GEN_8798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8800 = 8'h54 == local_offset_4 ? phv_data_84 : _GEN_8799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8801 = 8'h55 == local_offset_4 ? phv_data_85 : _GEN_8800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8802 = 8'h56 == local_offset_4 ? phv_data_86 : _GEN_8801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8803 = 8'h57 == local_offset_4 ? phv_data_87 : _GEN_8802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8804 = 8'h58 == local_offset_4 ? phv_data_88 : _GEN_8803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8805 = 8'h59 == local_offset_4 ? phv_data_89 : _GEN_8804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8806 = 8'h5a == local_offset_4 ? phv_data_90 : _GEN_8805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8807 = 8'h5b == local_offset_4 ? phv_data_91 : _GEN_8806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8808 = 8'h5c == local_offset_4 ? phv_data_92 : _GEN_8807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8809 = 8'h5d == local_offset_4 ? phv_data_93 : _GEN_8808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8810 = 8'h5e == local_offset_4 ? phv_data_94 : _GEN_8809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8811 = 8'h5f == local_offset_4 ? phv_data_95 : _GEN_8810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8812 = 8'h60 == local_offset_4 ? phv_data_96 : _GEN_8811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8813 = 8'h61 == local_offset_4 ? phv_data_97 : _GEN_8812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8814 = 8'h62 == local_offset_4 ? phv_data_98 : _GEN_8813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8815 = 8'h63 == local_offset_4 ? phv_data_99 : _GEN_8814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8816 = 8'h64 == local_offset_4 ? phv_data_100 : _GEN_8815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8817 = 8'h65 == local_offset_4 ? phv_data_101 : _GEN_8816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8818 = 8'h66 == local_offset_4 ? phv_data_102 : _GEN_8817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8819 = 8'h67 == local_offset_4 ? phv_data_103 : _GEN_8818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8820 = 8'h68 == local_offset_4 ? phv_data_104 : _GEN_8819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8821 = 8'h69 == local_offset_4 ? phv_data_105 : _GEN_8820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8822 = 8'h6a == local_offset_4 ? phv_data_106 : _GEN_8821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8823 = 8'h6b == local_offset_4 ? phv_data_107 : _GEN_8822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8824 = 8'h6c == local_offset_4 ? phv_data_108 : _GEN_8823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8825 = 8'h6d == local_offset_4 ? phv_data_109 : _GEN_8824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8826 = 8'h6e == local_offset_4 ? phv_data_110 : _GEN_8825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8827 = 8'h6f == local_offset_4 ? phv_data_111 : _GEN_8826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8828 = 8'h70 == local_offset_4 ? phv_data_112 : _GEN_8827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8829 = 8'h71 == local_offset_4 ? phv_data_113 : _GEN_8828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8830 = 8'h72 == local_offset_4 ? phv_data_114 : _GEN_8829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8831 = 8'h73 == local_offset_4 ? phv_data_115 : _GEN_8830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8832 = 8'h74 == local_offset_4 ? phv_data_116 : _GEN_8831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8833 = 8'h75 == local_offset_4 ? phv_data_117 : _GEN_8832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8834 = 8'h76 == local_offset_4 ? phv_data_118 : _GEN_8833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8835 = 8'h77 == local_offset_4 ? phv_data_119 : _GEN_8834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8836 = 8'h78 == local_offset_4 ? phv_data_120 : _GEN_8835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8837 = 8'h79 == local_offset_4 ? phv_data_121 : _GEN_8836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8838 = 8'h7a == local_offset_4 ? phv_data_122 : _GEN_8837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8839 = 8'h7b == local_offset_4 ? phv_data_123 : _GEN_8838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8840 = 8'h7c == local_offset_4 ? phv_data_124 : _GEN_8839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8841 = 8'h7d == local_offset_4 ? phv_data_125 : _GEN_8840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8842 = 8'h7e == local_offset_4 ? phv_data_126 : _GEN_8841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8843 = 8'h7f == local_offset_4 ? phv_data_127 : _GEN_8842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8844 = 8'h80 == local_offset_4 ? phv_data_128 : _GEN_8843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8845 = 8'h81 == local_offset_4 ? phv_data_129 : _GEN_8844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8846 = 8'h82 == local_offset_4 ? phv_data_130 : _GEN_8845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8847 = 8'h83 == local_offset_4 ? phv_data_131 : _GEN_8846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8848 = 8'h84 == local_offset_4 ? phv_data_132 : _GEN_8847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8849 = 8'h85 == local_offset_4 ? phv_data_133 : _GEN_8848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8850 = 8'h86 == local_offset_4 ? phv_data_134 : _GEN_8849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8851 = 8'h87 == local_offset_4 ? phv_data_135 : _GEN_8850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8852 = 8'h88 == local_offset_4 ? phv_data_136 : _GEN_8851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8853 = 8'h89 == local_offset_4 ? phv_data_137 : _GEN_8852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8854 = 8'h8a == local_offset_4 ? phv_data_138 : _GEN_8853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8855 = 8'h8b == local_offset_4 ? phv_data_139 : _GEN_8854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8856 = 8'h8c == local_offset_4 ? phv_data_140 : _GEN_8855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8857 = 8'h8d == local_offset_4 ? phv_data_141 : _GEN_8856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8858 = 8'h8e == local_offset_4 ? phv_data_142 : _GEN_8857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8859 = 8'h8f == local_offset_4 ? phv_data_143 : _GEN_8858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8860 = 8'h90 == local_offset_4 ? phv_data_144 : _GEN_8859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8861 = 8'h91 == local_offset_4 ? phv_data_145 : _GEN_8860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8862 = 8'h92 == local_offset_4 ? phv_data_146 : _GEN_8861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8863 = 8'h93 == local_offset_4 ? phv_data_147 : _GEN_8862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8864 = 8'h94 == local_offset_4 ? phv_data_148 : _GEN_8863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8865 = 8'h95 == local_offset_4 ? phv_data_149 : _GEN_8864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8866 = 8'h96 == local_offset_4 ? phv_data_150 : _GEN_8865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8867 = 8'h97 == local_offset_4 ? phv_data_151 : _GEN_8866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8868 = 8'h98 == local_offset_4 ? phv_data_152 : _GEN_8867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8869 = 8'h99 == local_offset_4 ? phv_data_153 : _GEN_8868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8870 = 8'h9a == local_offset_4 ? phv_data_154 : _GEN_8869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8871 = 8'h9b == local_offset_4 ? phv_data_155 : _GEN_8870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8872 = 8'h9c == local_offset_4 ? phv_data_156 : _GEN_8871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8873 = 8'h9d == local_offset_4 ? phv_data_157 : _GEN_8872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8874 = 8'h9e == local_offset_4 ? phv_data_158 : _GEN_8873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8875 = 8'h9f == local_offset_4 ? phv_data_159 : _GEN_8874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8876 = 8'ha0 == local_offset_4 ? phv_data_160 : _GEN_8875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8877 = 8'ha1 == local_offset_4 ? phv_data_161 : _GEN_8876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8878 = 8'ha2 == local_offset_4 ? phv_data_162 : _GEN_8877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8879 = 8'ha3 == local_offset_4 ? phv_data_163 : _GEN_8878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8880 = 8'ha4 == local_offset_4 ? phv_data_164 : _GEN_8879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8881 = 8'ha5 == local_offset_4 ? phv_data_165 : _GEN_8880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8882 = 8'ha6 == local_offset_4 ? phv_data_166 : _GEN_8881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8883 = 8'ha7 == local_offset_4 ? phv_data_167 : _GEN_8882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8884 = 8'ha8 == local_offset_4 ? phv_data_168 : _GEN_8883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8885 = 8'ha9 == local_offset_4 ? phv_data_169 : _GEN_8884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8886 = 8'haa == local_offset_4 ? phv_data_170 : _GEN_8885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8887 = 8'hab == local_offset_4 ? phv_data_171 : _GEN_8886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8888 = 8'hac == local_offset_4 ? phv_data_172 : _GEN_8887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8889 = 8'had == local_offset_4 ? phv_data_173 : _GEN_8888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8890 = 8'hae == local_offset_4 ? phv_data_174 : _GEN_8889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8891 = 8'haf == local_offset_4 ? phv_data_175 : _GEN_8890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8892 = 8'hb0 == local_offset_4 ? phv_data_176 : _GEN_8891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8893 = 8'hb1 == local_offset_4 ? phv_data_177 : _GEN_8892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8894 = 8'hb2 == local_offset_4 ? phv_data_178 : _GEN_8893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8895 = 8'hb3 == local_offset_4 ? phv_data_179 : _GEN_8894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8896 = 8'hb4 == local_offset_4 ? phv_data_180 : _GEN_8895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8897 = 8'hb5 == local_offset_4 ? phv_data_181 : _GEN_8896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8898 = 8'hb6 == local_offset_4 ? phv_data_182 : _GEN_8897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8899 = 8'hb7 == local_offset_4 ? phv_data_183 : _GEN_8898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8900 = 8'hb8 == local_offset_4 ? phv_data_184 : _GEN_8899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8901 = 8'hb9 == local_offset_4 ? phv_data_185 : _GEN_8900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8902 = 8'hba == local_offset_4 ? phv_data_186 : _GEN_8901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8903 = 8'hbb == local_offset_4 ? phv_data_187 : _GEN_8902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8904 = 8'hbc == local_offset_4 ? phv_data_188 : _GEN_8903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8905 = 8'hbd == local_offset_4 ? phv_data_189 : _GEN_8904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8906 = 8'hbe == local_offset_4 ? phv_data_190 : _GEN_8905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8907 = 8'hbf == local_offset_4 ? phv_data_191 : _GEN_8906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8908 = 8'hc0 == local_offset_4 ? phv_data_192 : _GEN_8907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8909 = 8'hc1 == local_offset_4 ? phv_data_193 : _GEN_8908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8910 = 8'hc2 == local_offset_4 ? phv_data_194 : _GEN_8909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8911 = 8'hc3 == local_offset_4 ? phv_data_195 : _GEN_8910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8912 = 8'hc4 == local_offset_4 ? phv_data_196 : _GEN_8911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8913 = 8'hc5 == local_offset_4 ? phv_data_197 : _GEN_8912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8914 = 8'hc6 == local_offset_4 ? phv_data_198 : _GEN_8913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8915 = 8'hc7 == local_offset_4 ? phv_data_199 : _GEN_8914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8916 = 8'hc8 == local_offset_4 ? phv_data_200 : _GEN_8915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8917 = 8'hc9 == local_offset_4 ? phv_data_201 : _GEN_8916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8918 = 8'hca == local_offset_4 ? phv_data_202 : _GEN_8917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8919 = 8'hcb == local_offset_4 ? phv_data_203 : _GEN_8918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8920 = 8'hcc == local_offset_4 ? phv_data_204 : _GEN_8919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8921 = 8'hcd == local_offset_4 ? phv_data_205 : _GEN_8920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8922 = 8'hce == local_offset_4 ? phv_data_206 : _GEN_8921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8923 = 8'hcf == local_offset_4 ? phv_data_207 : _GEN_8922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8924 = 8'hd0 == local_offset_4 ? phv_data_208 : _GEN_8923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8925 = 8'hd1 == local_offset_4 ? phv_data_209 : _GEN_8924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8926 = 8'hd2 == local_offset_4 ? phv_data_210 : _GEN_8925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8927 = 8'hd3 == local_offset_4 ? phv_data_211 : _GEN_8926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8928 = 8'hd4 == local_offset_4 ? phv_data_212 : _GEN_8927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8929 = 8'hd5 == local_offset_4 ? phv_data_213 : _GEN_8928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8930 = 8'hd6 == local_offset_4 ? phv_data_214 : _GEN_8929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8931 = 8'hd7 == local_offset_4 ? phv_data_215 : _GEN_8930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8932 = 8'hd8 == local_offset_4 ? phv_data_216 : _GEN_8931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8933 = 8'hd9 == local_offset_4 ? phv_data_217 : _GEN_8932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8934 = 8'hda == local_offset_4 ? phv_data_218 : _GEN_8933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8935 = 8'hdb == local_offset_4 ? phv_data_219 : _GEN_8934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8936 = 8'hdc == local_offset_4 ? phv_data_220 : _GEN_8935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8937 = 8'hdd == local_offset_4 ? phv_data_221 : _GEN_8936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8938 = 8'hde == local_offset_4 ? phv_data_222 : _GEN_8937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8939 = 8'hdf == local_offset_4 ? phv_data_223 : _GEN_8938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8940 = 8'he0 == local_offset_4 ? phv_data_224 : _GEN_8939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8941 = 8'he1 == local_offset_4 ? phv_data_225 : _GEN_8940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8942 = 8'he2 == local_offset_4 ? phv_data_226 : _GEN_8941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8943 = 8'he3 == local_offset_4 ? phv_data_227 : _GEN_8942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8944 = 8'he4 == local_offset_4 ? phv_data_228 : _GEN_8943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8945 = 8'he5 == local_offset_4 ? phv_data_229 : _GEN_8944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8946 = 8'he6 == local_offset_4 ? phv_data_230 : _GEN_8945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8947 = 8'he7 == local_offset_4 ? phv_data_231 : _GEN_8946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8948 = 8'he8 == local_offset_4 ? phv_data_232 : _GEN_8947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8949 = 8'he9 == local_offset_4 ? phv_data_233 : _GEN_8948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8950 = 8'hea == local_offset_4 ? phv_data_234 : _GEN_8949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8951 = 8'heb == local_offset_4 ? phv_data_235 : _GEN_8950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8952 = 8'hec == local_offset_4 ? phv_data_236 : _GEN_8951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8953 = 8'hed == local_offset_4 ? phv_data_237 : _GEN_8952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8954 = 8'hee == local_offset_4 ? phv_data_238 : _GEN_8953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8955 = 8'hef == local_offset_4 ? phv_data_239 : _GEN_8954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8956 = 8'hf0 == local_offset_4 ? phv_data_240 : _GEN_8955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8957 = 8'hf1 == local_offset_4 ? phv_data_241 : _GEN_8956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8958 = 8'hf2 == local_offset_4 ? phv_data_242 : _GEN_8957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8959 = 8'hf3 == local_offset_4 ? phv_data_243 : _GEN_8958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8960 = 8'hf4 == local_offset_4 ? phv_data_244 : _GEN_8959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8961 = 8'hf5 == local_offset_4 ? phv_data_245 : _GEN_8960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8962 = 8'hf6 == local_offset_4 ? phv_data_246 : _GEN_8961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8963 = 8'hf7 == local_offset_4 ? phv_data_247 : _GEN_8962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8964 = 8'hf8 == local_offset_4 ? phv_data_248 : _GEN_8963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8965 = 8'hf9 == local_offset_4 ? phv_data_249 : _GEN_8964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8966 = 8'hfa == local_offset_4 ? phv_data_250 : _GEN_8965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8967 = 8'hfb == local_offset_4 ? phv_data_251 : _GEN_8966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8968 = 8'hfc == local_offset_4 ? phv_data_252 : _GEN_8967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8969 = 8'hfd == local_offset_4 ? phv_data_253 : _GEN_8968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8970 = 8'hfe == local_offset_4 ? phv_data_254 : _GEN_8969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8971 = 8'hff == local_offset_4 ? phv_data_255 : _GEN_8970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_16678 = {{1'd0}, local_offset_4}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8972 = 9'h100 == _GEN_16678 ? phv_data_256 : _GEN_8971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8973 = 9'h101 == _GEN_16678 ? phv_data_257 : _GEN_8972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8974 = 9'h102 == _GEN_16678 ? phv_data_258 : _GEN_8973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8975 = 9'h103 == _GEN_16678 ? phv_data_259 : _GEN_8974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8976 = 9'h104 == _GEN_16678 ? phv_data_260 : _GEN_8975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8977 = 9'h105 == _GEN_16678 ? phv_data_261 : _GEN_8976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8978 = 9'h106 == _GEN_16678 ? phv_data_262 : _GEN_8977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8979 = 9'h107 == _GEN_16678 ? phv_data_263 : _GEN_8978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8980 = 9'h108 == _GEN_16678 ? phv_data_264 : _GEN_8979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8981 = 9'h109 == _GEN_16678 ? phv_data_265 : _GEN_8980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8982 = 9'h10a == _GEN_16678 ? phv_data_266 : _GEN_8981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8983 = 9'h10b == _GEN_16678 ? phv_data_267 : _GEN_8982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8984 = 9'h10c == _GEN_16678 ? phv_data_268 : _GEN_8983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8985 = 9'h10d == _GEN_16678 ? phv_data_269 : _GEN_8984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8986 = 9'h10e == _GEN_16678 ? phv_data_270 : _GEN_8985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8987 = 9'h10f == _GEN_16678 ? phv_data_271 : _GEN_8986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8988 = 9'h110 == _GEN_16678 ? phv_data_272 : _GEN_8987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8989 = 9'h111 == _GEN_16678 ? phv_data_273 : _GEN_8988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8990 = 9'h112 == _GEN_16678 ? phv_data_274 : _GEN_8989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8991 = 9'h113 == _GEN_16678 ? phv_data_275 : _GEN_8990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8992 = 9'h114 == _GEN_16678 ? phv_data_276 : _GEN_8991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8993 = 9'h115 == _GEN_16678 ? phv_data_277 : _GEN_8992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8994 = 9'h116 == _GEN_16678 ? phv_data_278 : _GEN_8993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8995 = 9'h117 == _GEN_16678 ? phv_data_279 : _GEN_8994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8996 = 9'h118 == _GEN_16678 ? phv_data_280 : _GEN_8995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8997 = 9'h119 == _GEN_16678 ? phv_data_281 : _GEN_8996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8998 = 9'h11a == _GEN_16678 ? phv_data_282 : _GEN_8997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8999 = 9'h11b == _GEN_16678 ? phv_data_283 : _GEN_8998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9000 = 9'h11c == _GEN_16678 ? phv_data_284 : _GEN_8999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9001 = 9'h11d == _GEN_16678 ? phv_data_285 : _GEN_9000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9002 = 9'h11e == _GEN_16678 ? phv_data_286 : _GEN_9001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9003 = 9'h11f == _GEN_16678 ? phv_data_287 : _GEN_9002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9004 = 9'h120 == _GEN_16678 ? phv_data_288 : _GEN_9003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9005 = 9'h121 == _GEN_16678 ? phv_data_289 : _GEN_9004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9006 = 9'h122 == _GEN_16678 ? phv_data_290 : _GEN_9005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9007 = 9'h123 == _GEN_16678 ? phv_data_291 : _GEN_9006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9008 = 9'h124 == _GEN_16678 ? phv_data_292 : _GEN_9007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9009 = 9'h125 == _GEN_16678 ? phv_data_293 : _GEN_9008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9010 = 9'h126 == _GEN_16678 ? phv_data_294 : _GEN_9009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9011 = 9'h127 == _GEN_16678 ? phv_data_295 : _GEN_9010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9012 = 9'h128 == _GEN_16678 ? phv_data_296 : _GEN_9011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9013 = 9'h129 == _GEN_16678 ? phv_data_297 : _GEN_9012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9014 = 9'h12a == _GEN_16678 ? phv_data_298 : _GEN_9013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9015 = 9'h12b == _GEN_16678 ? phv_data_299 : _GEN_9014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9016 = 9'h12c == _GEN_16678 ? phv_data_300 : _GEN_9015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9017 = 9'h12d == _GEN_16678 ? phv_data_301 : _GEN_9016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9018 = 9'h12e == _GEN_16678 ? phv_data_302 : _GEN_9017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9019 = 9'h12f == _GEN_16678 ? phv_data_303 : _GEN_9018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9020 = 9'h130 == _GEN_16678 ? phv_data_304 : _GEN_9019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9021 = 9'h131 == _GEN_16678 ? phv_data_305 : _GEN_9020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9022 = 9'h132 == _GEN_16678 ? phv_data_306 : _GEN_9021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9023 = 9'h133 == _GEN_16678 ? phv_data_307 : _GEN_9022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9024 = 9'h134 == _GEN_16678 ? phv_data_308 : _GEN_9023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9025 = 9'h135 == _GEN_16678 ? phv_data_309 : _GEN_9024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9026 = 9'h136 == _GEN_16678 ? phv_data_310 : _GEN_9025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9027 = 9'h137 == _GEN_16678 ? phv_data_311 : _GEN_9026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9028 = 9'h138 == _GEN_16678 ? phv_data_312 : _GEN_9027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9029 = 9'h139 == _GEN_16678 ? phv_data_313 : _GEN_9028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9030 = 9'h13a == _GEN_16678 ? phv_data_314 : _GEN_9029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9031 = 9'h13b == _GEN_16678 ? phv_data_315 : _GEN_9030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9032 = 9'h13c == _GEN_16678 ? phv_data_316 : _GEN_9031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9033 = 9'h13d == _GEN_16678 ? phv_data_317 : _GEN_9032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9034 = 9'h13e == _GEN_16678 ? phv_data_318 : _GEN_9033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9035 = 9'h13f == _GEN_16678 ? phv_data_319 : _GEN_9034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9036 = 9'h140 == _GEN_16678 ? phv_data_320 : _GEN_9035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9037 = 9'h141 == _GEN_16678 ? phv_data_321 : _GEN_9036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9038 = 9'h142 == _GEN_16678 ? phv_data_322 : _GEN_9037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9039 = 9'h143 == _GEN_16678 ? phv_data_323 : _GEN_9038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9040 = 9'h144 == _GEN_16678 ? phv_data_324 : _GEN_9039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9041 = 9'h145 == _GEN_16678 ? phv_data_325 : _GEN_9040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9042 = 9'h146 == _GEN_16678 ? phv_data_326 : _GEN_9041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9043 = 9'h147 == _GEN_16678 ? phv_data_327 : _GEN_9042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9044 = 9'h148 == _GEN_16678 ? phv_data_328 : _GEN_9043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9045 = 9'h149 == _GEN_16678 ? phv_data_329 : _GEN_9044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9046 = 9'h14a == _GEN_16678 ? phv_data_330 : _GEN_9045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9047 = 9'h14b == _GEN_16678 ? phv_data_331 : _GEN_9046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9048 = 9'h14c == _GEN_16678 ? phv_data_332 : _GEN_9047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9049 = 9'h14d == _GEN_16678 ? phv_data_333 : _GEN_9048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9050 = 9'h14e == _GEN_16678 ? phv_data_334 : _GEN_9049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9051 = 9'h14f == _GEN_16678 ? phv_data_335 : _GEN_9050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9052 = 9'h150 == _GEN_16678 ? phv_data_336 : _GEN_9051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9053 = 9'h151 == _GEN_16678 ? phv_data_337 : _GEN_9052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9054 = 9'h152 == _GEN_16678 ? phv_data_338 : _GEN_9053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9055 = 9'h153 == _GEN_16678 ? phv_data_339 : _GEN_9054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9056 = 9'h154 == _GEN_16678 ? phv_data_340 : _GEN_9055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9057 = 9'h155 == _GEN_16678 ? phv_data_341 : _GEN_9056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9058 = 9'h156 == _GEN_16678 ? phv_data_342 : _GEN_9057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9059 = 9'h157 == _GEN_16678 ? phv_data_343 : _GEN_9058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9060 = 9'h158 == _GEN_16678 ? phv_data_344 : _GEN_9059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9061 = 9'h159 == _GEN_16678 ? phv_data_345 : _GEN_9060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9062 = 9'h15a == _GEN_16678 ? phv_data_346 : _GEN_9061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9063 = 9'h15b == _GEN_16678 ? phv_data_347 : _GEN_9062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9064 = 9'h15c == _GEN_16678 ? phv_data_348 : _GEN_9063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9065 = 9'h15d == _GEN_16678 ? phv_data_349 : _GEN_9064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9066 = 9'h15e == _GEN_16678 ? phv_data_350 : _GEN_9065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9067 = 9'h15f == _GEN_16678 ? phv_data_351 : _GEN_9066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9068 = 9'h160 == _GEN_16678 ? phv_data_352 : _GEN_9067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9069 = 9'h161 == _GEN_16678 ? phv_data_353 : _GEN_9068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9070 = 9'h162 == _GEN_16678 ? phv_data_354 : _GEN_9069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9071 = 9'h163 == _GEN_16678 ? phv_data_355 : _GEN_9070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9072 = 9'h164 == _GEN_16678 ? phv_data_356 : _GEN_9071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9073 = 9'h165 == _GEN_16678 ? phv_data_357 : _GEN_9072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9074 = 9'h166 == _GEN_16678 ? phv_data_358 : _GEN_9073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9075 = 9'h167 == _GEN_16678 ? phv_data_359 : _GEN_9074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9076 = 9'h168 == _GEN_16678 ? phv_data_360 : _GEN_9075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9077 = 9'h169 == _GEN_16678 ? phv_data_361 : _GEN_9076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9078 = 9'h16a == _GEN_16678 ? phv_data_362 : _GEN_9077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9079 = 9'h16b == _GEN_16678 ? phv_data_363 : _GEN_9078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9080 = 9'h16c == _GEN_16678 ? phv_data_364 : _GEN_9079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9081 = 9'h16d == _GEN_16678 ? phv_data_365 : _GEN_9080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9082 = 9'h16e == _GEN_16678 ? phv_data_366 : _GEN_9081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9083 = 9'h16f == _GEN_16678 ? phv_data_367 : _GEN_9082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9084 = 9'h170 == _GEN_16678 ? phv_data_368 : _GEN_9083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9085 = 9'h171 == _GEN_16678 ? phv_data_369 : _GEN_9084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9086 = 9'h172 == _GEN_16678 ? phv_data_370 : _GEN_9085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9087 = 9'h173 == _GEN_16678 ? phv_data_371 : _GEN_9086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9088 = 9'h174 == _GEN_16678 ? phv_data_372 : _GEN_9087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9089 = 9'h175 == _GEN_16678 ? phv_data_373 : _GEN_9088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9090 = 9'h176 == _GEN_16678 ? phv_data_374 : _GEN_9089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9091 = 9'h177 == _GEN_16678 ? phv_data_375 : _GEN_9090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9092 = 9'h178 == _GEN_16678 ? phv_data_376 : _GEN_9091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9093 = 9'h179 == _GEN_16678 ? phv_data_377 : _GEN_9092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9094 = 9'h17a == _GEN_16678 ? phv_data_378 : _GEN_9093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9095 = 9'h17b == _GEN_16678 ? phv_data_379 : _GEN_9094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9096 = 9'h17c == _GEN_16678 ? phv_data_380 : _GEN_9095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9097 = 9'h17d == _GEN_16678 ? phv_data_381 : _GEN_9096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9098 = 9'h17e == _GEN_16678 ? phv_data_382 : _GEN_9097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9099 = 9'h17f == _GEN_16678 ? phv_data_383 : _GEN_9098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9100 = 9'h180 == _GEN_16678 ? phv_data_384 : _GEN_9099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9101 = 9'h181 == _GEN_16678 ? phv_data_385 : _GEN_9100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9102 = 9'h182 == _GEN_16678 ? phv_data_386 : _GEN_9101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9103 = 9'h183 == _GEN_16678 ? phv_data_387 : _GEN_9102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9104 = 9'h184 == _GEN_16678 ? phv_data_388 : _GEN_9103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9105 = 9'h185 == _GEN_16678 ? phv_data_389 : _GEN_9104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9106 = 9'h186 == _GEN_16678 ? phv_data_390 : _GEN_9105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9107 = 9'h187 == _GEN_16678 ? phv_data_391 : _GEN_9106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9108 = 9'h188 == _GEN_16678 ? phv_data_392 : _GEN_9107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9109 = 9'h189 == _GEN_16678 ? phv_data_393 : _GEN_9108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9110 = 9'h18a == _GEN_16678 ? phv_data_394 : _GEN_9109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9111 = 9'h18b == _GEN_16678 ? phv_data_395 : _GEN_9110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9112 = 9'h18c == _GEN_16678 ? phv_data_396 : _GEN_9111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9113 = 9'h18d == _GEN_16678 ? phv_data_397 : _GEN_9112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9114 = 9'h18e == _GEN_16678 ? phv_data_398 : _GEN_9113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9115 = 9'h18f == _GEN_16678 ? phv_data_399 : _GEN_9114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9116 = 9'h190 == _GEN_16678 ? phv_data_400 : _GEN_9115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9117 = 9'h191 == _GEN_16678 ? phv_data_401 : _GEN_9116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9118 = 9'h192 == _GEN_16678 ? phv_data_402 : _GEN_9117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9119 = 9'h193 == _GEN_16678 ? phv_data_403 : _GEN_9118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9120 = 9'h194 == _GEN_16678 ? phv_data_404 : _GEN_9119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9121 = 9'h195 == _GEN_16678 ? phv_data_405 : _GEN_9120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9122 = 9'h196 == _GEN_16678 ? phv_data_406 : _GEN_9121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9123 = 9'h197 == _GEN_16678 ? phv_data_407 : _GEN_9122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9124 = 9'h198 == _GEN_16678 ? phv_data_408 : _GEN_9123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9125 = 9'h199 == _GEN_16678 ? phv_data_409 : _GEN_9124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9126 = 9'h19a == _GEN_16678 ? phv_data_410 : _GEN_9125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9127 = 9'h19b == _GEN_16678 ? phv_data_411 : _GEN_9126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9128 = 9'h19c == _GEN_16678 ? phv_data_412 : _GEN_9127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9129 = 9'h19d == _GEN_16678 ? phv_data_413 : _GEN_9128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9130 = 9'h19e == _GEN_16678 ? phv_data_414 : _GEN_9129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9131 = 9'h19f == _GEN_16678 ? phv_data_415 : _GEN_9130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9132 = 9'h1a0 == _GEN_16678 ? phv_data_416 : _GEN_9131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9133 = 9'h1a1 == _GEN_16678 ? phv_data_417 : _GEN_9132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9134 = 9'h1a2 == _GEN_16678 ? phv_data_418 : _GEN_9133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9135 = 9'h1a3 == _GEN_16678 ? phv_data_419 : _GEN_9134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9136 = 9'h1a4 == _GEN_16678 ? phv_data_420 : _GEN_9135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9137 = 9'h1a5 == _GEN_16678 ? phv_data_421 : _GEN_9136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9138 = 9'h1a6 == _GEN_16678 ? phv_data_422 : _GEN_9137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9139 = 9'h1a7 == _GEN_16678 ? phv_data_423 : _GEN_9138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9140 = 9'h1a8 == _GEN_16678 ? phv_data_424 : _GEN_9139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9141 = 9'h1a9 == _GEN_16678 ? phv_data_425 : _GEN_9140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9142 = 9'h1aa == _GEN_16678 ? phv_data_426 : _GEN_9141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9143 = 9'h1ab == _GEN_16678 ? phv_data_427 : _GEN_9142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9144 = 9'h1ac == _GEN_16678 ? phv_data_428 : _GEN_9143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9145 = 9'h1ad == _GEN_16678 ? phv_data_429 : _GEN_9144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9146 = 9'h1ae == _GEN_16678 ? phv_data_430 : _GEN_9145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9147 = 9'h1af == _GEN_16678 ? phv_data_431 : _GEN_9146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9148 = 9'h1b0 == _GEN_16678 ? phv_data_432 : _GEN_9147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9149 = 9'h1b1 == _GEN_16678 ? phv_data_433 : _GEN_9148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9150 = 9'h1b2 == _GEN_16678 ? phv_data_434 : _GEN_9149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9151 = 9'h1b3 == _GEN_16678 ? phv_data_435 : _GEN_9150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9152 = 9'h1b4 == _GEN_16678 ? phv_data_436 : _GEN_9151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9153 = 9'h1b5 == _GEN_16678 ? phv_data_437 : _GEN_9152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9154 = 9'h1b6 == _GEN_16678 ? phv_data_438 : _GEN_9153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9155 = 9'h1b7 == _GEN_16678 ? phv_data_439 : _GEN_9154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9156 = 9'h1b8 == _GEN_16678 ? phv_data_440 : _GEN_9155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9157 = 9'h1b9 == _GEN_16678 ? phv_data_441 : _GEN_9156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9158 = 9'h1ba == _GEN_16678 ? phv_data_442 : _GEN_9157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9159 = 9'h1bb == _GEN_16678 ? phv_data_443 : _GEN_9158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9160 = 9'h1bc == _GEN_16678 ? phv_data_444 : _GEN_9159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9161 = 9'h1bd == _GEN_16678 ? phv_data_445 : _GEN_9160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9162 = 9'h1be == _GEN_16678 ? phv_data_446 : _GEN_9161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9163 = 9'h1bf == _GEN_16678 ? phv_data_447 : _GEN_9162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9164 = 9'h1c0 == _GEN_16678 ? phv_data_448 : _GEN_9163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9165 = 9'h1c1 == _GEN_16678 ? phv_data_449 : _GEN_9164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9166 = 9'h1c2 == _GEN_16678 ? phv_data_450 : _GEN_9165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9167 = 9'h1c3 == _GEN_16678 ? phv_data_451 : _GEN_9166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9168 = 9'h1c4 == _GEN_16678 ? phv_data_452 : _GEN_9167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9169 = 9'h1c5 == _GEN_16678 ? phv_data_453 : _GEN_9168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9170 = 9'h1c6 == _GEN_16678 ? phv_data_454 : _GEN_9169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9171 = 9'h1c7 == _GEN_16678 ? phv_data_455 : _GEN_9170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9172 = 9'h1c8 == _GEN_16678 ? phv_data_456 : _GEN_9171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9173 = 9'h1c9 == _GEN_16678 ? phv_data_457 : _GEN_9172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9174 = 9'h1ca == _GEN_16678 ? phv_data_458 : _GEN_9173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9175 = 9'h1cb == _GEN_16678 ? phv_data_459 : _GEN_9174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9176 = 9'h1cc == _GEN_16678 ? phv_data_460 : _GEN_9175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9177 = 9'h1cd == _GEN_16678 ? phv_data_461 : _GEN_9176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9178 = 9'h1ce == _GEN_16678 ? phv_data_462 : _GEN_9177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9179 = 9'h1cf == _GEN_16678 ? phv_data_463 : _GEN_9178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9180 = 9'h1d0 == _GEN_16678 ? phv_data_464 : _GEN_9179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9181 = 9'h1d1 == _GEN_16678 ? phv_data_465 : _GEN_9180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9182 = 9'h1d2 == _GEN_16678 ? phv_data_466 : _GEN_9181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9183 = 9'h1d3 == _GEN_16678 ? phv_data_467 : _GEN_9182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9184 = 9'h1d4 == _GEN_16678 ? phv_data_468 : _GEN_9183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9185 = 9'h1d5 == _GEN_16678 ? phv_data_469 : _GEN_9184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9186 = 9'h1d6 == _GEN_16678 ? phv_data_470 : _GEN_9185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9187 = 9'h1d7 == _GEN_16678 ? phv_data_471 : _GEN_9186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9188 = 9'h1d8 == _GEN_16678 ? phv_data_472 : _GEN_9187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9189 = 9'h1d9 == _GEN_16678 ? phv_data_473 : _GEN_9188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9190 = 9'h1da == _GEN_16678 ? phv_data_474 : _GEN_9189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9191 = 9'h1db == _GEN_16678 ? phv_data_475 : _GEN_9190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9192 = 9'h1dc == _GEN_16678 ? phv_data_476 : _GEN_9191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9193 = 9'h1dd == _GEN_16678 ? phv_data_477 : _GEN_9192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9194 = 9'h1de == _GEN_16678 ? phv_data_478 : _GEN_9193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9195 = 9'h1df == _GEN_16678 ? phv_data_479 : _GEN_9194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9196 = 9'h1e0 == _GEN_16678 ? phv_data_480 : _GEN_9195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9197 = 9'h1e1 == _GEN_16678 ? phv_data_481 : _GEN_9196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9198 = 9'h1e2 == _GEN_16678 ? phv_data_482 : _GEN_9197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9199 = 9'h1e3 == _GEN_16678 ? phv_data_483 : _GEN_9198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9200 = 9'h1e4 == _GEN_16678 ? phv_data_484 : _GEN_9199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9201 = 9'h1e5 == _GEN_16678 ? phv_data_485 : _GEN_9200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9202 = 9'h1e6 == _GEN_16678 ? phv_data_486 : _GEN_9201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9203 = 9'h1e7 == _GEN_16678 ? phv_data_487 : _GEN_9202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9204 = 9'h1e8 == _GEN_16678 ? phv_data_488 : _GEN_9203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9205 = 9'h1e9 == _GEN_16678 ? phv_data_489 : _GEN_9204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9206 = 9'h1ea == _GEN_16678 ? phv_data_490 : _GEN_9205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9207 = 9'h1eb == _GEN_16678 ? phv_data_491 : _GEN_9206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9208 = 9'h1ec == _GEN_16678 ? phv_data_492 : _GEN_9207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9209 = 9'h1ed == _GEN_16678 ? phv_data_493 : _GEN_9208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9210 = 9'h1ee == _GEN_16678 ? phv_data_494 : _GEN_9209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9211 = 9'h1ef == _GEN_16678 ? phv_data_495 : _GEN_9210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9212 = 9'h1f0 == _GEN_16678 ? phv_data_496 : _GEN_9211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9213 = 9'h1f1 == _GEN_16678 ? phv_data_497 : _GEN_9212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9214 = 9'h1f2 == _GEN_16678 ? phv_data_498 : _GEN_9213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9215 = 9'h1f3 == _GEN_16678 ? phv_data_499 : _GEN_9214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9216 = 9'h1f4 == _GEN_16678 ? phv_data_500 : _GEN_9215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9217 = 9'h1f5 == _GEN_16678 ? phv_data_501 : _GEN_9216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9218 = 9'h1f6 == _GEN_16678 ? phv_data_502 : _GEN_9217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9219 = 9'h1f7 == _GEN_16678 ? phv_data_503 : _GEN_9218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9220 = 9'h1f8 == _GEN_16678 ? phv_data_504 : _GEN_9219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9221 = 9'h1f9 == _GEN_16678 ? phv_data_505 : _GEN_9220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9222 = 9'h1fa == _GEN_16678 ? phv_data_506 : _GEN_9221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9223 = 9'h1fb == _GEN_16678 ? phv_data_507 : _GEN_9222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9224 = 9'h1fc == _GEN_16678 ? phv_data_508 : _GEN_9223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9225 = 9'h1fd == _GEN_16678 ? phv_data_509 : _GEN_9224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9226 = 9'h1fe == _GEN_16678 ? phv_data_510 : _GEN_9225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9227 = 9'h1ff == _GEN_16678 ? phv_data_511 : _GEN_9226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9229 = 8'h1 == _match_key_qbytes_4_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9230 = 8'h2 == _match_key_qbytes_4_T ? phv_data_2 : _GEN_9229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9231 = 8'h3 == _match_key_qbytes_4_T ? phv_data_3 : _GEN_9230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9232 = 8'h4 == _match_key_qbytes_4_T ? phv_data_4 : _GEN_9231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9233 = 8'h5 == _match_key_qbytes_4_T ? phv_data_5 : _GEN_9232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9234 = 8'h6 == _match_key_qbytes_4_T ? phv_data_6 : _GEN_9233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9235 = 8'h7 == _match_key_qbytes_4_T ? phv_data_7 : _GEN_9234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9236 = 8'h8 == _match_key_qbytes_4_T ? phv_data_8 : _GEN_9235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9237 = 8'h9 == _match_key_qbytes_4_T ? phv_data_9 : _GEN_9236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9238 = 8'ha == _match_key_qbytes_4_T ? phv_data_10 : _GEN_9237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9239 = 8'hb == _match_key_qbytes_4_T ? phv_data_11 : _GEN_9238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9240 = 8'hc == _match_key_qbytes_4_T ? phv_data_12 : _GEN_9239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9241 = 8'hd == _match_key_qbytes_4_T ? phv_data_13 : _GEN_9240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9242 = 8'he == _match_key_qbytes_4_T ? phv_data_14 : _GEN_9241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9243 = 8'hf == _match_key_qbytes_4_T ? phv_data_15 : _GEN_9242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9244 = 8'h10 == _match_key_qbytes_4_T ? phv_data_16 : _GEN_9243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9245 = 8'h11 == _match_key_qbytes_4_T ? phv_data_17 : _GEN_9244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9246 = 8'h12 == _match_key_qbytes_4_T ? phv_data_18 : _GEN_9245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9247 = 8'h13 == _match_key_qbytes_4_T ? phv_data_19 : _GEN_9246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9248 = 8'h14 == _match_key_qbytes_4_T ? phv_data_20 : _GEN_9247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9249 = 8'h15 == _match_key_qbytes_4_T ? phv_data_21 : _GEN_9248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9250 = 8'h16 == _match_key_qbytes_4_T ? phv_data_22 : _GEN_9249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9251 = 8'h17 == _match_key_qbytes_4_T ? phv_data_23 : _GEN_9250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9252 = 8'h18 == _match_key_qbytes_4_T ? phv_data_24 : _GEN_9251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9253 = 8'h19 == _match_key_qbytes_4_T ? phv_data_25 : _GEN_9252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9254 = 8'h1a == _match_key_qbytes_4_T ? phv_data_26 : _GEN_9253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9255 = 8'h1b == _match_key_qbytes_4_T ? phv_data_27 : _GEN_9254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9256 = 8'h1c == _match_key_qbytes_4_T ? phv_data_28 : _GEN_9255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9257 = 8'h1d == _match_key_qbytes_4_T ? phv_data_29 : _GEN_9256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9258 = 8'h1e == _match_key_qbytes_4_T ? phv_data_30 : _GEN_9257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9259 = 8'h1f == _match_key_qbytes_4_T ? phv_data_31 : _GEN_9258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9260 = 8'h20 == _match_key_qbytes_4_T ? phv_data_32 : _GEN_9259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9261 = 8'h21 == _match_key_qbytes_4_T ? phv_data_33 : _GEN_9260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9262 = 8'h22 == _match_key_qbytes_4_T ? phv_data_34 : _GEN_9261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9263 = 8'h23 == _match_key_qbytes_4_T ? phv_data_35 : _GEN_9262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9264 = 8'h24 == _match_key_qbytes_4_T ? phv_data_36 : _GEN_9263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9265 = 8'h25 == _match_key_qbytes_4_T ? phv_data_37 : _GEN_9264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9266 = 8'h26 == _match_key_qbytes_4_T ? phv_data_38 : _GEN_9265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9267 = 8'h27 == _match_key_qbytes_4_T ? phv_data_39 : _GEN_9266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9268 = 8'h28 == _match_key_qbytes_4_T ? phv_data_40 : _GEN_9267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9269 = 8'h29 == _match_key_qbytes_4_T ? phv_data_41 : _GEN_9268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9270 = 8'h2a == _match_key_qbytes_4_T ? phv_data_42 : _GEN_9269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9271 = 8'h2b == _match_key_qbytes_4_T ? phv_data_43 : _GEN_9270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9272 = 8'h2c == _match_key_qbytes_4_T ? phv_data_44 : _GEN_9271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9273 = 8'h2d == _match_key_qbytes_4_T ? phv_data_45 : _GEN_9272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9274 = 8'h2e == _match_key_qbytes_4_T ? phv_data_46 : _GEN_9273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9275 = 8'h2f == _match_key_qbytes_4_T ? phv_data_47 : _GEN_9274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9276 = 8'h30 == _match_key_qbytes_4_T ? phv_data_48 : _GEN_9275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9277 = 8'h31 == _match_key_qbytes_4_T ? phv_data_49 : _GEN_9276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9278 = 8'h32 == _match_key_qbytes_4_T ? phv_data_50 : _GEN_9277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9279 = 8'h33 == _match_key_qbytes_4_T ? phv_data_51 : _GEN_9278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9280 = 8'h34 == _match_key_qbytes_4_T ? phv_data_52 : _GEN_9279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9281 = 8'h35 == _match_key_qbytes_4_T ? phv_data_53 : _GEN_9280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9282 = 8'h36 == _match_key_qbytes_4_T ? phv_data_54 : _GEN_9281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9283 = 8'h37 == _match_key_qbytes_4_T ? phv_data_55 : _GEN_9282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9284 = 8'h38 == _match_key_qbytes_4_T ? phv_data_56 : _GEN_9283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9285 = 8'h39 == _match_key_qbytes_4_T ? phv_data_57 : _GEN_9284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9286 = 8'h3a == _match_key_qbytes_4_T ? phv_data_58 : _GEN_9285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9287 = 8'h3b == _match_key_qbytes_4_T ? phv_data_59 : _GEN_9286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9288 = 8'h3c == _match_key_qbytes_4_T ? phv_data_60 : _GEN_9287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9289 = 8'h3d == _match_key_qbytes_4_T ? phv_data_61 : _GEN_9288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9290 = 8'h3e == _match_key_qbytes_4_T ? phv_data_62 : _GEN_9289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9291 = 8'h3f == _match_key_qbytes_4_T ? phv_data_63 : _GEN_9290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9292 = 8'h40 == _match_key_qbytes_4_T ? phv_data_64 : _GEN_9291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9293 = 8'h41 == _match_key_qbytes_4_T ? phv_data_65 : _GEN_9292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9294 = 8'h42 == _match_key_qbytes_4_T ? phv_data_66 : _GEN_9293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9295 = 8'h43 == _match_key_qbytes_4_T ? phv_data_67 : _GEN_9294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9296 = 8'h44 == _match_key_qbytes_4_T ? phv_data_68 : _GEN_9295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9297 = 8'h45 == _match_key_qbytes_4_T ? phv_data_69 : _GEN_9296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9298 = 8'h46 == _match_key_qbytes_4_T ? phv_data_70 : _GEN_9297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9299 = 8'h47 == _match_key_qbytes_4_T ? phv_data_71 : _GEN_9298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9300 = 8'h48 == _match_key_qbytes_4_T ? phv_data_72 : _GEN_9299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9301 = 8'h49 == _match_key_qbytes_4_T ? phv_data_73 : _GEN_9300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9302 = 8'h4a == _match_key_qbytes_4_T ? phv_data_74 : _GEN_9301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9303 = 8'h4b == _match_key_qbytes_4_T ? phv_data_75 : _GEN_9302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9304 = 8'h4c == _match_key_qbytes_4_T ? phv_data_76 : _GEN_9303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9305 = 8'h4d == _match_key_qbytes_4_T ? phv_data_77 : _GEN_9304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9306 = 8'h4e == _match_key_qbytes_4_T ? phv_data_78 : _GEN_9305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9307 = 8'h4f == _match_key_qbytes_4_T ? phv_data_79 : _GEN_9306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9308 = 8'h50 == _match_key_qbytes_4_T ? phv_data_80 : _GEN_9307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9309 = 8'h51 == _match_key_qbytes_4_T ? phv_data_81 : _GEN_9308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9310 = 8'h52 == _match_key_qbytes_4_T ? phv_data_82 : _GEN_9309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9311 = 8'h53 == _match_key_qbytes_4_T ? phv_data_83 : _GEN_9310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9312 = 8'h54 == _match_key_qbytes_4_T ? phv_data_84 : _GEN_9311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9313 = 8'h55 == _match_key_qbytes_4_T ? phv_data_85 : _GEN_9312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9314 = 8'h56 == _match_key_qbytes_4_T ? phv_data_86 : _GEN_9313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9315 = 8'h57 == _match_key_qbytes_4_T ? phv_data_87 : _GEN_9314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9316 = 8'h58 == _match_key_qbytes_4_T ? phv_data_88 : _GEN_9315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9317 = 8'h59 == _match_key_qbytes_4_T ? phv_data_89 : _GEN_9316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9318 = 8'h5a == _match_key_qbytes_4_T ? phv_data_90 : _GEN_9317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9319 = 8'h5b == _match_key_qbytes_4_T ? phv_data_91 : _GEN_9318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9320 = 8'h5c == _match_key_qbytes_4_T ? phv_data_92 : _GEN_9319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9321 = 8'h5d == _match_key_qbytes_4_T ? phv_data_93 : _GEN_9320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9322 = 8'h5e == _match_key_qbytes_4_T ? phv_data_94 : _GEN_9321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9323 = 8'h5f == _match_key_qbytes_4_T ? phv_data_95 : _GEN_9322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9324 = 8'h60 == _match_key_qbytes_4_T ? phv_data_96 : _GEN_9323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9325 = 8'h61 == _match_key_qbytes_4_T ? phv_data_97 : _GEN_9324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9326 = 8'h62 == _match_key_qbytes_4_T ? phv_data_98 : _GEN_9325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9327 = 8'h63 == _match_key_qbytes_4_T ? phv_data_99 : _GEN_9326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9328 = 8'h64 == _match_key_qbytes_4_T ? phv_data_100 : _GEN_9327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9329 = 8'h65 == _match_key_qbytes_4_T ? phv_data_101 : _GEN_9328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9330 = 8'h66 == _match_key_qbytes_4_T ? phv_data_102 : _GEN_9329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9331 = 8'h67 == _match_key_qbytes_4_T ? phv_data_103 : _GEN_9330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9332 = 8'h68 == _match_key_qbytes_4_T ? phv_data_104 : _GEN_9331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9333 = 8'h69 == _match_key_qbytes_4_T ? phv_data_105 : _GEN_9332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9334 = 8'h6a == _match_key_qbytes_4_T ? phv_data_106 : _GEN_9333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9335 = 8'h6b == _match_key_qbytes_4_T ? phv_data_107 : _GEN_9334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9336 = 8'h6c == _match_key_qbytes_4_T ? phv_data_108 : _GEN_9335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9337 = 8'h6d == _match_key_qbytes_4_T ? phv_data_109 : _GEN_9336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9338 = 8'h6e == _match_key_qbytes_4_T ? phv_data_110 : _GEN_9337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9339 = 8'h6f == _match_key_qbytes_4_T ? phv_data_111 : _GEN_9338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9340 = 8'h70 == _match_key_qbytes_4_T ? phv_data_112 : _GEN_9339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9341 = 8'h71 == _match_key_qbytes_4_T ? phv_data_113 : _GEN_9340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9342 = 8'h72 == _match_key_qbytes_4_T ? phv_data_114 : _GEN_9341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9343 = 8'h73 == _match_key_qbytes_4_T ? phv_data_115 : _GEN_9342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9344 = 8'h74 == _match_key_qbytes_4_T ? phv_data_116 : _GEN_9343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9345 = 8'h75 == _match_key_qbytes_4_T ? phv_data_117 : _GEN_9344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9346 = 8'h76 == _match_key_qbytes_4_T ? phv_data_118 : _GEN_9345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9347 = 8'h77 == _match_key_qbytes_4_T ? phv_data_119 : _GEN_9346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9348 = 8'h78 == _match_key_qbytes_4_T ? phv_data_120 : _GEN_9347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9349 = 8'h79 == _match_key_qbytes_4_T ? phv_data_121 : _GEN_9348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9350 = 8'h7a == _match_key_qbytes_4_T ? phv_data_122 : _GEN_9349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9351 = 8'h7b == _match_key_qbytes_4_T ? phv_data_123 : _GEN_9350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9352 = 8'h7c == _match_key_qbytes_4_T ? phv_data_124 : _GEN_9351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9353 = 8'h7d == _match_key_qbytes_4_T ? phv_data_125 : _GEN_9352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9354 = 8'h7e == _match_key_qbytes_4_T ? phv_data_126 : _GEN_9353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9355 = 8'h7f == _match_key_qbytes_4_T ? phv_data_127 : _GEN_9354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9356 = 8'h80 == _match_key_qbytes_4_T ? phv_data_128 : _GEN_9355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9357 = 8'h81 == _match_key_qbytes_4_T ? phv_data_129 : _GEN_9356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9358 = 8'h82 == _match_key_qbytes_4_T ? phv_data_130 : _GEN_9357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9359 = 8'h83 == _match_key_qbytes_4_T ? phv_data_131 : _GEN_9358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9360 = 8'h84 == _match_key_qbytes_4_T ? phv_data_132 : _GEN_9359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9361 = 8'h85 == _match_key_qbytes_4_T ? phv_data_133 : _GEN_9360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9362 = 8'h86 == _match_key_qbytes_4_T ? phv_data_134 : _GEN_9361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9363 = 8'h87 == _match_key_qbytes_4_T ? phv_data_135 : _GEN_9362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9364 = 8'h88 == _match_key_qbytes_4_T ? phv_data_136 : _GEN_9363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9365 = 8'h89 == _match_key_qbytes_4_T ? phv_data_137 : _GEN_9364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9366 = 8'h8a == _match_key_qbytes_4_T ? phv_data_138 : _GEN_9365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9367 = 8'h8b == _match_key_qbytes_4_T ? phv_data_139 : _GEN_9366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9368 = 8'h8c == _match_key_qbytes_4_T ? phv_data_140 : _GEN_9367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9369 = 8'h8d == _match_key_qbytes_4_T ? phv_data_141 : _GEN_9368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9370 = 8'h8e == _match_key_qbytes_4_T ? phv_data_142 : _GEN_9369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9371 = 8'h8f == _match_key_qbytes_4_T ? phv_data_143 : _GEN_9370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9372 = 8'h90 == _match_key_qbytes_4_T ? phv_data_144 : _GEN_9371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9373 = 8'h91 == _match_key_qbytes_4_T ? phv_data_145 : _GEN_9372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9374 = 8'h92 == _match_key_qbytes_4_T ? phv_data_146 : _GEN_9373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9375 = 8'h93 == _match_key_qbytes_4_T ? phv_data_147 : _GEN_9374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9376 = 8'h94 == _match_key_qbytes_4_T ? phv_data_148 : _GEN_9375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9377 = 8'h95 == _match_key_qbytes_4_T ? phv_data_149 : _GEN_9376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9378 = 8'h96 == _match_key_qbytes_4_T ? phv_data_150 : _GEN_9377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9379 = 8'h97 == _match_key_qbytes_4_T ? phv_data_151 : _GEN_9378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9380 = 8'h98 == _match_key_qbytes_4_T ? phv_data_152 : _GEN_9379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9381 = 8'h99 == _match_key_qbytes_4_T ? phv_data_153 : _GEN_9380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9382 = 8'h9a == _match_key_qbytes_4_T ? phv_data_154 : _GEN_9381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9383 = 8'h9b == _match_key_qbytes_4_T ? phv_data_155 : _GEN_9382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9384 = 8'h9c == _match_key_qbytes_4_T ? phv_data_156 : _GEN_9383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9385 = 8'h9d == _match_key_qbytes_4_T ? phv_data_157 : _GEN_9384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9386 = 8'h9e == _match_key_qbytes_4_T ? phv_data_158 : _GEN_9385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9387 = 8'h9f == _match_key_qbytes_4_T ? phv_data_159 : _GEN_9386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9388 = 8'ha0 == _match_key_qbytes_4_T ? phv_data_160 : _GEN_9387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9389 = 8'ha1 == _match_key_qbytes_4_T ? phv_data_161 : _GEN_9388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9390 = 8'ha2 == _match_key_qbytes_4_T ? phv_data_162 : _GEN_9389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9391 = 8'ha3 == _match_key_qbytes_4_T ? phv_data_163 : _GEN_9390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9392 = 8'ha4 == _match_key_qbytes_4_T ? phv_data_164 : _GEN_9391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9393 = 8'ha5 == _match_key_qbytes_4_T ? phv_data_165 : _GEN_9392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9394 = 8'ha6 == _match_key_qbytes_4_T ? phv_data_166 : _GEN_9393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9395 = 8'ha7 == _match_key_qbytes_4_T ? phv_data_167 : _GEN_9394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9396 = 8'ha8 == _match_key_qbytes_4_T ? phv_data_168 : _GEN_9395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9397 = 8'ha9 == _match_key_qbytes_4_T ? phv_data_169 : _GEN_9396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9398 = 8'haa == _match_key_qbytes_4_T ? phv_data_170 : _GEN_9397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9399 = 8'hab == _match_key_qbytes_4_T ? phv_data_171 : _GEN_9398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9400 = 8'hac == _match_key_qbytes_4_T ? phv_data_172 : _GEN_9399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9401 = 8'had == _match_key_qbytes_4_T ? phv_data_173 : _GEN_9400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9402 = 8'hae == _match_key_qbytes_4_T ? phv_data_174 : _GEN_9401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9403 = 8'haf == _match_key_qbytes_4_T ? phv_data_175 : _GEN_9402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9404 = 8'hb0 == _match_key_qbytes_4_T ? phv_data_176 : _GEN_9403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9405 = 8'hb1 == _match_key_qbytes_4_T ? phv_data_177 : _GEN_9404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9406 = 8'hb2 == _match_key_qbytes_4_T ? phv_data_178 : _GEN_9405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9407 = 8'hb3 == _match_key_qbytes_4_T ? phv_data_179 : _GEN_9406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9408 = 8'hb4 == _match_key_qbytes_4_T ? phv_data_180 : _GEN_9407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9409 = 8'hb5 == _match_key_qbytes_4_T ? phv_data_181 : _GEN_9408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9410 = 8'hb6 == _match_key_qbytes_4_T ? phv_data_182 : _GEN_9409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9411 = 8'hb7 == _match_key_qbytes_4_T ? phv_data_183 : _GEN_9410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9412 = 8'hb8 == _match_key_qbytes_4_T ? phv_data_184 : _GEN_9411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9413 = 8'hb9 == _match_key_qbytes_4_T ? phv_data_185 : _GEN_9412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9414 = 8'hba == _match_key_qbytes_4_T ? phv_data_186 : _GEN_9413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9415 = 8'hbb == _match_key_qbytes_4_T ? phv_data_187 : _GEN_9414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9416 = 8'hbc == _match_key_qbytes_4_T ? phv_data_188 : _GEN_9415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9417 = 8'hbd == _match_key_qbytes_4_T ? phv_data_189 : _GEN_9416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9418 = 8'hbe == _match_key_qbytes_4_T ? phv_data_190 : _GEN_9417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9419 = 8'hbf == _match_key_qbytes_4_T ? phv_data_191 : _GEN_9418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9420 = 8'hc0 == _match_key_qbytes_4_T ? phv_data_192 : _GEN_9419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9421 = 8'hc1 == _match_key_qbytes_4_T ? phv_data_193 : _GEN_9420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9422 = 8'hc2 == _match_key_qbytes_4_T ? phv_data_194 : _GEN_9421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9423 = 8'hc3 == _match_key_qbytes_4_T ? phv_data_195 : _GEN_9422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9424 = 8'hc4 == _match_key_qbytes_4_T ? phv_data_196 : _GEN_9423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9425 = 8'hc5 == _match_key_qbytes_4_T ? phv_data_197 : _GEN_9424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9426 = 8'hc6 == _match_key_qbytes_4_T ? phv_data_198 : _GEN_9425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9427 = 8'hc7 == _match_key_qbytes_4_T ? phv_data_199 : _GEN_9426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9428 = 8'hc8 == _match_key_qbytes_4_T ? phv_data_200 : _GEN_9427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9429 = 8'hc9 == _match_key_qbytes_4_T ? phv_data_201 : _GEN_9428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9430 = 8'hca == _match_key_qbytes_4_T ? phv_data_202 : _GEN_9429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9431 = 8'hcb == _match_key_qbytes_4_T ? phv_data_203 : _GEN_9430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9432 = 8'hcc == _match_key_qbytes_4_T ? phv_data_204 : _GEN_9431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9433 = 8'hcd == _match_key_qbytes_4_T ? phv_data_205 : _GEN_9432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9434 = 8'hce == _match_key_qbytes_4_T ? phv_data_206 : _GEN_9433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9435 = 8'hcf == _match_key_qbytes_4_T ? phv_data_207 : _GEN_9434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9436 = 8'hd0 == _match_key_qbytes_4_T ? phv_data_208 : _GEN_9435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9437 = 8'hd1 == _match_key_qbytes_4_T ? phv_data_209 : _GEN_9436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9438 = 8'hd2 == _match_key_qbytes_4_T ? phv_data_210 : _GEN_9437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9439 = 8'hd3 == _match_key_qbytes_4_T ? phv_data_211 : _GEN_9438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9440 = 8'hd4 == _match_key_qbytes_4_T ? phv_data_212 : _GEN_9439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9441 = 8'hd5 == _match_key_qbytes_4_T ? phv_data_213 : _GEN_9440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9442 = 8'hd6 == _match_key_qbytes_4_T ? phv_data_214 : _GEN_9441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9443 = 8'hd7 == _match_key_qbytes_4_T ? phv_data_215 : _GEN_9442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9444 = 8'hd8 == _match_key_qbytes_4_T ? phv_data_216 : _GEN_9443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9445 = 8'hd9 == _match_key_qbytes_4_T ? phv_data_217 : _GEN_9444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9446 = 8'hda == _match_key_qbytes_4_T ? phv_data_218 : _GEN_9445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9447 = 8'hdb == _match_key_qbytes_4_T ? phv_data_219 : _GEN_9446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9448 = 8'hdc == _match_key_qbytes_4_T ? phv_data_220 : _GEN_9447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9449 = 8'hdd == _match_key_qbytes_4_T ? phv_data_221 : _GEN_9448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9450 = 8'hde == _match_key_qbytes_4_T ? phv_data_222 : _GEN_9449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9451 = 8'hdf == _match_key_qbytes_4_T ? phv_data_223 : _GEN_9450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9452 = 8'he0 == _match_key_qbytes_4_T ? phv_data_224 : _GEN_9451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9453 = 8'he1 == _match_key_qbytes_4_T ? phv_data_225 : _GEN_9452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9454 = 8'he2 == _match_key_qbytes_4_T ? phv_data_226 : _GEN_9453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9455 = 8'he3 == _match_key_qbytes_4_T ? phv_data_227 : _GEN_9454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9456 = 8'he4 == _match_key_qbytes_4_T ? phv_data_228 : _GEN_9455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9457 = 8'he5 == _match_key_qbytes_4_T ? phv_data_229 : _GEN_9456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9458 = 8'he6 == _match_key_qbytes_4_T ? phv_data_230 : _GEN_9457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9459 = 8'he7 == _match_key_qbytes_4_T ? phv_data_231 : _GEN_9458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9460 = 8'he8 == _match_key_qbytes_4_T ? phv_data_232 : _GEN_9459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9461 = 8'he9 == _match_key_qbytes_4_T ? phv_data_233 : _GEN_9460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9462 = 8'hea == _match_key_qbytes_4_T ? phv_data_234 : _GEN_9461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9463 = 8'heb == _match_key_qbytes_4_T ? phv_data_235 : _GEN_9462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9464 = 8'hec == _match_key_qbytes_4_T ? phv_data_236 : _GEN_9463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9465 = 8'hed == _match_key_qbytes_4_T ? phv_data_237 : _GEN_9464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9466 = 8'hee == _match_key_qbytes_4_T ? phv_data_238 : _GEN_9465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9467 = 8'hef == _match_key_qbytes_4_T ? phv_data_239 : _GEN_9466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9468 = 8'hf0 == _match_key_qbytes_4_T ? phv_data_240 : _GEN_9467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9469 = 8'hf1 == _match_key_qbytes_4_T ? phv_data_241 : _GEN_9468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9470 = 8'hf2 == _match_key_qbytes_4_T ? phv_data_242 : _GEN_9469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9471 = 8'hf3 == _match_key_qbytes_4_T ? phv_data_243 : _GEN_9470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9472 = 8'hf4 == _match_key_qbytes_4_T ? phv_data_244 : _GEN_9471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9473 = 8'hf5 == _match_key_qbytes_4_T ? phv_data_245 : _GEN_9472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9474 = 8'hf6 == _match_key_qbytes_4_T ? phv_data_246 : _GEN_9473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9475 = 8'hf7 == _match_key_qbytes_4_T ? phv_data_247 : _GEN_9474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9476 = 8'hf8 == _match_key_qbytes_4_T ? phv_data_248 : _GEN_9475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9477 = 8'hf9 == _match_key_qbytes_4_T ? phv_data_249 : _GEN_9476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9478 = 8'hfa == _match_key_qbytes_4_T ? phv_data_250 : _GEN_9477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9479 = 8'hfb == _match_key_qbytes_4_T ? phv_data_251 : _GEN_9478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9480 = 8'hfc == _match_key_qbytes_4_T ? phv_data_252 : _GEN_9479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9481 = 8'hfd == _match_key_qbytes_4_T ? phv_data_253 : _GEN_9480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9482 = 8'hfe == _match_key_qbytes_4_T ? phv_data_254 : _GEN_9481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9483 = 8'hff == _match_key_qbytes_4_T ? phv_data_255 : _GEN_9482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_16934 = {{1'd0}, _match_key_qbytes_4_T}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9484 = 9'h100 == _GEN_16934 ? phv_data_256 : _GEN_9483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9485 = 9'h101 == _GEN_16934 ? phv_data_257 : _GEN_9484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9486 = 9'h102 == _GEN_16934 ? phv_data_258 : _GEN_9485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9487 = 9'h103 == _GEN_16934 ? phv_data_259 : _GEN_9486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9488 = 9'h104 == _GEN_16934 ? phv_data_260 : _GEN_9487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9489 = 9'h105 == _GEN_16934 ? phv_data_261 : _GEN_9488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9490 = 9'h106 == _GEN_16934 ? phv_data_262 : _GEN_9489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9491 = 9'h107 == _GEN_16934 ? phv_data_263 : _GEN_9490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9492 = 9'h108 == _GEN_16934 ? phv_data_264 : _GEN_9491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9493 = 9'h109 == _GEN_16934 ? phv_data_265 : _GEN_9492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9494 = 9'h10a == _GEN_16934 ? phv_data_266 : _GEN_9493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9495 = 9'h10b == _GEN_16934 ? phv_data_267 : _GEN_9494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9496 = 9'h10c == _GEN_16934 ? phv_data_268 : _GEN_9495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9497 = 9'h10d == _GEN_16934 ? phv_data_269 : _GEN_9496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9498 = 9'h10e == _GEN_16934 ? phv_data_270 : _GEN_9497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9499 = 9'h10f == _GEN_16934 ? phv_data_271 : _GEN_9498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9500 = 9'h110 == _GEN_16934 ? phv_data_272 : _GEN_9499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9501 = 9'h111 == _GEN_16934 ? phv_data_273 : _GEN_9500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9502 = 9'h112 == _GEN_16934 ? phv_data_274 : _GEN_9501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9503 = 9'h113 == _GEN_16934 ? phv_data_275 : _GEN_9502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9504 = 9'h114 == _GEN_16934 ? phv_data_276 : _GEN_9503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9505 = 9'h115 == _GEN_16934 ? phv_data_277 : _GEN_9504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9506 = 9'h116 == _GEN_16934 ? phv_data_278 : _GEN_9505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9507 = 9'h117 == _GEN_16934 ? phv_data_279 : _GEN_9506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9508 = 9'h118 == _GEN_16934 ? phv_data_280 : _GEN_9507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9509 = 9'h119 == _GEN_16934 ? phv_data_281 : _GEN_9508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9510 = 9'h11a == _GEN_16934 ? phv_data_282 : _GEN_9509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9511 = 9'h11b == _GEN_16934 ? phv_data_283 : _GEN_9510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9512 = 9'h11c == _GEN_16934 ? phv_data_284 : _GEN_9511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9513 = 9'h11d == _GEN_16934 ? phv_data_285 : _GEN_9512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9514 = 9'h11e == _GEN_16934 ? phv_data_286 : _GEN_9513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9515 = 9'h11f == _GEN_16934 ? phv_data_287 : _GEN_9514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9516 = 9'h120 == _GEN_16934 ? phv_data_288 : _GEN_9515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9517 = 9'h121 == _GEN_16934 ? phv_data_289 : _GEN_9516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9518 = 9'h122 == _GEN_16934 ? phv_data_290 : _GEN_9517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9519 = 9'h123 == _GEN_16934 ? phv_data_291 : _GEN_9518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9520 = 9'h124 == _GEN_16934 ? phv_data_292 : _GEN_9519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9521 = 9'h125 == _GEN_16934 ? phv_data_293 : _GEN_9520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9522 = 9'h126 == _GEN_16934 ? phv_data_294 : _GEN_9521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9523 = 9'h127 == _GEN_16934 ? phv_data_295 : _GEN_9522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9524 = 9'h128 == _GEN_16934 ? phv_data_296 : _GEN_9523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9525 = 9'h129 == _GEN_16934 ? phv_data_297 : _GEN_9524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9526 = 9'h12a == _GEN_16934 ? phv_data_298 : _GEN_9525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9527 = 9'h12b == _GEN_16934 ? phv_data_299 : _GEN_9526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9528 = 9'h12c == _GEN_16934 ? phv_data_300 : _GEN_9527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9529 = 9'h12d == _GEN_16934 ? phv_data_301 : _GEN_9528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9530 = 9'h12e == _GEN_16934 ? phv_data_302 : _GEN_9529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9531 = 9'h12f == _GEN_16934 ? phv_data_303 : _GEN_9530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9532 = 9'h130 == _GEN_16934 ? phv_data_304 : _GEN_9531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9533 = 9'h131 == _GEN_16934 ? phv_data_305 : _GEN_9532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9534 = 9'h132 == _GEN_16934 ? phv_data_306 : _GEN_9533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9535 = 9'h133 == _GEN_16934 ? phv_data_307 : _GEN_9534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9536 = 9'h134 == _GEN_16934 ? phv_data_308 : _GEN_9535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9537 = 9'h135 == _GEN_16934 ? phv_data_309 : _GEN_9536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9538 = 9'h136 == _GEN_16934 ? phv_data_310 : _GEN_9537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9539 = 9'h137 == _GEN_16934 ? phv_data_311 : _GEN_9538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9540 = 9'h138 == _GEN_16934 ? phv_data_312 : _GEN_9539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9541 = 9'h139 == _GEN_16934 ? phv_data_313 : _GEN_9540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9542 = 9'h13a == _GEN_16934 ? phv_data_314 : _GEN_9541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9543 = 9'h13b == _GEN_16934 ? phv_data_315 : _GEN_9542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9544 = 9'h13c == _GEN_16934 ? phv_data_316 : _GEN_9543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9545 = 9'h13d == _GEN_16934 ? phv_data_317 : _GEN_9544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9546 = 9'h13e == _GEN_16934 ? phv_data_318 : _GEN_9545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9547 = 9'h13f == _GEN_16934 ? phv_data_319 : _GEN_9546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9548 = 9'h140 == _GEN_16934 ? phv_data_320 : _GEN_9547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9549 = 9'h141 == _GEN_16934 ? phv_data_321 : _GEN_9548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9550 = 9'h142 == _GEN_16934 ? phv_data_322 : _GEN_9549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9551 = 9'h143 == _GEN_16934 ? phv_data_323 : _GEN_9550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9552 = 9'h144 == _GEN_16934 ? phv_data_324 : _GEN_9551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9553 = 9'h145 == _GEN_16934 ? phv_data_325 : _GEN_9552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9554 = 9'h146 == _GEN_16934 ? phv_data_326 : _GEN_9553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9555 = 9'h147 == _GEN_16934 ? phv_data_327 : _GEN_9554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9556 = 9'h148 == _GEN_16934 ? phv_data_328 : _GEN_9555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9557 = 9'h149 == _GEN_16934 ? phv_data_329 : _GEN_9556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9558 = 9'h14a == _GEN_16934 ? phv_data_330 : _GEN_9557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9559 = 9'h14b == _GEN_16934 ? phv_data_331 : _GEN_9558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9560 = 9'h14c == _GEN_16934 ? phv_data_332 : _GEN_9559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9561 = 9'h14d == _GEN_16934 ? phv_data_333 : _GEN_9560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9562 = 9'h14e == _GEN_16934 ? phv_data_334 : _GEN_9561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9563 = 9'h14f == _GEN_16934 ? phv_data_335 : _GEN_9562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9564 = 9'h150 == _GEN_16934 ? phv_data_336 : _GEN_9563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9565 = 9'h151 == _GEN_16934 ? phv_data_337 : _GEN_9564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9566 = 9'h152 == _GEN_16934 ? phv_data_338 : _GEN_9565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9567 = 9'h153 == _GEN_16934 ? phv_data_339 : _GEN_9566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9568 = 9'h154 == _GEN_16934 ? phv_data_340 : _GEN_9567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9569 = 9'h155 == _GEN_16934 ? phv_data_341 : _GEN_9568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9570 = 9'h156 == _GEN_16934 ? phv_data_342 : _GEN_9569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9571 = 9'h157 == _GEN_16934 ? phv_data_343 : _GEN_9570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9572 = 9'h158 == _GEN_16934 ? phv_data_344 : _GEN_9571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9573 = 9'h159 == _GEN_16934 ? phv_data_345 : _GEN_9572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9574 = 9'h15a == _GEN_16934 ? phv_data_346 : _GEN_9573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9575 = 9'h15b == _GEN_16934 ? phv_data_347 : _GEN_9574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9576 = 9'h15c == _GEN_16934 ? phv_data_348 : _GEN_9575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9577 = 9'h15d == _GEN_16934 ? phv_data_349 : _GEN_9576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9578 = 9'h15e == _GEN_16934 ? phv_data_350 : _GEN_9577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9579 = 9'h15f == _GEN_16934 ? phv_data_351 : _GEN_9578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9580 = 9'h160 == _GEN_16934 ? phv_data_352 : _GEN_9579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9581 = 9'h161 == _GEN_16934 ? phv_data_353 : _GEN_9580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9582 = 9'h162 == _GEN_16934 ? phv_data_354 : _GEN_9581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9583 = 9'h163 == _GEN_16934 ? phv_data_355 : _GEN_9582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9584 = 9'h164 == _GEN_16934 ? phv_data_356 : _GEN_9583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9585 = 9'h165 == _GEN_16934 ? phv_data_357 : _GEN_9584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9586 = 9'h166 == _GEN_16934 ? phv_data_358 : _GEN_9585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9587 = 9'h167 == _GEN_16934 ? phv_data_359 : _GEN_9586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9588 = 9'h168 == _GEN_16934 ? phv_data_360 : _GEN_9587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9589 = 9'h169 == _GEN_16934 ? phv_data_361 : _GEN_9588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9590 = 9'h16a == _GEN_16934 ? phv_data_362 : _GEN_9589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9591 = 9'h16b == _GEN_16934 ? phv_data_363 : _GEN_9590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9592 = 9'h16c == _GEN_16934 ? phv_data_364 : _GEN_9591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9593 = 9'h16d == _GEN_16934 ? phv_data_365 : _GEN_9592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9594 = 9'h16e == _GEN_16934 ? phv_data_366 : _GEN_9593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9595 = 9'h16f == _GEN_16934 ? phv_data_367 : _GEN_9594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9596 = 9'h170 == _GEN_16934 ? phv_data_368 : _GEN_9595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9597 = 9'h171 == _GEN_16934 ? phv_data_369 : _GEN_9596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9598 = 9'h172 == _GEN_16934 ? phv_data_370 : _GEN_9597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9599 = 9'h173 == _GEN_16934 ? phv_data_371 : _GEN_9598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9600 = 9'h174 == _GEN_16934 ? phv_data_372 : _GEN_9599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9601 = 9'h175 == _GEN_16934 ? phv_data_373 : _GEN_9600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9602 = 9'h176 == _GEN_16934 ? phv_data_374 : _GEN_9601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9603 = 9'h177 == _GEN_16934 ? phv_data_375 : _GEN_9602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9604 = 9'h178 == _GEN_16934 ? phv_data_376 : _GEN_9603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9605 = 9'h179 == _GEN_16934 ? phv_data_377 : _GEN_9604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9606 = 9'h17a == _GEN_16934 ? phv_data_378 : _GEN_9605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9607 = 9'h17b == _GEN_16934 ? phv_data_379 : _GEN_9606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9608 = 9'h17c == _GEN_16934 ? phv_data_380 : _GEN_9607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9609 = 9'h17d == _GEN_16934 ? phv_data_381 : _GEN_9608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9610 = 9'h17e == _GEN_16934 ? phv_data_382 : _GEN_9609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9611 = 9'h17f == _GEN_16934 ? phv_data_383 : _GEN_9610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9612 = 9'h180 == _GEN_16934 ? phv_data_384 : _GEN_9611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9613 = 9'h181 == _GEN_16934 ? phv_data_385 : _GEN_9612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9614 = 9'h182 == _GEN_16934 ? phv_data_386 : _GEN_9613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9615 = 9'h183 == _GEN_16934 ? phv_data_387 : _GEN_9614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9616 = 9'h184 == _GEN_16934 ? phv_data_388 : _GEN_9615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9617 = 9'h185 == _GEN_16934 ? phv_data_389 : _GEN_9616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9618 = 9'h186 == _GEN_16934 ? phv_data_390 : _GEN_9617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9619 = 9'h187 == _GEN_16934 ? phv_data_391 : _GEN_9618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9620 = 9'h188 == _GEN_16934 ? phv_data_392 : _GEN_9619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9621 = 9'h189 == _GEN_16934 ? phv_data_393 : _GEN_9620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9622 = 9'h18a == _GEN_16934 ? phv_data_394 : _GEN_9621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9623 = 9'h18b == _GEN_16934 ? phv_data_395 : _GEN_9622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9624 = 9'h18c == _GEN_16934 ? phv_data_396 : _GEN_9623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9625 = 9'h18d == _GEN_16934 ? phv_data_397 : _GEN_9624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9626 = 9'h18e == _GEN_16934 ? phv_data_398 : _GEN_9625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9627 = 9'h18f == _GEN_16934 ? phv_data_399 : _GEN_9626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9628 = 9'h190 == _GEN_16934 ? phv_data_400 : _GEN_9627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9629 = 9'h191 == _GEN_16934 ? phv_data_401 : _GEN_9628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9630 = 9'h192 == _GEN_16934 ? phv_data_402 : _GEN_9629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9631 = 9'h193 == _GEN_16934 ? phv_data_403 : _GEN_9630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9632 = 9'h194 == _GEN_16934 ? phv_data_404 : _GEN_9631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9633 = 9'h195 == _GEN_16934 ? phv_data_405 : _GEN_9632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9634 = 9'h196 == _GEN_16934 ? phv_data_406 : _GEN_9633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9635 = 9'h197 == _GEN_16934 ? phv_data_407 : _GEN_9634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9636 = 9'h198 == _GEN_16934 ? phv_data_408 : _GEN_9635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9637 = 9'h199 == _GEN_16934 ? phv_data_409 : _GEN_9636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9638 = 9'h19a == _GEN_16934 ? phv_data_410 : _GEN_9637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9639 = 9'h19b == _GEN_16934 ? phv_data_411 : _GEN_9638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9640 = 9'h19c == _GEN_16934 ? phv_data_412 : _GEN_9639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9641 = 9'h19d == _GEN_16934 ? phv_data_413 : _GEN_9640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9642 = 9'h19e == _GEN_16934 ? phv_data_414 : _GEN_9641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9643 = 9'h19f == _GEN_16934 ? phv_data_415 : _GEN_9642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9644 = 9'h1a0 == _GEN_16934 ? phv_data_416 : _GEN_9643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9645 = 9'h1a1 == _GEN_16934 ? phv_data_417 : _GEN_9644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9646 = 9'h1a2 == _GEN_16934 ? phv_data_418 : _GEN_9645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9647 = 9'h1a3 == _GEN_16934 ? phv_data_419 : _GEN_9646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9648 = 9'h1a4 == _GEN_16934 ? phv_data_420 : _GEN_9647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9649 = 9'h1a5 == _GEN_16934 ? phv_data_421 : _GEN_9648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9650 = 9'h1a6 == _GEN_16934 ? phv_data_422 : _GEN_9649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9651 = 9'h1a7 == _GEN_16934 ? phv_data_423 : _GEN_9650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9652 = 9'h1a8 == _GEN_16934 ? phv_data_424 : _GEN_9651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9653 = 9'h1a9 == _GEN_16934 ? phv_data_425 : _GEN_9652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9654 = 9'h1aa == _GEN_16934 ? phv_data_426 : _GEN_9653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9655 = 9'h1ab == _GEN_16934 ? phv_data_427 : _GEN_9654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9656 = 9'h1ac == _GEN_16934 ? phv_data_428 : _GEN_9655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9657 = 9'h1ad == _GEN_16934 ? phv_data_429 : _GEN_9656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9658 = 9'h1ae == _GEN_16934 ? phv_data_430 : _GEN_9657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9659 = 9'h1af == _GEN_16934 ? phv_data_431 : _GEN_9658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9660 = 9'h1b0 == _GEN_16934 ? phv_data_432 : _GEN_9659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9661 = 9'h1b1 == _GEN_16934 ? phv_data_433 : _GEN_9660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9662 = 9'h1b2 == _GEN_16934 ? phv_data_434 : _GEN_9661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9663 = 9'h1b3 == _GEN_16934 ? phv_data_435 : _GEN_9662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9664 = 9'h1b4 == _GEN_16934 ? phv_data_436 : _GEN_9663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9665 = 9'h1b5 == _GEN_16934 ? phv_data_437 : _GEN_9664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9666 = 9'h1b6 == _GEN_16934 ? phv_data_438 : _GEN_9665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9667 = 9'h1b7 == _GEN_16934 ? phv_data_439 : _GEN_9666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9668 = 9'h1b8 == _GEN_16934 ? phv_data_440 : _GEN_9667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9669 = 9'h1b9 == _GEN_16934 ? phv_data_441 : _GEN_9668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9670 = 9'h1ba == _GEN_16934 ? phv_data_442 : _GEN_9669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9671 = 9'h1bb == _GEN_16934 ? phv_data_443 : _GEN_9670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9672 = 9'h1bc == _GEN_16934 ? phv_data_444 : _GEN_9671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9673 = 9'h1bd == _GEN_16934 ? phv_data_445 : _GEN_9672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9674 = 9'h1be == _GEN_16934 ? phv_data_446 : _GEN_9673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9675 = 9'h1bf == _GEN_16934 ? phv_data_447 : _GEN_9674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9676 = 9'h1c0 == _GEN_16934 ? phv_data_448 : _GEN_9675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9677 = 9'h1c1 == _GEN_16934 ? phv_data_449 : _GEN_9676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9678 = 9'h1c2 == _GEN_16934 ? phv_data_450 : _GEN_9677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9679 = 9'h1c3 == _GEN_16934 ? phv_data_451 : _GEN_9678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9680 = 9'h1c4 == _GEN_16934 ? phv_data_452 : _GEN_9679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9681 = 9'h1c5 == _GEN_16934 ? phv_data_453 : _GEN_9680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9682 = 9'h1c6 == _GEN_16934 ? phv_data_454 : _GEN_9681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9683 = 9'h1c7 == _GEN_16934 ? phv_data_455 : _GEN_9682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9684 = 9'h1c8 == _GEN_16934 ? phv_data_456 : _GEN_9683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9685 = 9'h1c9 == _GEN_16934 ? phv_data_457 : _GEN_9684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9686 = 9'h1ca == _GEN_16934 ? phv_data_458 : _GEN_9685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9687 = 9'h1cb == _GEN_16934 ? phv_data_459 : _GEN_9686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9688 = 9'h1cc == _GEN_16934 ? phv_data_460 : _GEN_9687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9689 = 9'h1cd == _GEN_16934 ? phv_data_461 : _GEN_9688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9690 = 9'h1ce == _GEN_16934 ? phv_data_462 : _GEN_9689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9691 = 9'h1cf == _GEN_16934 ? phv_data_463 : _GEN_9690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9692 = 9'h1d0 == _GEN_16934 ? phv_data_464 : _GEN_9691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9693 = 9'h1d1 == _GEN_16934 ? phv_data_465 : _GEN_9692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9694 = 9'h1d2 == _GEN_16934 ? phv_data_466 : _GEN_9693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9695 = 9'h1d3 == _GEN_16934 ? phv_data_467 : _GEN_9694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9696 = 9'h1d4 == _GEN_16934 ? phv_data_468 : _GEN_9695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9697 = 9'h1d5 == _GEN_16934 ? phv_data_469 : _GEN_9696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9698 = 9'h1d6 == _GEN_16934 ? phv_data_470 : _GEN_9697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9699 = 9'h1d7 == _GEN_16934 ? phv_data_471 : _GEN_9698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9700 = 9'h1d8 == _GEN_16934 ? phv_data_472 : _GEN_9699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9701 = 9'h1d9 == _GEN_16934 ? phv_data_473 : _GEN_9700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9702 = 9'h1da == _GEN_16934 ? phv_data_474 : _GEN_9701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9703 = 9'h1db == _GEN_16934 ? phv_data_475 : _GEN_9702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9704 = 9'h1dc == _GEN_16934 ? phv_data_476 : _GEN_9703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9705 = 9'h1dd == _GEN_16934 ? phv_data_477 : _GEN_9704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9706 = 9'h1de == _GEN_16934 ? phv_data_478 : _GEN_9705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9707 = 9'h1df == _GEN_16934 ? phv_data_479 : _GEN_9706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9708 = 9'h1e0 == _GEN_16934 ? phv_data_480 : _GEN_9707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9709 = 9'h1e1 == _GEN_16934 ? phv_data_481 : _GEN_9708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9710 = 9'h1e2 == _GEN_16934 ? phv_data_482 : _GEN_9709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9711 = 9'h1e3 == _GEN_16934 ? phv_data_483 : _GEN_9710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9712 = 9'h1e4 == _GEN_16934 ? phv_data_484 : _GEN_9711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9713 = 9'h1e5 == _GEN_16934 ? phv_data_485 : _GEN_9712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9714 = 9'h1e6 == _GEN_16934 ? phv_data_486 : _GEN_9713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9715 = 9'h1e7 == _GEN_16934 ? phv_data_487 : _GEN_9714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9716 = 9'h1e8 == _GEN_16934 ? phv_data_488 : _GEN_9715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9717 = 9'h1e9 == _GEN_16934 ? phv_data_489 : _GEN_9716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9718 = 9'h1ea == _GEN_16934 ? phv_data_490 : _GEN_9717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9719 = 9'h1eb == _GEN_16934 ? phv_data_491 : _GEN_9718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9720 = 9'h1ec == _GEN_16934 ? phv_data_492 : _GEN_9719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9721 = 9'h1ed == _GEN_16934 ? phv_data_493 : _GEN_9720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9722 = 9'h1ee == _GEN_16934 ? phv_data_494 : _GEN_9721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9723 = 9'h1ef == _GEN_16934 ? phv_data_495 : _GEN_9722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9724 = 9'h1f0 == _GEN_16934 ? phv_data_496 : _GEN_9723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9725 = 9'h1f1 == _GEN_16934 ? phv_data_497 : _GEN_9724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9726 = 9'h1f2 == _GEN_16934 ? phv_data_498 : _GEN_9725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9727 = 9'h1f3 == _GEN_16934 ? phv_data_499 : _GEN_9726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9728 = 9'h1f4 == _GEN_16934 ? phv_data_500 : _GEN_9727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9729 = 9'h1f5 == _GEN_16934 ? phv_data_501 : _GEN_9728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9730 = 9'h1f6 == _GEN_16934 ? phv_data_502 : _GEN_9729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9731 = 9'h1f7 == _GEN_16934 ? phv_data_503 : _GEN_9730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9732 = 9'h1f8 == _GEN_16934 ? phv_data_504 : _GEN_9731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9733 = 9'h1f9 == _GEN_16934 ? phv_data_505 : _GEN_9732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9734 = 9'h1fa == _GEN_16934 ? phv_data_506 : _GEN_9733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9735 = 9'h1fb == _GEN_16934 ? phv_data_507 : _GEN_9734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9736 = 9'h1fc == _GEN_16934 ? phv_data_508 : _GEN_9735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9737 = 9'h1fd == _GEN_16934 ? phv_data_509 : _GEN_9736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9738 = 9'h1fe == _GEN_16934 ? phv_data_510 : _GEN_9737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9739 = 9'h1ff == _GEN_16934 ? phv_data_511 : _GEN_9738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9741 = 8'h1 == _match_key_qbytes_4_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9742 = 8'h2 == _match_key_qbytes_4_T_1 ? phv_data_2 : _GEN_9741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9743 = 8'h3 == _match_key_qbytes_4_T_1 ? phv_data_3 : _GEN_9742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9744 = 8'h4 == _match_key_qbytes_4_T_1 ? phv_data_4 : _GEN_9743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9745 = 8'h5 == _match_key_qbytes_4_T_1 ? phv_data_5 : _GEN_9744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9746 = 8'h6 == _match_key_qbytes_4_T_1 ? phv_data_6 : _GEN_9745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9747 = 8'h7 == _match_key_qbytes_4_T_1 ? phv_data_7 : _GEN_9746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9748 = 8'h8 == _match_key_qbytes_4_T_1 ? phv_data_8 : _GEN_9747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9749 = 8'h9 == _match_key_qbytes_4_T_1 ? phv_data_9 : _GEN_9748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9750 = 8'ha == _match_key_qbytes_4_T_1 ? phv_data_10 : _GEN_9749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9751 = 8'hb == _match_key_qbytes_4_T_1 ? phv_data_11 : _GEN_9750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9752 = 8'hc == _match_key_qbytes_4_T_1 ? phv_data_12 : _GEN_9751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9753 = 8'hd == _match_key_qbytes_4_T_1 ? phv_data_13 : _GEN_9752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9754 = 8'he == _match_key_qbytes_4_T_1 ? phv_data_14 : _GEN_9753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9755 = 8'hf == _match_key_qbytes_4_T_1 ? phv_data_15 : _GEN_9754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9756 = 8'h10 == _match_key_qbytes_4_T_1 ? phv_data_16 : _GEN_9755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9757 = 8'h11 == _match_key_qbytes_4_T_1 ? phv_data_17 : _GEN_9756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9758 = 8'h12 == _match_key_qbytes_4_T_1 ? phv_data_18 : _GEN_9757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9759 = 8'h13 == _match_key_qbytes_4_T_1 ? phv_data_19 : _GEN_9758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9760 = 8'h14 == _match_key_qbytes_4_T_1 ? phv_data_20 : _GEN_9759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9761 = 8'h15 == _match_key_qbytes_4_T_1 ? phv_data_21 : _GEN_9760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9762 = 8'h16 == _match_key_qbytes_4_T_1 ? phv_data_22 : _GEN_9761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9763 = 8'h17 == _match_key_qbytes_4_T_1 ? phv_data_23 : _GEN_9762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9764 = 8'h18 == _match_key_qbytes_4_T_1 ? phv_data_24 : _GEN_9763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9765 = 8'h19 == _match_key_qbytes_4_T_1 ? phv_data_25 : _GEN_9764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9766 = 8'h1a == _match_key_qbytes_4_T_1 ? phv_data_26 : _GEN_9765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9767 = 8'h1b == _match_key_qbytes_4_T_1 ? phv_data_27 : _GEN_9766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9768 = 8'h1c == _match_key_qbytes_4_T_1 ? phv_data_28 : _GEN_9767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9769 = 8'h1d == _match_key_qbytes_4_T_1 ? phv_data_29 : _GEN_9768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9770 = 8'h1e == _match_key_qbytes_4_T_1 ? phv_data_30 : _GEN_9769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9771 = 8'h1f == _match_key_qbytes_4_T_1 ? phv_data_31 : _GEN_9770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9772 = 8'h20 == _match_key_qbytes_4_T_1 ? phv_data_32 : _GEN_9771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9773 = 8'h21 == _match_key_qbytes_4_T_1 ? phv_data_33 : _GEN_9772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9774 = 8'h22 == _match_key_qbytes_4_T_1 ? phv_data_34 : _GEN_9773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9775 = 8'h23 == _match_key_qbytes_4_T_1 ? phv_data_35 : _GEN_9774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9776 = 8'h24 == _match_key_qbytes_4_T_1 ? phv_data_36 : _GEN_9775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9777 = 8'h25 == _match_key_qbytes_4_T_1 ? phv_data_37 : _GEN_9776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9778 = 8'h26 == _match_key_qbytes_4_T_1 ? phv_data_38 : _GEN_9777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9779 = 8'h27 == _match_key_qbytes_4_T_1 ? phv_data_39 : _GEN_9778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9780 = 8'h28 == _match_key_qbytes_4_T_1 ? phv_data_40 : _GEN_9779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9781 = 8'h29 == _match_key_qbytes_4_T_1 ? phv_data_41 : _GEN_9780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9782 = 8'h2a == _match_key_qbytes_4_T_1 ? phv_data_42 : _GEN_9781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9783 = 8'h2b == _match_key_qbytes_4_T_1 ? phv_data_43 : _GEN_9782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9784 = 8'h2c == _match_key_qbytes_4_T_1 ? phv_data_44 : _GEN_9783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9785 = 8'h2d == _match_key_qbytes_4_T_1 ? phv_data_45 : _GEN_9784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9786 = 8'h2e == _match_key_qbytes_4_T_1 ? phv_data_46 : _GEN_9785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9787 = 8'h2f == _match_key_qbytes_4_T_1 ? phv_data_47 : _GEN_9786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9788 = 8'h30 == _match_key_qbytes_4_T_1 ? phv_data_48 : _GEN_9787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9789 = 8'h31 == _match_key_qbytes_4_T_1 ? phv_data_49 : _GEN_9788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9790 = 8'h32 == _match_key_qbytes_4_T_1 ? phv_data_50 : _GEN_9789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9791 = 8'h33 == _match_key_qbytes_4_T_1 ? phv_data_51 : _GEN_9790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9792 = 8'h34 == _match_key_qbytes_4_T_1 ? phv_data_52 : _GEN_9791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9793 = 8'h35 == _match_key_qbytes_4_T_1 ? phv_data_53 : _GEN_9792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9794 = 8'h36 == _match_key_qbytes_4_T_1 ? phv_data_54 : _GEN_9793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9795 = 8'h37 == _match_key_qbytes_4_T_1 ? phv_data_55 : _GEN_9794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9796 = 8'h38 == _match_key_qbytes_4_T_1 ? phv_data_56 : _GEN_9795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9797 = 8'h39 == _match_key_qbytes_4_T_1 ? phv_data_57 : _GEN_9796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9798 = 8'h3a == _match_key_qbytes_4_T_1 ? phv_data_58 : _GEN_9797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9799 = 8'h3b == _match_key_qbytes_4_T_1 ? phv_data_59 : _GEN_9798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9800 = 8'h3c == _match_key_qbytes_4_T_1 ? phv_data_60 : _GEN_9799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9801 = 8'h3d == _match_key_qbytes_4_T_1 ? phv_data_61 : _GEN_9800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9802 = 8'h3e == _match_key_qbytes_4_T_1 ? phv_data_62 : _GEN_9801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9803 = 8'h3f == _match_key_qbytes_4_T_1 ? phv_data_63 : _GEN_9802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9804 = 8'h40 == _match_key_qbytes_4_T_1 ? phv_data_64 : _GEN_9803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9805 = 8'h41 == _match_key_qbytes_4_T_1 ? phv_data_65 : _GEN_9804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9806 = 8'h42 == _match_key_qbytes_4_T_1 ? phv_data_66 : _GEN_9805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9807 = 8'h43 == _match_key_qbytes_4_T_1 ? phv_data_67 : _GEN_9806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9808 = 8'h44 == _match_key_qbytes_4_T_1 ? phv_data_68 : _GEN_9807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9809 = 8'h45 == _match_key_qbytes_4_T_1 ? phv_data_69 : _GEN_9808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9810 = 8'h46 == _match_key_qbytes_4_T_1 ? phv_data_70 : _GEN_9809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9811 = 8'h47 == _match_key_qbytes_4_T_1 ? phv_data_71 : _GEN_9810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9812 = 8'h48 == _match_key_qbytes_4_T_1 ? phv_data_72 : _GEN_9811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9813 = 8'h49 == _match_key_qbytes_4_T_1 ? phv_data_73 : _GEN_9812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9814 = 8'h4a == _match_key_qbytes_4_T_1 ? phv_data_74 : _GEN_9813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9815 = 8'h4b == _match_key_qbytes_4_T_1 ? phv_data_75 : _GEN_9814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9816 = 8'h4c == _match_key_qbytes_4_T_1 ? phv_data_76 : _GEN_9815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9817 = 8'h4d == _match_key_qbytes_4_T_1 ? phv_data_77 : _GEN_9816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9818 = 8'h4e == _match_key_qbytes_4_T_1 ? phv_data_78 : _GEN_9817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9819 = 8'h4f == _match_key_qbytes_4_T_1 ? phv_data_79 : _GEN_9818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9820 = 8'h50 == _match_key_qbytes_4_T_1 ? phv_data_80 : _GEN_9819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9821 = 8'h51 == _match_key_qbytes_4_T_1 ? phv_data_81 : _GEN_9820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9822 = 8'h52 == _match_key_qbytes_4_T_1 ? phv_data_82 : _GEN_9821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9823 = 8'h53 == _match_key_qbytes_4_T_1 ? phv_data_83 : _GEN_9822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9824 = 8'h54 == _match_key_qbytes_4_T_1 ? phv_data_84 : _GEN_9823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9825 = 8'h55 == _match_key_qbytes_4_T_1 ? phv_data_85 : _GEN_9824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9826 = 8'h56 == _match_key_qbytes_4_T_1 ? phv_data_86 : _GEN_9825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9827 = 8'h57 == _match_key_qbytes_4_T_1 ? phv_data_87 : _GEN_9826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9828 = 8'h58 == _match_key_qbytes_4_T_1 ? phv_data_88 : _GEN_9827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9829 = 8'h59 == _match_key_qbytes_4_T_1 ? phv_data_89 : _GEN_9828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9830 = 8'h5a == _match_key_qbytes_4_T_1 ? phv_data_90 : _GEN_9829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9831 = 8'h5b == _match_key_qbytes_4_T_1 ? phv_data_91 : _GEN_9830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9832 = 8'h5c == _match_key_qbytes_4_T_1 ? phv_data_92 : _GEN_9831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9833 = 8'h5d == _match_key_qbytes_4_T_1 ? phv_data_93 : _GEN_9832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9834 = 8'h5e == _match_key_qbytes_4_T_1 ? phv_data_94 : _GEN_9833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9835 = 8'h5f == _match_key_qbytes_4_T_1 ? phv_data_95 : _GEN_9834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9836 = 8'h60 == _match_key_qbytes_4_T_1 ? phv_data_96 : _GEN_9835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9837 = 8'h61 == _match_key_qbytes_4_T_1 ? phv_data_97 : _GEN_9836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9838 = 8'h62 == _match_key_qbytes_4_T_1 ? phv_data_98 : _GEN_9837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9839 = 8'h63 == _match_key_qbytes_4_T_1 ? phv_data_99 : _GEN_9838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9840 = 8'h64 == _match_key_qbytes_4_T_1 ? phv_data_100 : _GEN_9839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9841 = 8'h65 == _match_key_qbytes_4_T_1 ? phv_data_101 : _GEN_9840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9842 = 8'h66 == _match_key_qbytes_4_T_1 ? phv_data_102 : _GEN_9841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9843 = 8'h67 == _match_key_qbytes_4_T_1 ? phv_data_103 : _GEN_9842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9844 = 8'h68 == _match_key_qbytes_4_T_1 ? phv_data_104 : _GEN_9843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9845 = 8'h69 == _match_key_qbytes_4_T_1 ? phv_data_105 : _GEN_9844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9846 = 8'h6a == _match_key_qbytes_4_T_1 ? phv_data_106 : _GEN_9845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9847 = 8'h6b == _match_key_qbytes_4_T_1 ? phv_data_107 : _GEN_9846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9848 = 8'h6c == _match_key_qbytes_4_T_1 ? phv_data_108 : _GEN_9847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9849 = 8'h6d == _match_key_qbytes_4_T_1 ? phv_data_109 : _GEN_9848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9850 = 8'h6e == _match_key_qbytes_4_T_1 ? phv_data_110 : _GEN_9849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9851 = 8'h6f == _match_key_qbytes_4_T_1 ? phv_data_111 : _GEN_9850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9852 = 8'h70 == _match_key_qbytes_4_T_1 ? phv_data_112 : _GEN_9851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9853 = 8'h71 == _match_key_qbytes_4_T_1 ? phv_data_113 : _GEN_9852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9854 = 8'h72 == _match_key_qbytes_4_T_1 ? phv_data_114 : _GEN_9853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9855 = 8'h73 == _match_key_qbytes_4_T_1 ? phv_data_115 : _GEN_9854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9856 = 8'h74 == _match_key_qbytes_4_T_1 ? phv_data_116 : _GEN_9855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9857 = 8'h75 == _match_key_qbytes_4_T_1 ? phv_data_117 : _GEN_9856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9858 = 8'h76 == _match_key_qbytes_4_T_1 ? phv_data_118 : _GEN_9857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9859 = 8'h77 == _match_key_qbytes_4_T_1 ? phv_data_119 : _GEN_9858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9860 = 8'h78 == _match_key_qbytes_4_T_1 ? phv_data_120 : _GEN_9859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9861 = 8'h79 == _match_key_qbytes_4_T_1 ? phv_data_121 : _GEN_9860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9862 = 8'h7a == _match_key_qbytes_4_T_1 ? phv_data_122 : _GEN_9861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9863 = 8'h7b == _match_key_qbytes_4_T_1 ? phv_data_123 : _GEN_9862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9864 = 8'h7c == _match_key_qbytes_4_T_1 ? phv_data_124 : _GEN_9863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9865 = 8'h7d == _match_key_qbytes_4_T_1 ? phv_data_125 : _GEN_9864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9866 = 8'h7e == _match_key_qbytes_4_T_1 ? phv_data_126 : _GEN_9865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9867 = 8'h7f == _match_key_qbytes_4_T_1 ? phv_data_127 : _GEN_9866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9868 = 8'h80 == _match_key_qbytes_4_T_1 ? phv_data_128 : _GEN_9867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9869 = 8'h81 == _match_key_qbytes_4_T_1 ? phv_data_129 : _GEN_9868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9870 = 8'h82 == _match_key_qbytes_4_T_1 ? phv_data_130 : _GEN_9869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9871 = 8'h83 == _match_key_qbytes_4_T_1 ? phv_data_131 : _GEN_9870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9872 = 8'h84 == _match_key_qbytes_4_T_1 ? phv_data_132 : _GEN_9871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9873 = 8'h85 == _match_key_qbytes_4_T_1 ? phv_data_133 : _GEN_9872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9874 = 8'h86 == _match_key_qbytes_4_T_1 ? phv_data_134 : _GEN_9873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9875 = 8'h87 == _match_key_qbytes_4_T_1 ? phv_data_135 : _GEN_9874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9876 = 8'h88 == _match_key_qbytes_4_T_1 ? phv_data_136 : _GEN_9875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9877 = 8'h89 == _match_key_qbytes_4_T_1 ? phv_data_137 : _GEN_9876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9878 = 8'h8a == _match_key_qbytes_4_T_1 ? phv_data_138 : _GEN_9877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9879 = 8'h8b == _match_key_qbytes_4_T_1 ? phv_data_139 : _GEN_9878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9880 = 8'h8c == _match_key_qbytes_4_T_1 ? phv_data_140 : _GEN_9879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9881 = 8'h8d == _match_key_qbytes_4_T_1 ? phv_data_141 : _GEN_9880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9882 = 8'h8e == _match_key_qbytes_4_T_1 ? phv_data_142 : _GEN_9881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9883 = 8'h8f == _match_key_qbytes_4_T_1 ? phv_data_143 : _GEN_9882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9884 = 8'h90 == _match_key_qbytes_4_T_1 ? phv_data_144 : _GEN_9883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9885 = 8'h91 == _match_key_qbytes_4_T_1 ? phv_data_145 : _GEN_9884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9886 = 8'h92 == _match_key_qbytes_4_T_1 ? phv_data_146 : _GEN_9885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9887 = 8'h93 == _match_key_qbytes_4_T_1 ? phv_data_147 : _GEN_9886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9888 = 8'h94 == _match_key_qbytes_4_T_1 ? phv_data_148 : _GEN_9887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9889 = 8'h95 == _match_key_qbytes_4_T_1 ? phv_data_149 : _GEN_9888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9890 = 8'h96 == _match_key_qbytes_4_T_1 ? phv_data_150 : _GEN_9889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9891 = 8'h97 == _match_key_qbytes_4_T_1 ? phv_data_151 : _GEN_9890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9892 = 8'h98 == _match_key_qbytes_4_T_1 ? phv_data_152 : _GEN_9891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9893 = 8'h99 == _match_key_qbytes_4_T_1 ? phv_data_153 : _GEN_9892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9894 = 8'h9a == _match_key_qbytes_4_T_1 ? phv_data_154 : _GEN_9893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9895 = 8'h9b == _match_key_qbytes_4_T_1 ? phv_data_155 : _GEN_9894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9896 = 8'h9c == _match_key_qbytes_4_T_1 ? phv_data_156 : _GEN_9895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9897 = 8'h9d == _match_key_qbytes_4_T_1 ? phv_data_157 : _GEN_9896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9898 = 8'h9e == _match_key_qbytes_4_T_1 ? phv_data_158 : _GEN_9897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9899 = 8'h9f == _match_key_qbytes_4_T_1 ? phv_data_159 : _GEN_9898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9900 = 8'ha0 == _match_key_qbytes_4_T_1 ? phv_data_160 : _GEN_9899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9901 = 8'ha1 == _match_key_qbytes_4_T_1 ? phv_data_161 : _GEN_9900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9902 = 8'ha2 == _match_key_qbytes_4_T_1 ? phv_data_162 : _GEN_9901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9903 = 8'ha3 == _match_key_qbytes_4_T_1 ? phv_data_163 : _GEN_9902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9904 = 8'ha4 == _match_key_qbytes_4_T_1 ? phv_data_164 : _GEN_9903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9905 = 8'ha5 == _match_key_qbytes_4_T_1 ? phv_data_165 : _GEN_9904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9906 = 8'ha6 == _match_key_qbytes_4_T_1 ? phv_data_166 : _GEN_9905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9907 = 8'ha7 == _match_key_qbytes_4_T_1 ? phv_data_167 : _GEN_9906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9908 = 8'ha8 == _match_key_qbytes_4_T_1 ? phv_data_168 : _GEN_9907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9909 = 8'ha9 == _match_key_qbytes_4_T_1 ? phv_data_169 : _GEN_9908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9910 = 8'haa == _match_key_qbytes_4_T_1 ? phv_data_170 : _GEN_9909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9911 = 8'hab == _match_key_qbytes_4_T_1 ? phv_data_171 : _GEN_9910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9912 = 8'hac == _match_key_qbytes_4_T_1 ? phv_data_172 : _GEN_9911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9913 = 8'had == _match_key_qbytes_4_T_1 ? phv_data_173 : _GEN_9912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9914 = 8'hae == _match_key_qbytes_4_T_1 ? phv_data_174 : _GEN_9913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9915 = 8'haf == _match_key_qbytes_4_T_1 ? phv_data_175 : _GEN_9914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9916 = 8'hb0 == _match_key_qbytes_4_T_1 ? phv_data_176 : _GEN_9915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9917 = 8'hb1 == _match_key_qbytes_4_T_1 ? phv_data_177 : _GEN_9916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9918 = 8'hb2 == _match_key_qbytes_4_T_1 ? phv_data_178 : _GEN_9917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9919 = 8'hb3 == _match_key_qbytes_4_T_1 ? phv_data_179 : _GEN_9918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9920 = 8'hb4 == _match_key_qbytes_4_T_1 ? phv_data_180 : _GEN_9919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9921 = 8'hb5 == _match_key_qbytes_4_T_1 ? phv_data_181 : _GEN_9920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9922 = 8'hb6 == _match_key_qbytes_4_T_1 ? phv_data_182 : _GEN_9921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9923 = 8'hb7 == _match_key_qbytes_4_T_1 ? phv_data_183 : _GEN_9922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9924 = 8'hb8 == _match_key_qbytes_4_T_1 ? phv_data_184 : _GEN_9923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9925 = 8'hb9 == _match_key_qbytes_4_T_1 ? phv_data_185 : _GEN_9924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9926 = 8'hba == _match_key_qbytes_4_T_1 ? phv_data_186 : _GEN_9925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9927 = 8'hbb == _match_key_qbytes_4_T_1 ? phv_data_187 : _GEN_9926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9928 = 8'hbc == _match_key_qbytes_4_T_1 ? phv_data_188 : _GEN_9927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9929 = 8'hbd == _match_key_qbytes_4_T_1 ? phv_data_189 : _GEN_9928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9930 = 8'hbe == _match_key_qbytes_4_T_1 ? phv_data_190 : _GEN_9929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9931 = 8'hbf == _match_key_qbytes_4_T_1 ? phv_data_191 : _GEN_9930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9932 = 8'hc0 == _match_key_qbytes_4_T_1 ? phv_data_192 : _GEN_9931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9933 = 8'hc1 == _match_key_qbytes_4_T_1 ? phv_data_193 : _GEN_9932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9934 = 8'hc2 == _match_key_qbytes_4_T_1 ? phv_data_194 : _GEN_9933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9935 = 8'hc3 == _match_key_qbytes_4_T_1 ? phv_data_195 : _GEN_9934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9936 = 8'hc4 == _match_key_qbytes_4_T_1 ? phv_data_196 : _GEN_9935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9937 = 8'hc5 == _match_key_qbytes_4_T_1 ? phv_data_197 : _GEN_9936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9938 = 8'hc6 == _match_key_qbytes_4_T_1 ? phv_data_198 : _GEN_9937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9939 = 8'hc7 == _match_key_qbytes_4_T_1 ? phv_data_199 : _GEN_9938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9940 = 8'hc8 == _match_key_qbytes_4_T_1 ? phv_data_200 : _GEN_9939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9941 = 8'hc9 == _match_key_qbytes_4_T_1 ? phv_data_201 : _GEN_9940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9942 = 8'hca == _match_key_qbytes_4_T_1 ? phv_data_202 : _GEN_9941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9943 = 8'hcb == _match_key_qbytes_4_T_1 ? phv_data_203 : _GEN_9942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9944 = 8'hcc == _match_key_qbytes_4_T_1 ? phv_data_204 : _GEN_9943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9945 = 8'hcd == _match_key_qbytes_4_T_1 ? phv_data_205 : _GEN_9944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9946 = 8'hce == _match_key_qbytes_4_T_1 ? phv_data_206 : _GEN_9945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9947 = 8'hcf == _match_key_qbytes_4_T_1 ? phv_data_207 : _GEN_9946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9948 = 8'hd0 == _match_key_qbytes_4_T_1 ? phv_data_208 : _GEN_9947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9949 = 8'hd1 == _match_key_qbytes_4_T_1 ? phv_data_209 : _GEN_9948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9950 = 8'hd2 == _match_key_qbytes_4_T_1 ? phv_data_210 : _GEN_9949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9951 = 8'hd3 == _match_key_qbytes_4_T_1 ? phv_data_211 : _GEN_9950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9952 = 8'hd4 == _match_key_qbytes_4_T_1 ? phv_data_212 : _GEN_9951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9953 = 8'hd5 == _match_key_qbytes_4_T_1 ? phv_data_213 : _GEN_9952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9954 = 8'hd6 == _match_key_qbytes_4_T_1 ? phv_data_214 : _GEN_9953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9955 = 8'hd7 == _match_key_qbytes_4_T_1 ? phv_data_215 : _GEN_9954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9956 = 8'hd8 == _match_key_qbytes_4_T_1 ? phv_data_216 : _GEN_9955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9957 = 8'hd9 == _match_key_qbytes_4_T_1 ? phv_data_217 : _GEN_9956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9958 = 8'hda == _match_key_qbytes_4_T_1 ? phv_data_218 : _GEN_9957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9959 = 8'hdb == _match_key_qbytes_4_T_1 ? phv_data_219 : _GEN_9958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9960 = 8'hdc == _match_key_qbytes_4_T_1 ? phv_data_220 : _GEN_9959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9961 = 8'hdd == _match_key_qbytes_4_T_1 ? phv_data_221 : _GEN_9960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9962 = 8'hde == _match_key_qbytes_4_T_1 ? phv_data_222 : _GEN_9961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9963 = 8'hdf == _match_key_qbytes_4_T_1 ? phv_data_223 : _GEN_9962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9964 = 8'he0 == _match_key_qbytes_4_T_1 ? phv_data_224 : _GEN_9963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9965 = 8'he1 == _match_key_qbytes_4_T_1 ? phv_data_225 : _GEN_9964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9966 = 8'he2 == _match_key_qbytes_4_T_1 ? phv_data_226 : _GEN_9965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9967 = 8'he3 == _match_key_qbytes_4_T_1 ? phv_data_227 : _GEN_9966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9968 = 8'he4 == _match_key_qbytes_4_T_1 ? phv_data_228 : _GEN_9967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9969 = 8'he5 == _match_key_qbytes_4_T_1 ? phv_data_229 : _GEN_9968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9970 = 8'he6 == _match_key_qbytes_4_T_1 ? phv_data_230 : _GEN_9969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9971 = 8'he7 == _match_key_qbytes_4_T_1 ? phv_data_231 : _GEN_9970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9972 = 8'he8 == _match_key_qbytes_4_T_1 ? phv_data_232 : _GEN_9971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9973 = 8'he9 == _match_key_qbytes_4_T_1 ? phv_data_233 : _GEN_9972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9974 = 8'hea == _match_key_qbytes_4_T_1 ? phv_data_234 : _GEN_9973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9975 = 8'heb == _match_key_qbytes_4_T_1 ? phv_data_235 : _GEN_9974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9976 = 8'hec == _match_key_qbytes_4_T_1 ? phv_data_236 : _GEN_9975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9977 = 8'hed == _match_key_qbytes_4_T_1 ? phv_data_237 : _GEN_9976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9978 = 8'hee == _match_key_qbytes_4_T_1 ? phv_data_238 : _GEN_9977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9979 = 8'hef == _match_key_qbytes_4_T_1 ? phv_data_239 : _GEN_9978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9980 = 8'hf0 == _match_key_qbytes_4_T_1 ? phv_data_240 : _GEN_9979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9981 = 8'hf1 == _match_key_qbytes_4_T_1 ? phv_data_241 : _GEN_9980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9982 = 8'hf2 == _match_key_qbytes_4_T_1 ? phv_data_242 : _GEN_9981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9983 = 8'hf3 == _match_key_qbytes_4_T_1 ? phv_data_243 : _GEN_9982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9984 = 8'hf4 == _match_key_qbytes_4_T_1 ? phv_data_244 : _GEN_9983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9985 = 8'hf5 == _match_key_qbytes_4_T_1 ? phv_data_245 : _GEN_9984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9986 = 8'hf6 == _match_key_qbytes_4_T_1 ? phv_data_246 : _GEN_9985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9987 = 8'hf7 == _match_key_qbytes_4_T_1 ? phv_data_247 : _GEN_9986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9988 = 8'hf8 == _match_key_qbytes_4_T_1 ? phv_data_248 : _GEN_9987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9989 = 8'hf9 == _match_key_qbytes_4_T_1 ? phv_data_249 : _GEN_9988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9990 = 8'hfa == _match_key_qbytes_4_T_1 ? phv_data_250 : _GEN_9989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9991 = 8'hfb == _match_key_qbytes_4_T_1 ? phv_data_251 : _GEN_9990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9992 = 8'hfc == _match_key_qbytes_4_T_1 ? phv_data_252 : _GEN_9991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9993 = 8'hfd == _match_key_qbytes_4_T_1 ? phv_data_253 : _GEN_9992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9994 = 8'hfe == _match_key_qbytes_4_T_1 ? phv_data_254 : _GEN_9993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9995 = 8'hff == _match_key_qbytes_4_T_1 ? phv_data_255 : _GEN_9994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_17190 = {{1'd0}, _match_key_qbytes_4_T_1}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9996 = 9'h100 == _GEN_17190 ? phv_data_256 : _GEN_9995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9997 = 9'h101 == _GEN_17190 ? phv_data_257 : _GEN_9996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9998 = 9'h102 == _GEN_17190 ? phv_data_258 : _GEN_9997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9999 = 9'h103 == _GEN_17190 ? phv_data_259 : _GEN_9998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10000 = 9'h104 == _GEN_17190 ? phv_data_260 : _GEN_9999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10001 = 9'h105 == _GEN_17190 ? phv_data_261 : _GEN_10000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10002 = 9'h106 == _GEN_17190 ? phv_data_262 : _GEN_10001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10003 = 9'h107 == _GEN_17190 ? phv_data_263 : _GEN_10002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10004 = 9'h108 == _GEN_17190 ? phv_data_264 : _GEN_10003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10005 = 9'h109 == _GEN_17190 ? phv_data_265 : _GEN_10004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10006 = 9'h10a == _GEN_17190 ? phv_data_266 : _GEN_10005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10007 = 9'h10b == _GEN_17190 ? phv_data_267 : _GEN_10006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10008 = 9'h10c == _GEN_17190 ? phv_data_268 : _GEN_10007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10009 = 9'h10d == _GEN_17190 ? phv_data_269 : _GEN_10008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10010 = 9'h10e == _GEN_17190 ? phv_data_270 : _GEN_10009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10011 = 9'h10f == _GEN_17190 ? phv_data_271 : _GEN_10010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10012 = 9'h110 == _GEN_17190 ? phv_data_272 : _GEN_10011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10013 = 9'h111 == _GEN_17190 ? phv_data_273 : _GEN_10012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10014 = 9'h112 == _GEN_17190 ? phv_data_274 : _GEN_10013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10015 = 9'h113 == _GEN_17190 ? phv_data_275 : _GEN_10014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10016 = 9'h114 == _GEN_17190 ? phv_data_276 : _GEN_10015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10017 = 9'h115 == _GEN_17190 ? phv_data_277 : _GEN_10016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10018 = 9'h116 == _GEN_17190 ? phv_data_278 : _GEN_10017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10019 = 9'h117 == _GEN_17190 ? phv_data_279 : _GEN_10018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10020 = 9'h118 == _GEN_17190 ? phv_data_280 : _GEN_10019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10021 = 9'h119 == _GEN_17190 ? phv_data_281 : _GEN_10020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10022 = 9'h11a == _GEN_17190 ? phv_data_282 : _GEN_10021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10023 = 9'h11b == _GEN_17190 ? phv_data_283 : _GEN_10022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10024 = 9'h11c == _GEN_17190 ? phv_data_284 : _GEN_10023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10025 = 9'h11d == _GEN_17190 ? phv_data_285 : _GEN_10024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10026 = 9'h11e == _GEN_17190 ? phv_data_286 : _GEN_10025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10027 = 9'h11f == _GEN_17190 ? phv_data_287 : _GEN_10026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10028 = 9'h120 == _GEN_17190 ? phv_data_288 : _GEN_10027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10029 = 9'h121 == _GEN_17190 ? phv_data_289 : _GEN_10028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10030 = 9'h122 == _GEN_17190 ? phv_data_290 : _GEN_10029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10031 = 9'h123 == _GEN_17190 ? phv_data_291 : _GEN_10030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10032 = 9'h124 == _GEN_17190 ? phv_data_292 : _GEN_10031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10033 = 9'h125 == _GEN_17190 ? phv_data_293 : _GEN_10032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10034 = 9'h126 == _GEN_17190 ? phv_data_294 : _GEN_10033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10035 = 9'h127 == _GEN_17190 ? phv_data_295 : _GEN_10034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10036 = 9'h128 == _GEN_17190 ? phv_data_296 : _GEN_10035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10037 = 9'h129 == _GEN_17190 ? phv_data_297 : _GEN_10036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10038 = 9'h12a == _GEN_17190 ? phv_data_298 : _GEN_10037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10039 = 9'h12b == _GEN_17190 ? phv_data_299 : _GEN_10038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10040 = 9'h12c == _GEN_17190 ? phv_data_300 : _GEN_10039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10041 = 9'h12d == _GEN_17190 ? phv_data_301 : _GEN_10040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10042 = 9'h12e == _GEN_17190 ? phv_data_302 : _GEN_10041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10043 = 9'h12f == _GEN_17190 ? phv_data_303 : _GEN_10042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10044 = 9'h130 == _GEN_17190 ? phv_data_304 : _GEN_10043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10045 = 9'h131 == _GEN_17190 ? phv_data_305 : _GEN_10044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10046 = 9'h132 == _GEN_17190 ? phv_data_306 : _GEN_10045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10047 = 9'h133 == _GEN_17190 ? phv_data_307 : _GEN_10046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10048 = 9'h134 == _GEN_17190 ? phv_data_308 : _GEN_10047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10049 = 9'h135 == _GEN_17190 ? phv_data_309 : _GEN_10048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10050 = 9'h136 == _GEN_17190 ? phv_data_310 : _GEN_10049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10051 = 9'h137 == _GEN_17190 ? phv_data_311 : _GEN_10050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10052 = 9'h138 == _GEN_17190 ? phv_data_312 : _GEN_10051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10053 = 9'h139 == _GEN_17190 ? phv_data_313 : _GEN_10052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10054 = 9'h13a == _GEN_17190 ? phv_data_314 : _GEN_10053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10055 = 9'h13b == _GEN_17190 ? phv_data_315 : _GEN_10054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10056 = 9'h13c == _GEN_17190 ? phv_data_316 : _GEN_10055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10057 = 9'h13d == _GEN_17190 ? phv_data_317 : _GEN_10056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10058 = 9'h13e == _GEN_17190 ? phv_data_318 : _GEN_10057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10059 = 9'h13f == _GEN_17190 ? phv_data_319 : _GEN_10058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10060 = 9'h140 == _GEN_17190 ? phv_data_320 : _GEN_10059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10061 = 9'h141 == _GEN_17190 ? phv_data_321 : _GEN_10060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10062 = 9'h142 == _GEN_17190 ? phv_data_322 : _GEN_10061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10063 = 9'h143 == _GEN_17190 ? phv_data_323 : _GEN_10062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10064 = 9'h144 == _GEN_17190 ? phv_data_324 : _GEN_10063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10065 = 9'h145 == _GEN_17190 ? phv_data_325 : _GEN_10064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10066 = 9'h146 == _GEN_17190 ? phv_data_326 : _GEN_10065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10067 = 9'h147 == _GEN_17190 ? phv_data_327 : _GEN_10066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10068 = 9'h148 == _GEN_17190 ? phv_data_328 : _GEN_10067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10069 = 9'h149 == _GEN_17190 ? phv_data_329 : _GEN_10068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10070 = 9'h14a == _GEN_17190 ? phv_data_330 : _GEN_10069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10071 = 9'h14b == _GEN_17190 ? phv_data_331 : _GEN_10070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10072 = 9'h14c == _GEN_17190 ? phv_data_332 : _GEN_10071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10073 = 9'h14d == _GEN_17190 ? phv_data_333 : _GEN_10072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10074 = 9'h14e == _GEN_17190 ? phv_data_334 : _GEN_10073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10075 = 9'h14f == _GEN_17190 ? phv_data_335 : _GEN_10074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10076 = 9'h150 == _GEN_17190 ? phv_data_336 : _GEN_10075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10077 = 9'h151 == _GEN_17190 ? phv_data_337 : _GEN_10076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10078 = 9'h152 == _GEN_17190 ? phv_data_338 : _GEN_10077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10079 = 9'h153 == _GEN_17190 ? phv_data_339 : _GEN_10078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10080 = 9'h154 == _GEN_17190 ? phv_data_340 : _GEN_10079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10081 = 9'h155 == _GEN_17190 ? phv_data_341 : _GEN_10080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10082 = 9'h156 == _GEN_17190 ? phv_data_342 : _GEN_10081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10083 = 9'h157 == _GEN_17190 ? phv_data_343 : _GEN_10082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10084 = 9'h158 == _GEN_17190 ? phv_data_344 : _GEN_10083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10085 = 9'h159 == _GEN_17190 ? phv_data_345 : _GEN_10084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10086 = 9'h15a == _GEN_17190 ? phv_data_346 : _GEN_10085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10087 = 9'h15b == _GEN_17190 ? phv_data_347 : _GEN_10086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10088 = 9'h15c == _GEN_17190 ? phv_data_348 : _GEN_10087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10089 = 9'h15d == _GEN_17190 ? phv_data_349 : _GEN_10088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10090 = 9'h15e == _GEN_17190 ? phv_data_350 : _GEN_10089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10091 = 9'h15f == _GEN_17190 ? phv_data_351 : _GEN_10090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10092 = 9'h160 == _GEN_17190 ? phv_data_352 : _GEN_10091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10093 = 9'h161 == _GEN_17190 ? phv_data_353 : _GEN_10092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10094 = 9'h162 == _GEN_17190 ? phv_data_354 : _GEN_10093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10095 = 9'h163 == _GEN_17190 ? phv_data_355 : _GEN_10094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10096 = 9'h164 == _GEN_17190 ? phv_data_356 : _GEN_10095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10097 = 9'h165 == _GEN_17190 ? phv_data_357 : _GEN_10096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10098 = 9'h166 == _GEN_17190 ? phv_data_358 : _GEN_10097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10099 = 9'h167 == _GEN_17190 ? phv_data_359 : _GEN_10098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10100 = 9'h168 == _GEN_17190 ? phv_data_360 : _GEN_10099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10101 = 9'h169 == _GEN_17190 ? phv_data_361 : _GEN_10100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10102 = 9'h16a == _GEN_17190 ? phv_data_362 : _GEN_10101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10103 = 9'h16b == _GEN_17190 ? phv_data_363 : _GEN_10102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10104 = 9'h16c == _GEN_17190 ? phv_data_364 : _GEN_10103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10105 = 9'h16d == _GEN_17190 ? phv_data_365 : _GEN_10104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10106 = 9'h16e == _GEN_17190 ? phv_data_366 : _GEN_10105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10107 = 9'h16f == _GEN_17190 ? phv_data_367 : _GEN_10106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10108 = 9'h170 == _GEN_17190 ? phv_data_368 : _GEN_10107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10109 = 9'h171 == _GEN_17190 ? phv_data_369 : _GEN_10108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10110 = 9'h172 == _GEN_17190 ? phv_data_370 : _GEN_10109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10111 = 9'h173 == _GEN_17190 ? phv_data_371 : _GEN_10110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10112 = 9'h174 == _GEN_17190 ? phv_data_372 : _GEN_10111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10113 = 9'h175 == _GEN_17190 ? phv_data_373 : _GEN_10112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10114 = 9'h176 == _GEN_17190 ? phv_data_374 : _GEN_10113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10115 = 9'h177 == _GEN_17190 ? phv_data_375 : _GEN_10114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10116 = 9'h178 == _GEN_17190 ? phv_data_376 : _GEN_10115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10117 = 9'h179 == _GEN_17190 ? phv_data_377 : _GEN_10116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10118 = 9'h17a == _GEN_17190 ? phv_data_378 : _GEN_10117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10119 = 9'h17b == _GEN_17190 ? phv_data_379 : _GEN_10118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10120 = 9'h17c == _GEN_17190 ? phv_data_380 : _GEN_10119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10121 = 9'h17d == _GEN_17190 ? phv_data_381 : _GEN_10120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10122 = 9'h17e == _GEN_17190 ? phv_data_382 : _GEN_10121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10123 = 9'h17f == _GEN_17190 ? phv_data_383 : _GEN_10122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10124 = 9'h180 == _GEN_17190 ? phv_data_384 : _GEN_10123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10125 = 9'h181 == _GEN_17190 ? phv_data_385 : _GEN_10124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10126 = 9'h182 == _GEN_17190 ? phv_data_386 : _GEN_10125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10127 = 9'h183 == _GEN_17190 ? phv_data_387 : _GEN_10126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10128 = 9'h184 == _GEN_17190 ? phv_data_388 : _GEN_10127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10129 = 9'h185 == _GEN_17190 ? phv_data_389 : _GEN_10128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10130 = 9'h186 == _GEN_17190 ? phv_data_390 : _GEN_10129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10131 = 9'h187 == _GEN_17190 ? phv_data_391 : _GEN_10130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10132 = 9'h188 == _GEN_17190 ? phv_data_392 : _GEN_10131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10133 = 9'h189 == _GEN_17190 ? phv_data_393 : _GEN_10132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10134 = 9'h18a == _GEN_17190 ? phv_data_394 : _GEN_10133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10135 = 9'h18b == _GEN_17190 ? phv_data_395 : _GEN_10134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10136 = 9'h18c == _GEN_17190 ? phv_data_396 : _GEN_10135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10137 = 9'h18d == _GEN_17190 ? phv_data_397 : _GEN_10136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10138 = 9'h18e == _GEN_17190 ? phv_data_398 : _GEN_10137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10139 = 9'h18f == _GEN_17190 ? phv_data_399 : _GEN_10138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10140 = 9'h190 == _GEN_17190 ? phv_data_400 : _GEN_10139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10141 = 9'h191 == _GEN_17190 ? phv_data_401 : _GEN_10140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10142 = 9'h192 == _GEN_17190 ? phv_data_402 : _GEN_10141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10143 = 9'h193 == _GEN_17190 ? phv_data_403 : _GEN_10142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10144 = 9'h194 == _GEN_17190 ? phv_data_404 : _GEN_10143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10145 = 9'h195 == _GEN_17190 ? phv_data_405 : _GEN_10144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10146 = 9'h196 == _GEN_17190 ? phv_data_406 : _GEN_10145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10147 = 9'h197 == _GEN_17190 ? phv_data_407 : _GEN_10146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10148 = 9'h198 == _GEN_17190 ? phv_data_408 : _GEN_10147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10149 = 9'h199 == _GEN_17190 ? phv_data_409 : _GEN_10148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10150 = 9'h19a == _GEN_17190 ? phv_data_410 : _GEN_10149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10151 = 9'h19b == _GEN_17190 ? phv_data_411 : _GEN_10150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10152 = 9'h19c == _GEN_17190 ? phv_data_412 : _GEN_10151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10153 = 9'h19d == _GEN_17190 ? phv_data_413 : _GEN_10152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10154 = 9'h19e == _GEN_17190 ? phv_data_414 : _GEN_10153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10155 = 9'h19f == _GEN_17190 ? phv_data_415 : _GEN_10154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10156 = 9'h1a0 == _GEN_17190 ? phv_data_416 : _GEN_10155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10157 = 9'h1a1 == _GEN_17190 ? phv_data_417 : _GEN_10156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10158 = 9'h1a2 == _GEN_17190 ? phv_data_418 : _GEN_10157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10159 = 9'h1a3 == _GEN_17190 ? phv_data_419 : _GEN_10158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10160 = 9'h1a4 == _GEN_17190 ? phv_data_420 : _GEN_10159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10161 = 9'h1a5 == _GEN_17190 ? phv_data_421 : _GEN_10160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10162 = 9'h1a6 == _GEN_17190 ? phv_data_422 : _GEN_10161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10163 = 9'h1a7 == _GEN_17190 ? phv_data_423 : _GEN_10162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10164 = 9'h1a8 == _GEN_17190 ? phv_data_424 : _GEN_10163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10165 = 9'h1a9 == _GEN_17190 ? phv_data_425 : _GEN_10164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10166 = 9'h1aa == _GEN_17190 ? phv_data_426 : _GEN_10165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10167 = 9'h1ab == _GEN_17190 ? phv_data_427 : _GEN_10166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10168 = 9'h1ac == _GEN_17190 ? phv_data_428 : _GEN_10167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10169 = 9'h1ad == _GEN_17190 ? phv_data_429 : _GEN_10168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10170 = 9'h1ae == _GEN_17190 ? phv_data_430 : _GEN_10169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10171 = 9'h1af == _GEN_17190 ? phv_data_431 : _GEN_10170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10172 = 9'h1b0 == _GEN_17190 ? phv_data_432 : _GEN_10171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10173 = 9'h1b1 == _GEN_17190 ? phv_data_433 : _GEN_10172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10174 = 9'h1b2 == _GEN_17190 ? phv_data_434 : _GEN_10173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10175 = 9'h1b3 == _GEN_17190 ? phv_data_435 : _GEN_10174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10176 = 9'h1b4 == _GEN_17190 ? phv_data_436 : _GEN_10175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10177 = 9'h1b5 == _GEN_17190 ? phv_data_437 : _GEN_10176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10178 = 9'h1b6 == _GEN_17190 ? phv_data_438 : _GEN_10177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10179 = 9'h1b7 == _GEN_17190 ? phv_data_439 : _GEN_10178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10180 = 9'h1b8 == _GEN_17190 ? phv_data_440 : _GEN_10179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10181 = 9'h1b9 == _GEN_17190 ? phv_data_441 : _GEN_10180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10182 = 9'h1ba == _GEN_17190 ? phv_data_442 : _GEN_10181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10183 = 9'h1bb == _GEN_17190 ? phv_data_443 : _GEN_10182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10184 = 9'h1bc == _GEN_17190 ? phv_data_444 : _GEN_10183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10185 = 9'h1bd == _GEN_17190 ? phv_data_445 : _GEN_10184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10186 = 9'h1be == _GEN_17190 ? phv_data_446 : _GEN_10185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10187 = 9'h1bf == _GEN_17190 ? phv_data_447 : _GEN_10186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10188 = 9'h1c0 == _GEN_17190 ? phv_data_448 : _GEN_10187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10189 = 9'h1c1 == _GEN_17190 ? phv_data_449 : _GEN_10188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10190 = 9'h1c2 == _GEN_17190 ? phv_data_450 : _GEN_10189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10191 = 9'h1c3 == _GEN_17190 ? phv_data_451 : _GEN_10190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10192 = 9'h1c4 == _GEN_17190 ? phv_data_452 : _GEN_10191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10193 = 9'h1c5 == _GEN_17190 ? phv_data_453 : _GEN_10192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10194 = 9'h1c6 == _GEN_17190 ? phv_data_454 : _GEN_10193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10195 = 9'h1c7 == _GEN_17190 ? phv_data_455 : _GEN_10194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10196 = 9'h1c8 == _GEN_17190 ? phv_data_456 : _GEN_10195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10197 = 9'h1c9 == _GEN_17190 ? phv_data_457 : _GEN_10196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10198 = 9'h1ca == _GEN_17190 ? phv_data_458 : _GEN_10197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10199 = 9'h1cb == _GEN_17190 ? phv_data_459 : _GEN_10198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10200 = 9'h1cc == _GEN_17190 ? phv_data_460 : _GEN_10199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10201 = 9'h1cd == _GEN_17190 ? phv_data_461 : _GEN_10200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10202 = 9'h1ce == _GEN_17190 ? phv_data_462 : _GEN_10201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10203 = 9'h1cf == _GEN_17190 ? phv_data_463 : _GEN_10202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10204 = 9'h1d0 == _GEN_17190 ? phv_data_464 : _GEN_10203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10205 = 9'h1d1 == _GEN_17190 ? phv_data_465 : _GEN_10204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10206 = 9'h1d2 == _GEN_17190 ? phv_data_466 : _GEN_10205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10207 = 9'h1d3 == _GEN_17190 ? phv_data_467 : _GEN_10206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10208 = 9'h1d4 == _GEN_17190 ? phv_data_468 : _GEN_10207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10209 = 9'h1d5 == _GEN_17190 ? phv_data_469 : _GEN_10208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10210 = 9'h1d6 == _GEN_17190 ? phv_data_470 : _GEN_10209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10211 = 9'h1d7 == _GEN_17190 ? phv_data_471 : _GEN_10210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10212 = 9'h1d8 == _GEN_17190 ? phv_data_472 : _GEN_10211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10213 = 9'h1d9 == _GEN_17190 ? phv_data_473 : _GEN_10212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10214 = 9'h1da == _GEN_17190 ? phv_data_474 : _GEN_10213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10215 = 9'h1db == _GEN_17190 ? phv_data_475 : _GEN_10214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10216 = 9'h1dc == _GEN_17190 ? phv_data_476 : _GEN_10215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10217 = 9'h1dd == _GEN_17190 ? phv_data_477 : _GEN_10216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10218 = 9'h1de == _GEN_17190 ? phv_data_478 : _GEN_10217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10219 = 9'h1df == _GEN_17190 ? phv_data_479 : _GEN_10218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10220 = 9'h1e0 == _GEN_17190 ? phv_data_480 : _GEN_10219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10221 = 9'h1e1 == _GEN_17190 ? phv_data_481 : _GEN_10220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10222 = 9'h1e2 == _GEN_17190 ? phv_data_482 : _GEN_10221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10223 = 9'h1e3 == _GEN_17190 ? phv_data_483 : _GEN_10222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10224 = 9'h1e4 == _GEN_17190 ? phv_data_484 : _GEN_10223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10225 = 9'h1e5 == _GEN_17190 ? phv_data_485 : _GEN_10224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10226 = 9'h1e6 == _GEN_17190 ? phv_data_486 : _GEN_10225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10227 = 9'h1e7 == _GEN_17190 ? phv_data_487 : _GEN_10226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10228 = 9'h1e8 == _GEN_17190 ? phv_data_488 : _GEN_10227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10229 = 9'h1e9 == _GEN_17190 ? phv_data_489 : _GEN_10228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10230 = 9'h1ea == _GEN_17190 ? phv_data_490 : _GEN_10229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10231 = 9'h1eb == _GEN_17190 ? phv_data_491 : _GEN_10230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10232 = 9'h1ec == _GEN_17190 ? phv_data_492 : _GEN_10231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10233 = 9'h1ed == _GEN_17190 ? phv_data_493 : _GEN_10232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10234 = 9'h1ee == _GEN_17190 ? phv_data_494 : _GEN_10233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10235 = 9'h1ef == _GEN_17190 ? phv_data_495 : _GEN_10234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10236 = 9'h1f0 == _GEN_17190 ? phv_data_496 : _GEN_10235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10237 = 9'h1f1 == _GEN_17190 ? phv_data_497 : _GEN_10236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10238 = 9'h1f2 == _GEN_17190 ? phv_data_498 : _GEN_10237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10239 = 9'h1f3 == _GEN_17190 ? phv_data_499 : _GEN_10238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10240 = 9'h1f4 == _GEN_17190 ? phv_data_500 : _GEN_10239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10241 = 9'h1f5 == _GEN_17190 ? phv_data_501 : _GEN_10240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10242 = 9'h1f6 == _GEN_17190 ? phv_data_502 : _GEN_10241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10243 = 9'h1f7 == _GEN_17190 ? phv_data_503 : _GEN_10242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10244 = 9'h1f8 == _GEN_17190 ? phv_data_504 : _GEN_10243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10245 = 9'h1f9 == _GEN_17190 ? phv_data_505 : _GEN_10244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10246 = 9'h1fa == _GEN_17190 ? phv_data_506 : _GEN_10245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10247 = 9'h1fb == _GEN_17190 ? phv_data_507 : _GEN_10246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10248 = 9'h1fc == _GEN_17190 ? phv_data_508 : _GEN_10247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10249 = 9'h1fd == _GEN_17190 ? phv_data_509 : _GEN_10248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10250 = 9'h1fe == _GEN_17190 ? phv_data_510 : _GEN_10249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10251 = 9'h1ff == _GEN_17190 ? phv_data_511 : _GEN_10250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_4_T_3 = {_GEN_9739,_GEN_10251,_GEN_8715,_GEN_9227}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_4 = local_offset_4 < end_offset ? _match_key_qbytes_4_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  wire [7:0] local_offset_5 = 8'h14 + read_key_offset; // @[matcher.scala 87:77]
  wire [5:0] match_key_qbytes_5_hi = local_offset_5[7:2]; // @[matcher.scala 91:54]
  wire [7:0] _match_key_qbytes_5_T = {match_key_qbytes_5_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_5_T_1 = {match_key_qbytes_5_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _match_key_qbytes_5_T_2 = {match_key_qbytes_5_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_10254 = 8'h1 == _match_key_qbytes_5_T_2 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10255 = 8'h2 == _match_key_qbytes_5_T_2 ? phv_data_2 : _GEN_10254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10256 = 8'h3 == _match_key_qbytes_5_T_2 ? phv_data_3 : _GEN_10255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10257 = 8'h4 == _match_key_qbytes_5_T_2 ? phv_data_4 : _GEN_10256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10258 = 8'h5 == _match_key_qbytes_5_T_2 ? phv_data_5 : _GEN_10257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10259 = 8'h6 == _match_key_qbytes_5_T_2 ? phv_data_6 : _GEN_10258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10260 = 8'h7 == _match_key_qbytes_5_T_2 ? phv_data_7 : _GEN_10259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10261 = 8'h8 == _match_key_qbytes_5_T_2 ? phv_data_8 : _GEN_10260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10262 = 8'h9 == _match_key_qbytes_5_T_2 ? phv_data_9 : _GEN_10261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10263 = 8'ha == _match_key_qbytes_5_T_2 ? phv_data_10 : _GEN_10262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10264 = 8'hb == _match_key_qbytes_5_T_2 ? phv_data_11 : _GEN_10263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10265 = 8'hc == _match_key_qbytes_5_T_2 ? phv_data_12 : _GEN_10264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10266 = 8'hd == _match_key_qbytes_5_T_2 ? phv_data_13 : _GEN_10265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10267 = 8'he == _match_key_qbytes_5_T_2 ? phv_data_14 : _GEN_10266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10268 = 8'hf == _match_key_qbytes_5_T_2 ? phv_data_15 : _GEN_10267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10269 = 8'h10 == _match_key_qbytes_5_T_2 ? phv_data_16 : _GEN_10268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10270 = 8'h11 == _match_key_qbytes_5_T_2 ? phv_data_17 : _GEN_10269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10271 = 8'h12 == _match_key_qbytes_5_T_2 ? phv_data_18 : _GEN_10270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10272 = 8'h13 == _match_key_qbytes_5_T_2 ? phv_data_19 : _GEN_10271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10273 = 8'h14 == _match_key_qbytes_5_T_2 ? phv_data_20 : _GEN_10272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10274 = 8'h15 == _match_key_qbytes_5_T_2 ? phv_data_21 : _GEN_10273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10275 = 8'h16 == _match_key_qbytes_5_T_2 ? phv_data_22 : _GEN_10274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10276 = 8'h17 == _match_key_qbytes_5_T_2 ? phv_data_23 : _GEN_10275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10277 = 8'h18 == _match_key_qbytes_5_T_2 ? phv_data_24 : _GEN_10276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10278 = 8'h19 == _match_key_qbytes_5_T_2 ? phv_data_25 : _GEN_10277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10279 = 8'h1a == _match_key_qbytes_5_T_2 ? phv_data_26 : _GEN_10278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10280 = 8'h1b == _match_key_qbytes_5_T_2 ? phv_data_27 : _GEN_10279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10281 = 8'h1c == _match_key_qbytes_5_T_2 ? phv_data_28 : _GEN_10280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10282 = 8'h1d == _match_key_qbytes_5_T_2 ? phv_data_29 : _GEN_10281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10283 = 8'h1e == _match_key_qbytes_5_T_2 ? phv_data_30 : _GEN_10282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10284 = 8'h1f == _match_key_qbytes_5_T_2 ? phv_data_31 : _GEN_10283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10285 = 8'h20 == _match_key_qbytes_5_T_2 ? phv_data_32 : _GEN_10284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10286 = 8'h21 == _match_key_qbytes_5_T_2 ? phv_data_33 : _GEN_10285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10287 = 8'h22 == _match_key_qbytes_5_T_2 ? phv_data_34 : _GEN_10286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10288 = 8'h23 == _match_key_qbytes_5_T_2 ? phv_data_35 : _GEN_10287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10289 = 8'h24 == _match_key_qbytes_5_T_2 ? phv_data_36 : _GEN_10288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10290 = 8'h25 == _match_key_qbytes_5_T_2 ? phv_data_37 : _GEN_10289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10291 = 8'h26 == _match_key_qbytes_5_T_2 ? phv_data_38 : _GEN_10290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10292 = 8'h27 == _match_key_qbytes_5_T_2 ? phv_data_39 : _GEN_10291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10293 = 8'h28 == _match_key_qbytes_5_T_2 ? phv_data_40 : _GEN_10292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10294 = 8'h29 == _match_key_qbytes_5_T_2 ? phv_data_41 : _GEN_10293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10295 = 8'h2a == _match_key_qbytes_5_T_2 ? phv_data_42 : _GEN_10294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10296 = 8'h2b == _match_key_qbytes_5_T_2 ? phv_data_43 : _GEN_10295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10297 = 8'h2c == _match_key_qbytes_5_T_2 ? phv_data_44 : _GEN_10296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10298 = 8'h2d == _match_key_qbytes_5_T_2 ? phv_data_45 : _GEN_10297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10299 = 8'h2e == _match_key_qbytes_5_T_2 ? phv_data_46 : _GEN_10298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10300 = 8'h2f == _match_key_qbytes_5_T_2 ? phv_data_47 : _GEN_10299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10301 = 8'h30 == _match_key_qbytes_5_T_2 ? phv_data_48 : _GEN_10300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10302 = 8'h31 == _match_key_qbytes_5_T_2 ? phv_data_49 : _GEN_10301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10303 = 8'h32 == _match_key_qbytes_5_T_2 ? phv_data_50 : _GEN_10302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10304 = 8'h33 == _match_key_qbytes_5_T_2 ? phv_data_51 : _GEN_10303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10305 = 8'h34 == _match_key_qbytes_5_T_2 ? phv_data_52 : _GEN_10304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10306 = 8'h35 == _match_key_qbytes_5_T_2 ? phv_data_53 : _GEN_10305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10307 = 8'h36 == _match_key_qbytes_5_T_2 ? phv_data_54 : _GEN_10306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10308 = 8'h37 == _match_key_qbytes_5_T_2 ? phv_data_55 : _GEN_10307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10309 = 8'h38 == _match_key_qbytes_5_T_2 ? phv_data_56 : _GEN_10308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10310 = 8'h39 == _match_key_qbytes_5_T_2 ? phv_data_57 : _GEN_10309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10311 = 8'h3a == _match_key_qbytes_5_T_2 ? phv_data_58 : _GEN_10310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10312 = 8'h3b == _match_key_qbytes_5_T_2 ? phv_data_59 : _GEN_10311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10313 = 8'h3c == _match_key_qbytes_5_T_2 ? phv_data_60 : _GEN_10312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10314 = 8'h3d == _match_key_qbytes_5_T_2 ? phv_data_61 : _GEN_10313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10315 = 8'h3e == _match_key_qbytes_5_T_2 ? phv_data_62 : _GEN_10314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10316 = 8'h3f == _match_key_qbytes_5_T_2 ? phv_data_63 : _GEN_10315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10317 = 8'h40 == _match_key_qbytes_5_T_2 ? phv_data_64 : _GEN_10316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10318 = 8'h41 == _match_key_qbytes_5_T_2 ? phv_data_65 : _GEN_10317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10319 = 8'h42 == _match_key_qbytes_5_T_2 ? phv_data_66 : _GEN_10318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10320 = 8'h43 == _match_key_qbytes_5_T_2 ? phv_data_67 : _GEN_10319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10321 = 8'h44 == _match_key_qbytes_5_T_2 ? phv_data_68 : _GEN_10320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10322 = 8'h45 == _match_key_qbytes_5_T_2 ? phv_data_69 : _GEN_10321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10323 = 8'h46 == _match_key_qbytes_5_T_2 ? phv_data_70 : _GEN_10322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10324 = 8'h47 == _match_key_qbytes_5_T_2 ? phv_data_71 : _GEN_10323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10325 = 8'h48 == _match_key_qbytes_5_T_2 ? phv_data_72 : _GEN_10324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10326 = 8'h49 == _match_key_qbytes_5_T_2 ? phv_data_73 : _GEN_10325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10327 = 8'h4a == _match_key_qbytes_5_T_2 ? phv_data_74 : _GEN_10326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10328 = 8'h4b == _match_key_qbytes_5_T_2 ? phv_data_75 : _GEN_10327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10329 = 8'h4c == _match_key_qbytes_5_T_2 ? phv_data_76 : _GEN_10328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10330 = 8'h4d == _match_key_qbytes_5_T_2 ? phv_data_77 : _GEN_10329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10331 = 8'h4e == _match_key_qbytes_5_T_2 ? phv_data_78 : _GEN_10330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10332 = 8'h4f == _match_key_qbytes_5_T_2 ? phv_data_79 : _GEN_10331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10333 = 8'h50 == _match_key_qbytes_5_T_2 ? phv_data_80 : _GEN_10332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10334 = 8'h51 == _match_key_qbytes_5_T_2 ? phv_data_81 : _GEN_10333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10335 = 8'h52 == _match_key_qbytes_5_T_2 ? phv_data_82 : _GEN_10334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10336 = 8'h53 == _match_key_qbytes_5_T_2 ? phv_data_83 : _GEN_10335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10337 = 8'h54 == _match_key_qbytes_5_T_2 ? phv_data_84 : _GEN_10336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10338 = 8'h55 == _match_key_qbytes_5_T_2 ? phv_data_85 : _GEN_10337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10339 = 8'h56 == _match_key_qbytes_5_T_2 ? phv_data_86 : _GEN_10338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10340 = 8'h57 == _match_key_qbytes_5_T_2 ? phv_data_87 : _GEN_10339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10341 = 8'h58 == _match_key_qbytes_5_T_2 ? phv_data_88 : _GEN_10340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10342 = 8'h59 == _match_key_qbytes_5_T_2 ? phv_data_89 : _GEN_10341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10343 = 8'h5a == _match_key_qbytes_5_T_2 ? phv_data_90 : _GEN_10342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10344 = 8'h5b == _match_key_qbytes_5_T_2 ? phv_data_91 : _GEN_10343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10345 = 8'h5c == _match_key_qbytes_5_T_2 ? phv_data_92 : _GEN_10344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10346 = 8'h5d == _match_key_qbytes_5_T_2 ? phv_data_93 : _GEN_10345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10347 = 8'h5e == _match_key_qbytes_5_T_2 ? phv_data_94 : _GEN_10346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10348 = 8'h5f == _match_key_qbytes_5_T_2 ? phv_data_95 : _GEN_10347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10349 = 8'h60 == _match_key_qbytes_5_T_2 ? phv_data_96 : _GEN_10348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10350 = 8'h61 == _match_key_qbytes_5_T_2 ? phv_data_97 : _GEN_10349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10351 = 8'h62 == _match_key_qbytes_5_T_2 ? phv_data_98 : _GEN_10350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10352 = 8'h63 == _match_key_qbytes_5_T_2 ? phv_data_99 : _GEN_10351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10353 = 8'h64 == _match_key_qbytes_5_T_2 ? phv_data_100 : _GEN_10352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10354 = 8'h65 == _match_key_qbytes_5_T_2 ? phv_data_101 : _GEN_10353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10355 = 8'h66 == _match_key_qbytes_5_T_2 ? phv_data_102 : _GEN_10354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10356 = 8'h67 == _match_key_qbytes_5_T_2 ? phv_data_103 : _GEN_10355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10357 = 8'h68 == _match_key_qbytes_5_T_2 ? phv_data_104 : _GEN_10356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10358 = 8'h69 == _match_key_qbytes_5_T_2 ? phv_data_105 : _GEN_10357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10359 = 8'h6a == _match_key_qbytes_5_T_2 ? phv_data_106 : _GEN_10358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10360 = 8'h6b == _match_key_qbytes_5_T_2 ? phv_data_107 : _GEN_10359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10361 = 8'h6c == _match_key_qbytes_5_T_2 ? phv_data_108 : _GEN_10360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10362 = 8'h6d == _match_key_qbytes_5_T_2 ? phv_data_109 : _GEN_10361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10363 = 8'h6e == _match_key_qbytes_5_T_2 ? phv_data_110 : _GEN_10362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10364 = 8'h6f == _match_key_qbytes_5_T_2 ? phv_data_111 : _GEN_10363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10365 = 8'h70 == _match_key_qbytes_5_T_2 ? phv_data_112 : _GEN_10364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10366 = 8'h71 == _match_key_qbytes_5_T_2 ? phv_data_113 : _GEN_10365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10367 = 8'h72 == _match_key_qbytes_5_T_2 ? phv_data_114 : _GEN_10366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10368 = 8'h73 == _match_key_qbytes_5_T_2 ? phv_data_115 : _GEN_10367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10369 = 8'h74 == _match_key_qbytes_5_T_2 ? phv_data_116 : _GEN_10368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10370 = 8'h75 == _match_key_qbytes_5_T_2 ? phv_data_117 : _GEN_10369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10371 = 8'h76 == _match_key_qbytes_5_T_2 ? phv_data_118 : _GEN_10370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10372 = 8'h77 == _match_key_qbytes_5_T_2 ? phv_data_119 : _GEN_10371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10373 = 8'h78 == _match_key_qbytes_5_T_2 ? phv_data_120 : _GEN_10372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10374 = 8'h79 == _match_key_qbytes_5_T_2 ? phv_data_121 : _GEN_10373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10375 = 8'h7a == _match_key_qbytes_5_T_2 ? phv_data_122 : _GEN_10374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10376 = 8'h7b == _match_key_qbytes_5_T_2 ? phv_data_123 : _GEN_10375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10377 = 8'h7c == _match_key_qbytes_5_T_2 ? phv_data_124 : _GEN_10376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10378 = 8'h7d == _match_key_qbytes_5_T_2 ? phv_data_125 : _GEN_10377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10379 = 8'h7e == _match_key_qbytes_5_T_2 ? phv_data_126 : _GEN_10378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10380 = 8'h7f == _match_key_qbytes_5_T_2 ? phv_data_127 : _GEN_10379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10381 = 8'h80 == _match_key_qbytes_5_T_2 ? phv_data_128 : _GEN_10380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10382 = 8'h81 == _match_key_qbytes_5_T_2 ? phv_data_129 : _GEN_10381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10383 = 8'h82 == _match_key_qbytes_5_T_2 ? phv_data_130 : _GEN_10382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10384 = 8'h83 == _match_key_qbytes_5_T_2 ? phv_data_131 : _GEN_10383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10385 = 8'h84 == _match_key_qbytes_5_T_2 ? phv_data_132 : _GEN_10384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10386 = 8'h85 == _match_key_qbytes_5_T_2 ? phv_data_133 : _GEN_10385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10387 = 8'h86 == _match_key_qbytes_5_T_2 ? phv_data_134 : _GEN_10386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10388 = 8'h87 == _match_key_qbytes_5_T_2 ? phv_data_135 : _GEN_10387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10389 = 8'h88 == _match_key_qbytes_5_T_2 ? phv_data_136 : _GEN_10388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10390 = 8'h89 == _match_key_qbytes_5_T_2 ? phv_data_137 : _GEN_10389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10391 = 8'h8a == _match_key_qbytes_5_T_2 ? phv_data_138 : _GEN_10390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10392 = 8'h8b == _match_key_qbytes_5_T_2 ? phv_data_139 : _GEN_10391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10393 = 8'h8c == _match_key_qbytes_5_T_2 ? phv_data_140 : _GEN_10392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10394 = 8'h8d == _match_key_qbytes_5_T_2 ? phv_data_141 : _GEN_10393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10395 = 8'h8e == _match_key_qbytes_5_T_2 ? phv_data_142 : _GEN_10394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10396 = 8'h8f == _match_key_qbytes_5_T_2 ? phv_data_143 : _GEN_10395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10397 = 8'h90 == _match_key_qbytes_5_T_2 ? phv_data_144 : _GEN_10396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10398 = 8'h91 == _match_key_qbytes_5_T_2 ? phv_data_145 : _GEN_10397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10399 = 8'h92 == _match_key_qbytes_5_T_2 ? phv_data_146 : _GEN_10398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10400 = 8'h93 == _match_key_qbytes_5_T_2 ? phv_data_147 : _GEN_10399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10401 = 8'h94 == _match_key_qbytes_5_T_2 ? phv_data_148 : _GEN_10400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10402 = 8'h95 == _match_key_qbytes_5_T_2 ? phv_data_149 : _GEN_10401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10403 = 8'h96 == _match_key_qbytes_5_T_2 ? phv_data_150 : _GEN_10402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10404 = 8'h97 == _match_key_qbytes_5_T_2 ? phv_data_151 : _GEN_10403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10405 = 8'h98 == _match_key_qbytes_5_T_2 ? phv_data_152 : _GEN_10404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10406 = 8'h99 == _match_key_qbytes_5_T_2 ? phv_data_153 : _GEN_10405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10407 = 8'h9a == _match_key_qbytes_5_T_2 ? phv_data_154 : _GEN_10406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10408 = 8'h9b == _match_key_qbytes_5_T_2 ? phv_data_155 : _GEN_10407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10409 = 8'h9c == _match_key_qbytes_5_T_2 ? phv_data_156 : _GEN_10408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10410 = 8'h9d == _match_key_qbytes_5_T_2 ? phv_data_157 : _GEN_10409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10411 = 8'h9e == _match_key_qbytes_5_T_2 ? phv_data_158 : _GEN_10410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10412 = 8'h9f == _match_key_qbytes_5_T_2 ? phv_data_159 : _GEN_10411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10413 = 8'ha0 == _match_key_qbytes_5_T_2 ? phv_data_160 : _GEN_10412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10414 = 8'ha1 == _match_key_qbytes_5_T_2 ? phv_data_161 : _GEN_10413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10415 = 8'ha2 == _match_key_qbytes_5_T_2 ? phv_data_162 : _GEN_10414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10416 = 8'ha3 == _match_key_qbytes_5_T_2 ? phv_data_163 : _GEN_10415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10417 = 8'ha4 == _match_key_qbytes_5_T_2 ? phv_data_164 : _GEN_10416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10418 = 8'ha5 == _match_key_qbytes_5_T_2 ? phv_data_165 : _GEN_10417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10419 = 8'ha6 == _match_key_qbytes_5_T_2 ? phv_data_166 : _GEN_10418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10420 = 8'ha7 == _match_key_qbytes_5_T_2 ? phv_data_167 : _GEN_10419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10421 = 8'ha8 == _match_key_qbytes_5_T_2 ? phv_data_168 : _GEN_10420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10422 = 8'ha9 == _match_key_qbytes_5_T_2 ? phv_data_169 : _GEN_10421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10423 = 8'haa == _match_key_qbytes_5_T_2 ? phv_data_170 : _GEN_10422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10424 = 8'hab == _match_key_qbytes_5_T_2 ? phv_data_171 : _GEN_10423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10425 = 8'hac == _match_key_qbytes_5_T_2 ? phv_data_172 : _GEN_10424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10426 = 8'had == _match_key_qbytes_5_T_2 ? phv_data_173 : _GEN_10425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10427 = 8'hae == _match_key_qbytes_5_T_2 ? phv_data_174 : _GEN_10426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10428 = 8'haf == _match_key_qbytes_5_T_2 ? phv_data_175 : _GEN_10427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10429 = 8'hb0 == _match_key_qbytes_5_T_2 ? phv_data_176 : _GEN_10428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10430 = 8'hb1 == _match_key_qbytes_5_T_2 ? phv_data_177 : _GEN_10429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10431 = 8'hb2 == _match_key_qbytes_5_T_2 ? phv_data_178 : _GEN_10430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10432 = 8'hb3 == _match_key_qbytes_5_T_2 ? phv_data_179 : _GEN_10431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10433 = 8'hb4 == _match_key_qbytes_5_T_2 ? phv_data_180 : _GEN_10432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10434 = 8'hb5 == _match_key_qbytes_5_T_2 ? phv_data_181 : _GEN_10433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10435 = 8'hb6 == _match_key_qbytes_5_T_2 ? phv_data_182 : _GEN_10434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10436 = 8'hb7 == _match_key_qbytes_5_T_2 ? phv_data_183 : _GEN_10435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10437 = 8'hb8 == _match_key_qbytes_5_T_2 ? phv_data_184 : _GEN_10436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10438 = 8'hb9 == _match_key_qbytes_5_T_2 ? phv_data_185 : _GEN_10437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10439 = 8'hba == _match_key_qbytes_5_T_2 ? phv_data_186 : _GEN_10438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10440 = 8'hbb == _match_key_qbytes_5_T_2 ? phv_data_187 : _GEN_10439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10441 = 8'hbc == _match_key_qbytes_5_T_2 ? phv_data_188 : _GEN_10440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10442 = 8'hbd == _match_key_qbytes_5_T_2 ? phv_data_189 : _GEN_10441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10443 = 8'hbe == _match_key_qbytes_5_T_2 ? phv_data_190 : _GEN_10442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10444 = 8'hbf == _match_key_qbytes_5_T_2 ? phv_data_191 : _GEN_10443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10445 = 8'hc0 == _match_key_qbytes_5_T_2 ? phv_data_192 : _GEN_10444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10446 = 8'hc1 == _match_key_qbytes_5_T_2 ? phv_data_193 : _GEN_10445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10447 = 8'hc2 == _match_key_qbytes_5_T_2 ? phv_data_194 : _GEN_10446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10448 = 8'hc3 == _match_key_qbytes_5_T_2 ? phv_data_195 : _GEN_10447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10449 = 8'hc4 == _match_key_qbytes_5_T_2 ? phv_data_196 : _GEN_10448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10450 = 8'hc5 == _match_key_qbytes_5_T_2 ? phv_data_197 : _GEN_10449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10451 = 8'hc6 == _match_key_qbytes_5_T_2 ? phv_data_198 : _GEN_10450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10452 = 8'hc7 == _match_key_qbytes_5_T_2 ? phv_data_199 : _GEN_10451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10453 = 8'hc8 == _match_key_qbytes_5_T_2 ? phv_data_200 : _GEN_10452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10454 = 8'hc9 == _match_key_qbytes_5_T_2 ? phv_data_201 : _GEN_10453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10455 = 8'hca == _match_key_qbytes_5_T_2 ? phv_data_202 : _GEN_10454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10456 = 8'hcb == _match_key_qbytes_5_T_2 ? phv_data_203 : _GEN_10455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10457 = 8'hcc == _match_key_qbytes_5_T_2 ? phv_data_204 : _GEN_10456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10458 = 8'hcd == _match_key_qbytes_5_T_2 ? phv_data_205 : _GEN_10457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10459 = 8'hce == _match_key_qbytes_5_T_2 ? phv_data_206 : _GEN_10458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10460 = 8'hcf == _match_key_qbytes_5_T_2 ? phv_data_207 : _GEN_10459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10461 = 8'hd0 == _match_key_qbytes_5_T_2 ? phv_data_208 : _GEN_10460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10462 = 8'hd1 == _match_key_qbytes_5_T_2 ? phv_data_209 : _GEN_10461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10463 = 8'hd2 == _match_key_qbytes_5_T_2 ? phv_data_210 : _GEN_10462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10464 = 8'hd3 == _match_key_qbytes_5_T_2 ? phv_data_211 : _GEN_10463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10465 = 8'hd4 == _match_key_qbytes_5_T_2 ? phv_data_212 : _GEN_10464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10466 = 8'hd5 == _match_key_qbytes_5_T_2 ? phv_data_213 : _GEN_10465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10467 = 8'hd6 == _match_key_qbytes_5_T_2 ? phv_data_214 : _GEN_10466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10468 = 8'hd7 == _match_key_qbytes_5_T_2 ? phv_data_215 : _GEN_10467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10469 = 8'hd8 == _match_key_qbytes_5_T_2 ? phv_data_216 : _GEN_10468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10470 = 8'hd9 == _match_key_qbytes_5_T_2 ? phv_data_217 : _GEN_10469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10471 = 8'hda == _match_key_qbytes_5_T_2 ? phv_data_218 : _GEN_10470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10472 = 8'hdb == _match_key_qbytes_5_T_2 ? phv_data_219 : _GEN_10471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10473 = 8'hdc == _match_key_qbytes_5_T_2 ? phv_data_220 : _GEN_10472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10474 = 8'hdd == _match_key_qbytes_5_T_2 ? phv_data_221 : _GEN_10473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10475 = 8'hde == _match_key_qbytes_5_T_2 ? phv_data_222 : _GEN_10474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10476 = 8'hdf == _match_key_qbytes_5_T_2 ? phv_data_223 : _GEN_10475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10477 = 8'he0 == _match_key_qbytes_5_T_2 ? phv_data_224 : _GEN_10476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10478 = 8'he1 == _match_key_qbytes_5_T_2 ? phv_data_225 : _GEN_10477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10479 = 8'he2 == _match_key_qbytes_5_T_2 ? phv_data_226 : _GEN_10478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10480 = 8'he3 == _match_key_qbytes_5_T_2 ? phv_data_227 : _GEN_10479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10481 = 8'he4 == _match_key_qbytes_5_T_2 ? phv_data_228 : _GEN_10480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10482 = 8'he5 == _match_key_qbytes_5_T_2 ? phv_data_229 : _GEN_10481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10483 = 8'he6 == _match_key_qbytes_5_T_2 ? phv_data_230 : _GEN_10482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10484 = 8'he7 == _match_key_qbytes_5_T_2 ? phv_data_231 : _GEN_10483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10485 = 8'he8 == _match_key_qbytes_5_T_2 ? phv_data_232 : _GEN_10484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10486 = 8'he9 == _match_key_qbytes_5_T_2 ? phv_data_233 : _GEN_10485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10487 = 8'hea == _match_key_qbytes_5_T_2 ? phv_data_234 : _GEN_10486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10488 = 8'heb == _match_key_qbytes_5_T_2 ? phv_data_235 : _GEN_10487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10489 = 8'hec == _match_key_qbytes_5_T_2 ? phv_data_236 : _GEN_10488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10490 = 8'hed == _match_key_qbytes_5_T_2 ? phv_data_237 : _GEN_10489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10491 = 8'hee == _match_key_qbytes_5_T_2 ? phv_data_238 : _GEN_10490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10492 = 8'hef == _match_key_qbytes_5_T_2 ? phv_data_239 : _GEN_10491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10493 = 8'hf0 == _match_key_qbytes_5_T_2 ? phv_data_240 : _GEN_10492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10494 = 8'hf1 == _match_key_qbytes_5_T_2 ? phv_data_241 : _GEN_10493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10495 = 8'hf2 == _match_key_qbytes_5_T_2 ? phv_data_242 : _GEN_10494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10496 = 8'hf3 == _match_key_qbytes_5_T_2 ? phv_data_243 : _GEN_10495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10497 = 8'hf4 == _match_key_qbytes_5_T_2 ? phv_data_244 : _GEN_10496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10498 = 8'hf5 == _match_key_qbytes_5_T_2 ? phv_data_245 : _GEN_10497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10499 = 8'hf6 == _match_key_qbytes_5_T_2 ? phv_data_246 : _GEN_10498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10500 = 8'hf7 == _match_key_qbytes_5_T_2 ? phv_data_247 : _GEN_10499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10501 = 8'hf8 == _match_key_qbytes_5_T_2 ? phv_data_248 : _GEN_10500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10502 = 8'hf9 == _match_key_qbytes_5_T_2 ? phv_data_249 : _GEN_10501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10503 = 8'hfa == _match_key_qbytes_5_T_2 ? phv_data_250 : _GEN_10502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10504 = 8'hfb == _match_key_qbytes_5_T_2 ? phv_data_251 : _GEN_10503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10505 = 8'hfc == _match_key_qbytes_5_T_2 ? phv_data_252 : _GEN_10504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10506 = 8'hfd == _match_key_qbytes_5_T_2 ? phv_data_253 : _GEN_10505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10507 = 8'hfe == _match_key_qbytes_5_T_2 ? phv_data_254 : _GEN_10506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10508 = 8'hff == _match_key_qbytes_5_T_2 ? phv_data_255 : _GEN_10507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_17446 = {{1'd0}, _match_key_qbytes_5_T_2}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10509 = 9'h100 == _GEN_17446 ? phv_data_256 : _GEN_10508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10510 = 9'h101 == _GEN_17446 ? phv_data_257 : _GEN_10509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10511 = 9'h102 == _GEN_17446 ? phv_data_258 : _GEN_10510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10512 = 9'h103 == _GEN_17446 ? phv_data_259 : _GEN_10511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10513 = 9'h104 == _GEN_17446 ? phv_data_260 : _GEN_10512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10514 = 9'h105 == _GEN_17446 ? phv_data_261 : _GEN_10513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10515 = 9'h106 == _GEN_17446 ? phv_data_262 : _GEN_10514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10516 = 9'h107 == _GEN_17446 ? phv_data_263 : _GEN_10515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10517 = 9'h108 == _GEN_17446 ? phv_data_264 : _GEN_10516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10518 = 9'h109 == _GEN_17446 ? phv_data_265 : _GEN_10517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10519 = 9'h10a == _GEN_17446 ? phv_data_266 : _GEN_10518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10520 = 9'h10b == _GEN_17446 ? phv_data_267 : _GEN_10519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10521 = 9'h10c == _GEN_17446 ? phv_data_268 : _GEN_10520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10522 = 9'h10d == _GEN_17446 ? phv_data_269 : _GEN_10521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10523 = 9'h10e == _GEN_17446 ? phv_data_270 : _GEN_10522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10524 = 9'h10f == _GEN_17446 ? phv_data_271 : _GEN_10523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10525 = 9'h110 == _GEN_17446 ? phv_data_272 : _GEN_10524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10526 = 9'h111 == _GEN_17446 ? phv_data_273 : _GEN_10525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10527 = 9'h112 == _GEN_17446 ? phv_data_274 : _GEN_10526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10528 = 9'h113 == _GEN_17446 ? phv_data_275 : _GEN_10527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10529 = 9'h114 == _GEN_17446 ? phv_data_276 : _GEN_10528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10530 = 9'h115 == _GEN_17446 ? phv_data_277 : _GEN_10529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10531 = 9'h116 == _GEN_17446 ? phv_data_278 : _GEN_10530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10532 = 9'h117 == _GEN_17446 ? phv_data_279 : _GEN_10531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10533 = 9'h118 == _GEN_17446 ? phv_data_280 : _GEN_10532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10534 = 9'h119 == _GEN_17446 ? phv_data_281 : _GEN_10533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10535 = 9'h11a == _GEN_17446 ? phv_data_282 : _GEN_10534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10536 = 9'h11b == _GEN_17446 ? phv_data_283 : _GEN_10535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10537 = 9'h11c == _GEN_17446 ? phv_data_284 : _GEN_10536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10538 = 9'h11d == _GEN_17446 ? phv_data_285 : _GEN_10537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10539 = 9'h11e == _GEN_17446 ? phv_data_286 : _GEN_10538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10540 = 9'h11f == _GEN_17446 ? phv_data_287 : _GEN_10539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10541 = 9'h120 == _GEN_17446 ? phv_data_288 : _GEN_10540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10542 = 9'h121 == _GEN_17446 ? phv_data_289 : _GEN_10541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10543 = 9'h122 == _GEN_17446 ? phv_data_290 : _GEN_10542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10544 = 9'h123 == _GEN_17446 ? phv_data_291 : _GEN_10543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10545 = 9'h124 == _GEN_17446 ? phv_data_292 : _GEN_10544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10546 = 9'h125 == _GEN_17446 ? phv_data_293 : _GEN_10545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10547 = 9'h126 == _GEN_17446 ? phv_data_294 : _GEN_10546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10548 = 9'h127 == _GEN_17446 ? phv_data_295 : _GEN_10547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10549 = 9'h128 == _GEN_17446 ? phv_data_296 : _GEN_10548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10550 = 9'h129 == _GEN_17446 ? phv_data_297 : _GEN_10549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10551 = 9'h12a == _GEN_17446 ? phv_data_298 : _GEN_10550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10552 = 9'h12b == _GEN_17446 ? phv_data_299 : _GEN_10551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10553 = 9'h12c == _GEN_17446 ? phv_data_300 : _GEN_10552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10554 = 9'h12d == _GEN_17446 ? phv_data_301 : _GEN_10553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10555 = 9'h12e == _GEN_17446 ? phv_data_302 : _GEN_10554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10556 = 9'h12f == _GEN_17446 ? phv_data_303 : _GEN_10555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10557 = 9'h130 == _GEN_17446 ? phv_data_304 : _GEN_10556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10558 = 9'h131 == _GEN_17446 ? phv_data_305 : _GEN_10557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10559 = 9'h132 == _GEN_17446 ? phv_data_306 : _GEN_10558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10560 = 9'h133 == _GEN_17446 ? phv_data_307 : _GEN_10559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10561 = 9'h134 == _GEN_17446 ? phv_data_308 : _GEN_10560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10562 = 9'h135 == _GEN_17446 ? phv_data_309 : _GEN_10561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10563 = 9'h136 == _GEN_17446 ? phv_data_310 : _GEN_10562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10564 = 9'h137 == _GEN_17446 ? phv_data_311 : _GEN_10563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10565 = 9'h138 == _GEN_17446 ? phv_data_312 : _GEN_10564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10566 = 9'h139 == _GEN_17446 ? phv_data_313 : _GEN_10565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10567 = 9'h13a == _GEN_17446 ? phv_data_314 : _GEN_10566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10568 = 9'h13b == _GEN_17446 ? phv_data_315 : _GEN_10567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10569 = 9'h13c == _GEN_17446 ? phv_data_316 : _GEN_10568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10570 = 9'h13d == _GEN_17446 ? phv_data_317 : _GEN_10569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10571 = 9'h13e == _GEN_17446 ? phv_data_318 : _GEN_10570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10572 = 9'h13f == _GEN_17446 ? phv_data_319 : _GEN_10571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10573 = 9'h140 == _GEN_17446 ? phv_data_320 : _GEN_10572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10574 = 9'h141 == _GEN_17446 ? phv_data_321 : _GEN_10573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10575 = 9'h142 == _GEN_17446 ? phv_data_322 : _GEN_10574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10576 = 9'h143 == _GEN_17446 ? phv_data_323 : _GEN_10575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10577 = 9'h144 == _GEN_17446 ? phv_data_324 : _GEN_10576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10578 = 9'h145 == _GEN_17446 ? phv_data_325 : _GEN_10577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10579 = 9'h146 == _GEN_17446 ? phv_data_326 : _GEN_10578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10580 = 9'h147 == _GEN_17446 ? phv_data_327 : _GEN_10579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10581 = 9'h148 == _GEN_17446 ? phv_data_328 : _GEN_10580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10582 = 9'h149 == _GEN_17446 ? phv_data_329 : _GEN_10581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10583 = 9'h14a == _GEN_17446 ? phv_data_330 : _GEN_10582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10584 = 9'h14b == _GEN_17446 ? phv_data_331 : _GEN_10583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10585 = 9'h14c == _GEN_17446 ? phv_data_332 : _GEN_10584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10586 = 9'h14d == _GEN_17446 ? phv_data_333 : _GEN_10585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10587 = 9'h14e == _GEN_17446 ? phv_data_334 : _GEN_10586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10588 = 9'h14f == _GEN_17446 ? phv_data_335 : _GEN_10587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10589 = 9'h150 == _GEN_17446 ? phv_data_336 : _GEN_10588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10590 = 9'h151 == _GEN_17446 ? phv_data_337 : _GEN_10589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10591 = 9'h152 == _GEN_17446 ? phv_data_338 : _GEN_10590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10592 = 9'h153 == _GEN_17446 ? phv_data_339 : _GEN_10591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10593 = 9'h154 == _GEN_17446 ? phv_data_340 : _GEN_10592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10594 = 9'h155 == _GEN_17446 ? phv_data_341 : _GEN_10593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10595 = 9'h156 == _GEN_17446 ? phv_data_342 : _GEN_10594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10596 = 9'h157 == _GEN_17446 ? phv_data_343 : _GEN_10595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10597 = 9'h158 == _GEN_17446 ? phv_data_344 : _GEN_10596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10598 = 9'h159 == _GEN_17446 ? phv_data_345 : _GEN_10597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10599 = 9'h15a == _GEN_17446 ? phv_data_346 : _GEN_10598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10600 = 9'h15b == _GEN_17446 ? phv_data_347 : _GEN_10599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10601 = 9'h15c == _GEN_17446 ? phv_data_348 : _GEN_10600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10602 = 9'h15d == _GEN_17446 ? phv_data_349 : _GEN_10601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10603 = 9'h15e == _GEN_17446 ? phv_data_350 : _GEN_10602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10604 = 9'h15f == _GEN_17446 ? phv_data_351 : _GEN_10603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10605 = 9'h160 == _GEN_17446 ? phv_data_352 : _GEN_10604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10606 = 9'h161 == _GEN_17446 ? phv_data_353 : _GEN_10605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10607 = 9'h162 == _GEN_17446 ? phv_data_354 : _GEN_10606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10608 = 9'h163 == _GEN_17446 ? phv_data_355 : _GEN_10607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10609 = 9'h164 == _GEN_17446 ? phv_data_356 : _GEN_10608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10610 = 9'h165 == _GEN_17446 ? phv_data_357 : _GEN_10609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10611 = 9'h166 == _GEN_17446 ? phv_data_358 : _GEN_10610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10612 = 9'h167 == _GEN_17446 ? phv_data_359 : _GEN_10611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10613 = 9'h168 == _GEN_17446 ? phv_data_360 : _GEN_10612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10614 = 9'h169 == _GEN_17446 ? phv_data_361 : _GEN_10613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10615 = 9'h16a == _GEN_17446 ? phv_data_362 : _GEN_10614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10616 = 9'h16b == _GEN_17446 ? phv_data_363 : _GEN_10615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10617 = 9'h16c == _GEN_17446 ? phv_data_364 : _GEN_10616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10618 = 9'h16d == _GEN_17446 ? phv_data_365 : _GEN_10617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10619 = 9'h16e == _GEN_17446 ? phv_data_366 : _GEN_10618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10620 = 9'h16f == _GEN_17446 ? phv_data_367 : _GEN_10619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10621 = 9'h170 == _GEN_17446 ? phv_data_368 : _GEN_10620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10622 = 9'h171 == _GEN_17446 ? phv_data_369 : _GEN_10621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10623 = 9'h172 == _GEN_17446 ? phv_data_370 : _GEN_10622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10624 = 9'h173 == _GEN_17446 ? phv_data_371 : _GEN_10623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10625 = 9'h174 == _GEN_17446 ? phv_data_372 : _GEN_10624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10626 = 9'h175 == _GEN_17446 ? phv_data_373 : _GEN_10625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10627 = 9'h176 == _GEN_17446 ? phv_data_374 : _GEN_10626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10628 = 9'h177 == _GEN_17446 ? phv_data_375 : _GEN_10627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10629 = 9'h178 == _GEN_17446 ? phv_data_376 : _GEN_10628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10630 = 9'h179 == _GEN_17446 ? phv_data_377 : _GEN_10629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10631 = 9'h17a == _GEN_17446 ? phv_data_378 : _GEN_10630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10632 = 9'h17b == _GEN_17446 ? phv_data_379 : _GEN_10631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10633 = 9'h17c == _GEN_17446 ? phv_data_380 : _GEN_10632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10634 = 9'h17d == _GEN_17446 ? phv_data_381 : _GEN_10633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10635 = 9'h17e == _GEN_17446 ? phv_data_382 : _GEN_10634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10636 = 9'h17f == _GEN_17446 ? phv_data_383 : _GEN_10635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10637 = 9'h180 == _GEN_17446 ? phv_data_384 : _GEN_10636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10638 = 9'h181 == _GEN_17446 ? phv_data_385 : _GEN_10637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10639 = 9'h182 == _GEN_17446 ? phv_data_386 : _GEN_10638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10640 = 9'h183 == _GEN_17446 ? phv_data_387 : _GEN_10639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10641 = 9'h184 == _GEN_17446 ? phv_data_388 : _GEN_10640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10642 = 9'h185 == _GEN_17446 ? phv_data_389 : _GEN_10641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10643 = 9'h186 == _GEN_17446 ? phv_data_390 : _GEN_10642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10644 = 9'h187 == _GEN_17446 ? phv_data_391 : _GEN_10643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10645 = 9'h188 == _GEN_17446 ? phv_data_392 : _GEN_10644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10646 = 9'h189 == _GEN_17446 ? phv_data_393 : _GEN_10645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10647 = 9'h18a == _GEN_17446 ? phv_data_394 : _GEN_10646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10648 = 9'h18b == _GEN_17446 ? phv_data_395 : _GEN_10647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10649 = 9'h18c == _GEN_17446 ? phv_data_396 : _GEN_10648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10650 = 9'h18d == _GEN_17446 ? phv_data_397 : _GEN_10649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10651 = 9'h18e == _GEN_17446 ? phv_data_398 : _GEN_10650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10652 = 9'h18f == _GEN_17446 ? phv_data_399 : _GEN_10651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10653 = 9'h190 == _GEN_17446 ? phv_data_400 : _GEN_10652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10654 = 9'h191 == _GEN_17446 ? phv_data_401 : _GEN_10653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10655 = 9'h192 == _GEN_17446 ? phv_data_402 : _GEN_10654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10656 = 9'h193 == _GEN_17446 ? phv_data_403 : _GEN_10655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10657 = 9'h194 == _GEN_17446 ? phv_data_404 : _GEN_10656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10658 = 9'h195 == _GEN_17446 ? phv_data_405 : _GEN_10657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10659 = 9'h196 == _GEN_17446 ? phv_data_406 : _GEN_10658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10660 = 9'h197 == _GEN_17446 ? phv_data_407 : _GEN_10659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10661 = 9'h198 == _GEN_17446 ? phv_data_408 : _GEN_10660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10662 = 9'h199 == _GEN_17446 ? phv_data_409 : _GEN_10661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10663 = 9'h19a == _GEN_17446 ? phv_data_410 : _GEN_10662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10664 = 9'h19b == _GEN_17446 ? phv_data_411 : _GEN_10663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10665 = 9'h19c == _GEN_17446 ? phv_data_412 : _GEN_10664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10666 = 9'h19d == _GEN_17446 ? phv_data_413 : _GEN_10665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10667 = 9'h19e == _GEN_17446 ? phv_data_414 : _GEN_10666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10668 = 9'h19f == _GEN_17446 ? phv_data_415 : _GEN_10667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10669 = 9'h1a0 == _GEN_17446 ? phv_data_416 : _GEN_10668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10670 = 9'h1a1 == _GEN_17446 ? phv_data_417 : _GEN_10669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10671 = 9'h1a2 == _GEN_17446 ? phv_data_418 : _GEN_10670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10672 = 9'h1a3 == _GEN_17446 ? phv_data_419 : _GEN_10671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10673 = 9'h1a4 == _GEN_17446 ? phv_data_420 : _GEN_10672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10674 = 9'h1a5 == _GEN_17446 ? phv_data_421 : _GEN_10673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10675 = 9'h1a6 == _GEN_17446 ? phv_data_422 : _GEN_10674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10676 = 9'h1a7 == _GEN_17446 ? phv_data_423 : _GEN_10675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10677 = 9'h1a8 == _GEN_17446 ? phv_data_424 : _GEN_10676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10678 = 9'h1a9 == _GEN_17446 ? phv_data_425 : _GEN_10677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10679 = 9'h1aa == _GEN_17446 ? phv_data_426 : _GEN_10678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10680 = 9'h1ab == _GEN_17446 ? phv_data_427 : _GEN_10679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10681 = 9'h1ac == _GEN_17446 ? phv_data_428 : _GEN_10680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10682 = 9'h1ad == _GEN_17446 ? phv_data_429 : _GEN_10681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10683 = 9'h1ae == _GEN_17446 ? phv_data_430 : _GEN_10682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10684 = 9'h1af == _GEN_17446 ? phv_data_431 : _GEN_10683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10685 = 9'h1b0 == _GEN_17446 ? phv_data_432 : _GEN_10684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10686 = 9'h1b1 == _GEN_17446 ? phv_data_433 : _GEN_10685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10687 = 9'h1b2 == _GEN_17446 ? phv_data_434 : _GEN_10686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10688 = 9'h1b3 == _GEN_17446 ? phv_data_435 : _GEN_10687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10689 = 9'h1b4 == _GEN_17446 ? phv_data_436 : _GEN_10688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10690 = 9'h1b5 == _GEN_17446 ? phv_data_437 : _GEN_10689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10691 = 9'h1b6 == _GEN_17446 ? phv_data_438 : _GEN_10690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10692 = 9'h1b7 == _GEN_17446 ? phv_data_439 : _GEN_10691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10693 = 9'h1b8 == _GEN_17446 ? phv_data_440 : _GEN_10692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10694 = 9'h1b9 == _GEN_17446 ? phv_data_441 : _GEN_10693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10695 = 9'h1ba == _GEN_17446 ? phv_data_442 : _GEN_10694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10696 = 9'h1bb == _GEN_17446 ? phv_data_443 : _GEN_10695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10697 = 9'h1bc == _GEN_17446 ? phv_data_444 : _GEN_10696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10698 = 9'h1bd == _GEN_17446 ? phv_data_445 : _GEN_10697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10699 = 9'h1be == _GEN_17446 ? phv_data_446 : _GEN_10698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10700 = 9'h1bf == _GEN_17446 ? phv_data_447 : _GEN_10699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10701 = 9'h1c0 == _GEN_17446 ? phv_data_448 : _GEN_10700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10702 = 9'h1c1 == _GEN_17446 ? phv_data_449 : _GEN_10701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10703 = 9'h1c2 == _GEN_17446 ? phv_data_450 : _GEN_10702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10704 = 9'h1c3 == _GEN_17446 ? phv_data_451 : _GEN_10703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10705 = 9'h1c4 == _GEN_17446 ? phv_data_452 : _GEN_10704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10706 = 9'h1c5 == _GEN_17446 ? phv_data_453 : _GEN_10705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10707 = 9'h1c6 == _GEN_17446 ? phv_data_454 : _GEN_10706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10708 = 9'h1c7 == _GEN_17446 ? phv_data_455 : _GEN_10707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10709 = 9'h1c8 == _GEN_17446 ? phv_data_456 : _GEN_10708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10710 = 9'h1c9 == _GEN_17446 ? phv_data_457 : _GEN_10709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10711 = 9'h1ca == _GEN_17446 ? phv_data_458 : _GEN_10710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10712 = 9'h1cb == _GEN_17446 ? phv_data_459 : _GEN_10711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10713 = 9'h1cc == _GEN_17446 ? phv_data_460 : _GEN_10712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10714 = 9'h1cd == _GEN_17446 ? phv_data_461 : _GEN_10713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10715 = 9'h1ce == _GEN_17446 ? phv_data_462 : _GEN_10714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10716 = 9'h1cf == _GEN_17446 ? phv_data_463 : _GEN_10715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10717 = 9'h1d0 == _GEN_17446 ? phv_data_464 : _GEN_10716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10718 = 9'h1d1 == _GEN_17446 ? phv_data_465 : _GEN_10717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10719 = 9'h1d2 == _GEN_17446 ? phv_data_466 : _GEN_10718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10720 = 9'h1d3 == _GEN_17446 ? phv_data_467 : _GEN_10719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10721 = 9'h1d4 == _GEN_17446 ? phv_data_468 : _GEN_10720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10722 = 9'h1d5 == _GEN_17446 ? phv_data_469 : _GEN_10721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10723 = 9'h1d6 == _GEN_17446 ? phv_data_470 : _GEN_10722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10724 = 9'h1d7 == _GEN_17446 ? phv_data_471 : _GEN_10723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10725 = 9'h1d8 == _GEN_17446 ? phv_data_472 : _GEN_10724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10726 = 9'h1d9 == _GEN_17446 ? phv_data_473 : _GEN_10725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10727 = 9'h1da == _GEN_17446 ? phv_data_474 : _GEN_10726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10728 = 9'h1db == _GEN_17446 ? phv_data_475 : _GEN_10727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10729 = 9'h1dc == _GEN_17446 ? phv_data_476 : _GEN_10728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10730 = 9'h1dd == _GEN_17446 ? phv_data_477 : _GEN_10729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10731 = 9'h1de == _GEN_17446 ? phv_data_478 : _GEN_10730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10732 = 9'h1df == _GEN_17446 ? phv_data_479 : _GEN_10731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10733 = 9'h1e0 == _GEN_17446 ? phv_data_480 : _GEN_10732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10734 = 9'h1e1 == _GEN_17446 ? phv_data_481 : _GEN_10733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10735 = 9'h1e2 == _GEN_17446 ? phv_data_482 : _GEN_10734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10736 = 9'h1e3 == _GEN_17446 ? phv_data_483 : _GEN_10735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10737 = 9'h1e4 == _GEN_17446 ? phv_data_484 : _GEN_10736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10738 = 9'h1e5 == _GEN_17446 ? phv_data_485 : _GEN_10737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10739 = 9'h1e6 == _GEN_17446 ? phv_data_486 : _GEN_10738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10740 = 9'h1e7 == _GEN_17446 ? phv_data_487 : _GEN_10739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10741 = 9'h1e8 == _GEN_17446 ? phv_data_488 : _GEN_10740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10742 = 9'h1e9 == _GEN_17446 ? phv_data_489 : _GEN_10741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10743 = 9'h1ea == _GEN_17446 ? phv_data_490 : _GEN_10742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10744 = 9'h1eb == _GEN_17446 ? phv_data_491 : _GEN_10743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10745 = 9'h1ec == _GEN_17446 ? phv_data_492 : _GEN_10744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10746 = 9'h1ed == _GEN_17446 ? phv_data_493 : _GEN_10745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10747 = 9'h1ee == _GEN_17446 ? phv_data_494 : _GEN_10746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10748 = 9'h1ef == _GEN_17446 ? phv_data_495 : _GEN_10747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10749 = 9'h1f0 == _GEN_17446 ? phv_data_496 : _GEN_10748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10750 = 9'h1f1 == _GEN_17446 ? phv_data_497 : _GEN_10749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10751 = 9'h1f2 == _GEN_17446 ? phv_data_498 : _GEN_10750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10752 = 9'h1f3 == _GEN_17446 ? phv_data_499 : _GEN_10751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10753 = 9'h1f4 == _GEN_17446 ? phv_data_500 : _GEN_10752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10754 = 9'h1f5 == _GEN_17446 ? phv_data_501 : _GEN_10753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10755 = 9'h1f6 == _GEN_17446 ? phv_data_502 : _GEN_10754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10756 = 9'h1f7 == _GEN_17446 ? phv_data_503 : _GEN_10755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10757 = 9'h1f8 == _GEN_17446 ? phv_data_504 : _GEN_10756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10758 = 9'h1f9 == _GEN_17446 ? phv_data_505 : _GEN_10757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10759 = 9'h1fa == _GEN_17446 ? phv_data_506 : _GEN_10758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10760 = 9'h1fb == _GEN_17446 ? phv_data_507 : _GEN_10759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10761 = 9'h1fc == _GEN_17446 ? phv_data_508 : _GEN_10760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10762 = 9'h1fd == _GEN_17446 ? phv_data_509 : _GEN_10761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10763 = 9'h1fe == _GEN_17446 ? phv_data_510 : _GEN_10762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10764 = 9'h1ff == _GEN_17446 ? phv_data_511 : _GEN_10763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10766 = 8'h1 == local_offset_5 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10767 = 8'h2 == local_offset_5 ? phv_data_2 : _GEN_10766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10768 = 8'h3 == local_offset_5 ? phv_data_3 : _GEN_10767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10769 = 8'h4 == local_offset_5 ? phv_data_4 : _GEN_10768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10770 = 8'h5 == local_offset_5 ? phv_data_5 : _GEN_10769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10771 = 8'h6 == local_offset_5 ? phv_data_6 : _GEN_10770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10772 = 8'h7 == local_offset_5 ? phv_data_7 : _GEN_10771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10773 = 8'h8 == local_offset_5 ? phv_data_8 : _GEN_10772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10774 = 8'h9 == local_offset_5 ? phv_data_9 : _GEN_10773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10775 = 8'ha == local_offset_5 ? phv_data_10 : _GEN_10774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10776 = 8'hb == local_offset_5 ? phv_data_11 : _GEN_10775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10777 = 8'hc == local_offset_5 ? phv_data_12 : _GEN_10776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10778 = 8'hd == local_offset_5 ? phv_data_13 : _GEN_10777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10779 = 8'he == local_offset_5 ? phv_data_14 : _GEN_10778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10780 = 8'hf == local_offset_5 ? phv_data_15 : _GEN_10779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10781 = 8'h10 == local_offset_5 ? phv_data_16 : _GEN_10780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10782 = 8'h11 == local_offset_5 ? phv_data_17 : _GEN_10781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10783 = 8'h12 == local_offset_5 ? phv_data_18 : _GEN_10782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10784 = 8'h13 == local_offset_5 ? phv_data_19 : _GEN_10783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10785 = 8'h14 == local_offset_5 ? phv_data_20 : _GEN_10784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10786 = 8'h15 == local_offset_5 ? phv_data_21 : _GEN_10785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10787 = 8'h16 == local_offset_5 ? phv_data_22 : _GEN_10786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10788 = 8'h17 == local_offset_5 ? phv_data_23 : _GEN_10787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10789 = 8'h18 == local_offset_5 ? phv_data_24 : _GEN_10788; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10790 = 8'h19 == local_offset_5 ? phv_data_25 : _GEN_10789; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10791 = 8'h1a == local_offset_5 ? phv_data_26 : _GEN_10790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10792 = 8'h1b == local_offset_5 ? phv_data_27 : _GEN_10791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10793 = 8'h1c == local_offset_5 ? phv_data_28 : _GEN_10792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10794 = 8'h1d == local_offset_5 ? phv_data_29 : _GEN_10793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10795 = 8'h1e == local_offset_5 ? phv_data_30 : _GEN_10794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10796 = 8'h1f == local_offset_5 ? phv_data_31 : _GEN_10795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10797 = 8'h20 == local_offset_5 ? phv_data_32 : _GEN_10796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10798 = 8'h21 == local_offset_5 ? phv_data_33 : _GEN_10797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10799 = 8'h22 == local_offset_5 ? phv_data_34 : _GEN_10798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10800 = 8'h23 == local_offset_5 ? phv_data_35 : _GEN_10799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10801 = 8'h24 == local_offset_5 ? phv_data_36 : _GEN_10800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10802 = 8'h25 == local_offset_5 ? phv_data_37 : _GEN_10801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10803 = 8'h26 == local_offset_5 ? phv_data_38 : _GEN_10802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10804 = 8'h27 == local_offset_5 ? phv_data_39 : _GEN_10803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10805 = 8'h28 == local_offset_5 ? phv_data_40 : _GEN_10804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10806 = 8'h29 == local_offset_5 ? phv_data_41 : _GEN_10805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10807 = 8'h2a == local_offset_5 ? phv_data_42 : _GEN_10806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10808 = 8'h2b == local_offset_5 ? phv_data_43 : _GEN_10807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10809 = 8'h2c == local_offset_5 ? phv_data_44 : _GEN_10808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10810 = 8'h2d == local_offset_5 ? phv_data_45 : _GEN_10809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10811 = 8'h2e == local_offset_5 ? phv_data_46 : _GEN_10810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10812 = 8'h2f == local_offset_5 ? phv_data_47 : _GEN_10811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10813 = 8'h30 == local_offset_5 ? phv_data_48 : _GEN_10812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10814 = 8'h31 == local_offset_5 ? phv_data_49 : _GEN_10813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10815 = 8'h32 == local_offset_5 ? phv_data_50 : _GEN_10814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10816 = 8'h33 == local_offset_5 ? phv_data_51 : _GEN_10815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10817 = 8'h34 == local_offset_5 ? phv_data_52 : _GEN_10816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10818 = 8'h35 == local_offset_5 ? phv_data_53 : _GEN_10817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10819 = 8'h36 == local_offset_5 ? phv_data_54 : _GEN_10818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10820 = 8'h37 == local_offset_5 ? phv_data_55 : _GEN_10819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10821 = 8'h38 == local_offset_5 ? phv_data_56 : _GEN_10820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10822 = 8'h39 == local_offset_5 ? phv_data_57 : _GEN_10821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10823 = 8'h3a == local_offset_5 ? phv_data_58 : _GEN_10822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10824 = 8'h3b == local_offset_5 ? phv_data_59 : _GEN_10823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10825 = 8'h3c == local_offset_5 ? phv_data_60 : _GEN_10824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10826 = 8'h3d == local_offset_5 ? phv_data_61 : _GEN_10825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10827 = 8'h3e == local_offset_5 ? phv_data_62 : _GEN_10826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10828 = 8'h3f == local_offset_5 ? phv_data_63 : _GEN_10827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10829 = 8'h40 == local_offset_5 ? phv_data_64 : _GEN_10828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10830 = 8'h41 == local_offset_5 ? phv_data_65 : _GEN_10829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10831 = 8'h42 == local_offset_5 ? phv_data_66 : _GEN_10830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10832 = 8'h43 == local_offset_5 ? phv_data_67 : _GEN_10831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10833 = 8'h44 == local_offset_5 ? phv_data_68 : _GEN_10832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10834 = 8'h45 == local_offset_5 ? phv_data_69 : _GEN_10833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10835 = 8'h46 == local_offset_5 ? phv_data_70 : _GEN_10834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10836 = 8'h47 == local_offset_5 ? phv_data_71 : _GEN_10835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10837 = 8'h48 == local_offset_5 ? phv_data_72 : _GEN_10836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10838 = 8'h49 == local_offset_5 ? phv_data_73 : _GEN_10837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10839 = 8'h4a == local_offset_5 ? phv_data_74 : _GEN_10838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10840 = 8'h4b == local_offset_5 ? phv_data_75 : _GEN_10839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10841 = 8'h4c == local_offset_5 ? phv_data_76 : _GEN_10840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10842 = 8'h4d == local_offset_5 ? phv_data_77 : _GEN_10841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10843 = 8'h4e == local_offset_5 ? phv_data_78 : _GEN_10842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10844 = 8'h4f == local_offset_5 ? phv_data_79 : _GEN_10843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10845 = 8'h50 == local_offset_5 ? phv_data_80 : _GEN_10844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10846 = 8'h51 == local_offset_5 ? phv_data_81 : _GEN_10845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10847 = 8'h52 == local_offset_5 ? phv_data_82 : _GEN_10846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10848 = 8'h53 == local_offset_5 ? phv_data_83 : _GEN_10847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10849 = 8'h54 == local_offset_5 ? phv_data_84 : _GEN_10848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10850 = 8'h55 == local_offset_5 ? phv_data_85 : _GEN_10849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10851 = 8'h56 == local_offset_5 ? phv_data_86 : _GEN_10850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10852 = 8'h57 == local_offset_5 ? phv_data_87 : _GEN_10851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10853 = 8'h58 == local_offset_5 ? phv_data_88 : _GEN_10852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10854 = 8'h59 == local_offset_5 ? phv_data_89 : _GEN_10853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10855 = 8'h5a == local_offset_5 ? phv_data_90 : _GEN_10854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10856 = 8'h5b == local_offset_5 ? phv_data_91 : _GEN_10855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10857 = 8'h5c == local_offset_5 ? phv_data_92 : _GEN_10856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10858 = 8'h5d == local_offset_5 ? phv_data_93 : _GEN_10857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10859 = 8'h5e == local_offset_5 ? phv_data_94 : _GEN_10858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10860 = 8'h5f == local_offset_5 ? phv_data_95 : _GEN_10859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10861 = 8'h60 == local_offset_5 ? phv_data_96 : _GEN_10860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10862 = 8'h61 == local_offset_5 ? phv_data_97 : _GEN_10861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10863 = 8'h62 == local_offset_5 ? phv_data_98 : _GEN_10862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10864 = 8'h63 == local_offset_5 ? phv_data_99 : _GEN_10863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10865 = 8'h64 == local_offset_5 ? phv_data_100 : _GEN_10864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10866 = 8'h65 == local_offset_5 ? phv_data_101 : _GEN_10865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10867 = 8'h66 == local_offset_5 ? phv_data_102 : _GEN_10866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10868 = 8'h67 == local_offset_5 ? phv_data_103 : _GEN_10867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10869 = 8'h68 == local_offset_5 ? phv_data_104 : _GEN_10868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10870 = 8'h69 == local_offset_5 ? phv_data_105 : _GEN_10869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10871 = 8'h6a == local_offset_5 ? phv_data_106 : _GEN_10870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10872 = 8'h6b == local_offset_5 ? phv_data_107 : _GEN_10871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10873 = 8'h6c == local_offset_5 ? phv_data_108 : _GEN_10872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10874 = 8'h6d == local_offset_5 ? phv_data_109 : _GEN_10873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10875 = 8'h6e == local_offset_5 ? phv_data_110 : _GEN_10874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10876 = 8'h6f == local_offset_5 ? phv_data_111 : _GEN_10875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10877 = 8'h70 == local_offset_5 ? phv_data_112 : _GEN_10876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10878 = 8'h71 == local_offset_5 ? phv_data_113 : _GEN_10877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10879 = 8'h72 == local_offset_5 ? phv_data_114 : _GEN_10878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10880 = 8'h73 == local_offset_5 ? phv_data_115 : _GEN_10879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10881 = 8'h74 == local_offset_5 ? phv_data_116 : _GEN_10880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10882 = 8'h75 == local_offset_5 ? phv_data_117 : _GEN_10881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10883 = 8'h76 == local_offset_5 ? phv_data_118 : _GEN_10882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10884 = 8'h77 == local_offset_5 ? phv_data_119 : _GEN_10883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10885 = 8'h78 == local_offset_5 ? phv_data_120 : _GEN_10884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10886 = 8'h79 == local_offset_5 ? phv_data_121 : _GEN_10885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10887 = 8'h7a == local_offset_5 ? phv_data_122 : _GEN_10886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10888 = 8'h7b == local_offset_5 ? phv_data_123 : _GEN_10887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10889 = 8'h7c == local_offset_5 ? phv_data_124 : _GEN_10888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10890 = 8'h7d == local_offset_5 ? phv_data_125 : _GEN_10889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10891 = 8'h7e == local_offset_5 ? phv_data_126 : _GEN_10890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10892 = 8'h7f == local_offset_5 ? phv_data_127 : _GEN_10891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10893 = 8'h80 == local_offset_5 ? phv_data_128 : _GEN_10892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10894 = 8'h81 == local_offset_5 ? phv_data_129 : _GEN_10893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10895 = 8'h82 == local_offset_5 ? phv_data_130 : _GEN_10894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10896 = 8'h83 == local_offset_5 ? phv_data_131 : _GEN_10895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10897 = 8'h84 == local_offset_5 ? phv_data_132 : _GEN_10896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10898 = 8'h85 == local_offset_5 ? phv_data_133 : _GEN_10897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10899 = 8'h86 == local_offset_5 ? phv_data_134 : _GEN_10898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10900 = 8'h87 == local_offset_5 ? phv_data_135 : _GEN_10899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10901 = 8'h88 == local_offset_5 ? phv_data_136 : _GEN_10900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10902 = 8'h89 == local_offset_5 ? phv_data_137 : _GEN_10901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10903 = 8'h8a == local_offset_5 ? phv_data_138 : _GEN_10902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10904 = 8'h8b == local_offset_5 ? phv_data_139 : _GEN_10903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10905 = 8'h8c == local_offset_5 ? phv_data_140 : _GEN_10904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10906 = 8'h8d == local_offset_5 ? phv_data_141 : _GEN_10905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10907 = 8'h8e == local_offset_5 ? phv_data_142 : _GEN_10906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10908 = 8'h8f == local_offset_5 ? phv_data_143 : _GEN_10907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10909 = 8'h90 == local_offset_5 ? phv_data_144 : _GEN_10908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10910 = 8'h91 == local_offset_5 ? phv_data_145 : _GEN_10909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10911 = 8'h92 == local_offset_5 ? phv_data_146 : _GEN_10910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10912 = 8'h93 == local_offset_5 ? phv_data_147 : _GEN_10911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10913 = 8'h94 == local_offset_5 ? phv_data_148 : _GEN_10912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10914 = 8'h95 == local_offset_5 ? phv_data_149 : _GEN_10913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10915 = 8'h96 == local_offset_5 ? phv_data_150 : _GEN_10914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10916 = 8'h97 == local_offset_5 ? phv_data_151 : _GEN_10915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10917 = 8'h98 == local_offset_5 ? phv_data_152 : _GEN_10916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10918 = 8'h99 == local_offset_5 ? phv_data_153 : _GEN_10917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10919 = 8'h9a == local_offset_5 ? phv_data_154 : _GEN_10918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10920 = 8'h9b == local_offset_5 ? phv_data_155 : _GEN_10919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10921 = 8'h9c == local_offset_5 ? phv_data_156 : _GEN_10920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10922 = 8'h9d == local_offset_5 ? phv_data_157 : _GEN_10921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10923 = 8'h9e == local_offset_5 ? phv_data_158 : _GEN_10922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10924 = 8'h9f == local_offset_5 ? phv_data_159 : _GEN_10923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10925 = 8'ha0 == local_offset_5 ? phv_data_160 : _GEN_10924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10926 = 8'ha1 == local_offset_5 ? phv_data_161 : _GEN_10925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10927 = 8'ha2 == local_offset_5 ? phv_data_162 : _GEN_10926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10928 = 8'ha3 == local_offset_5 ? phv_data_163 : _GEN_10927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10929 = 8'ha4 == local_offset_5 ? phv_data_164 : _GEN_10928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10930 = 8'ha5 == local_offset_5 ? phv_data_165 : _GEN_10929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10931 = 8'ha6 == local_offset_5 ? phv_data_166 : _GEN_10930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10932 = 8'ha7 == local_offset_5 ? phv_data_167 : _GEN_10931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10933 = 8'ha8 == local_offset_5 ? phv_data_168 : _GEN_10932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10934 = 8'ha9 == local_offset_5 ? phv_data_169 : _GEN_10933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10935 = 8'haa == local_offset_5 ? phv_data_170 : _GEN_10934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10936 = 8'hab == local_offset_5 ? phv_data_171 : _GEN_10935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10937 = 8'hac == local_offset_5 ? phv_data_172 : _GEN_10936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10938 = 8'had == local_offset_5 ? phv_data_173 : _GEN_10937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10939 = 8'hae == local_offset_5 ? phv_data_174 : _GEN_10938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10940 = 8'haf == local_offset_5 ? phv_data_175 : _GEN_10939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10941 = 8'hb0 == local_offset_5 ? phv_data_176 : _GEN_10940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10942 = 8'hb1 == local_offset_5 ? phv_data_177 : _GEN_10941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10943 = 8'hb2 == local_offset_5 ? phv_data_178 : _GEN_10942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10944 = 8'hb3 == local_offset_5 ? phv_data_179 : _GEN_10943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10945 = 8'hb4 == local_offset_5 ? phv_data_180 : _GEN_10944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10946 = 8'hb5 == local_offset_5 ? phv_data_181 : _GEN_10945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10947 = 8'hb6 == local_offset_5 ? phv_data_182 : _GEN_10946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10948 = 8'hb7 == local_offset_5 ? phv_data_183 : _GEN_10947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10949 = 8'hb8 == local_offset_5 ? phv_data_184 : _GEN_10948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10950 = 8'hb9 == local_offset_5 ? phv_data_185 : _GEN_10949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10951 = 8'hba == local_offset_5 ? phv_data_186 : _GEN_10950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10952 = 8'hbb == local_offset_5 ? phv_data_187 : _GEN_10951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10953 = 8'hbc == local_offset_5 ? phv_data_188 : _GEN_10952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10954 = 8'hbd == local_offset_5 ? phv_data_189 : _GEN_10953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10955 = 8'hbe == local_offset_5 ? phv_data_190 : _GEN_10954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10956 = 8'hbf == local_offset_5 ? phv_data_191 : _GEN_10955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10957 = 8'hc0 == local_offset_5 ? phv_data_192 : _GEN_10956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10958 = 8'hc1 == local_offset_5 ? phv_data_193 : _GEN_10957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10959 = 8'hc2 == local_offset_5 ? phv_data_194 : _GEN_10958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10960 = 8'hc3 == local_offset_5 ? phv_data_195 : _GEN_10959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10961 = 8'hc4 == local_offset_5 ? phv_data_196 : _GEN_10960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10962 = 8'hc5 == local_offset_5 ? phv_data_197 : _GEN_10961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10963 = 8'hc6 == local_offset_5 ? phv_data_198 : _GEN_10962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10964 = 8'hc7 == local_offset_5 ? phv_data_199 : _GEN_10963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10965 = 8'hc8 == local_offset_5 ? phv_data_200 : _GEN_10964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10966 = 8'hc9 == local_offset_5 ? phv_data_201 : _GEN_10965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10967 = 8'hca == local_offset_5 ? phv_data_202 : _GEN_10966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10968 = 8'hcb == local_offset_5 ? phv_data_203 : _GEN_10967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10969 = 8'hcc == local_offset_5 ? phv_data_204 : _GEN_10968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10970 = 8'hcd == local_offset_5 ? phv_data_205 : _GEN_10969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10971 = 8'hce == local_offset_5 ? phv_data_206 : _GEN_10970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10972 = 8'hcf == local_offset_5 ? phv_data_207 : _GEN_10971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10973 = 8'hd0 == local_offset_5 ? phv_data_208 : _GEN_10972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10974 = 8'hd1 == local_offset_5 ? phv_data_209 : _GEN_10973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10975 = 8'hd2 == local_offset_5 ? phv_data_210 : _GEN_10974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10976 = 8'hd3 == local_offset_5 ? phv_data_211 : _GEN_10975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10977 = 8'hd4 == local_offset_5 ? phv_data_212 : _GEN_10976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10978 = 8'hd5 == local_offset_5 ? phv_data_213 : _GEN_10977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10979 = 8'hd6 == local_offset_5 ? phv_data_214 : _GEN_10978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10980 = 8'hd7 == local_offset_5 ? phv_data_215 : _GEN_10979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10981 = 8'hd8 == local_offset_5 ? phv_data_216 : _GEN_10980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10982 = 8'hd9 == local_offset_5 ? phv_data_217 : _GEN_10981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10983 = 8'hda == local_offset_5 ? phv_data_218 : _GEN_10982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10984 = 8'hdb == local_offset_5 ? phv_data_219 : _GEN_10983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10985 = 8'hdc == local_offset_5 ? phv_data_220 : _GEN_10984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10986 = 8'hdd == local_offset_5 ? phv_data_221 : _GEN_10985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10987 = 8'hde == local_offset_5 ? phv_data_222 : _GEN_10986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10988 = 8'hdf == local_offset_5 ? phv_data_223 : _GEN_10987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10989 = 8'he0 == local_offset_5 ? phv_data_224 : _GEN_10988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10990 = 8'he1 == local_offset_5 ? phv_data_225 : _GEN_10989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10991 = 8'he2 == local_offset_5 ? phv_data_226 : _GEN_10990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10992 = 8'he3 == local_offset_5 ? phv_data_227 : _GEN_10991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10993 = 8'he4 == local_offset_5 ? phv_data_228 : _GEN_10992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10994 = 8'he5 == local_offset_5 ? phv_data_229 : _GEN_10993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10995 = 8'he6 == local_offset_5 ? phv_data_230 : _GEN_10994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10996 = 8'he7 == local_offset_5 ? phv_data_231 : _GEN_10995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10997 = 8'he8 == local_offset_5 ? phv_data_232 : _GEN_10996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10998 = 8'he9 == local_offset_5 ? phv_data_233 : _GEN_10997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10999 = 8'hea == local_offset_5 ? phv_data_234 : _GEN_10998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11000 = 8'heb == local_offset_5 ? phv_data_235 : _GEN_10999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11001 = 8'hec == local_offset_5 ? phv_data_236 : _GEN_11000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11002 = 8'hed == local_offset_5 ? phv_data_237 : _GEN_11001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11003 = 8'hee == local_offset_5 ? phv_data_238 : _GEN_11002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11004 = 8'hef == local_offset_5 ? phv_data_239 : _GEN_11003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11005 = 8'hf0 == local_offset_5 ? phv_data_240 : _GEN_11004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11006 = 8'hf1 == local_offset_5 ? phv_data_241 : _GEN_11005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11007 = 8'hf2 == local_offset_5 ? phv_data_242 : _GEN_11006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11008 = 8'hf3 == local_offset_5 ? phv_data_243 : _GEN_11007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11009 = 8'hf4 == local_offset_5 ? phv_data_244 : _GEN_11008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11010 = 8'hf5 == local_offset_5 ? phv_data_245 : _GEN_11009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11011 = 8'hf6 == local_offset_5 ? phv_data_246 : _GEN_11010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11012 = 8'hf7 == local_offset_5 ? phv_data_247 : _GEN_11011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11013 = 8'hf8 == local_offset_5 ? phv_data_248 : _GEN_11012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11014 = 8'hf9 == local_offset_5 ? phv_data_249 : _GEN_11013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11015 = 8'hfa == local_offset_5 ? phv_data_250 : _GEN_11014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11016 = 8'hfb == local_offset_5 ? phv_data_251 : _GEN_11015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11017 = 8'hfc == local_offset_5 ? phv_data_252 : _GEN_11016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11018 = 8'hfd == local_offset_5 ? phv_data_253 : _GEN_11017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11019 = 8'hfe == local_offset_5 ? phv_data_254 : _GEN_11018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11020 = 8'hff == local_offset_5 ? phv_data_255 : _GEN_11019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_17702 = {{1'd0}, local_offset_5}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11021 = 9'h100 == _GEN_17702 ? phv_data_256 : _GEN_11020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11022 = 9'h101 == _GEN_17702 ? phv_data_257 : _GEN_11021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11023 = 9'h102 == _GEN_17702 ? phv_data_258 : _GEN_11022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11024 = 9'h103 == _GEN_17702 ? phv_data_259 : _GEN_11023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11025 = 9'h104 == _GEN_17702 ? phv_data_260 : _GEN_11024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11026 = 9'h105 == _GEN_17702 ? phv_data_261 : _GEN_11025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11027 = 9'h106 == _GEN_17702 ? phv_data_262 : _GEN_11026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11028 = 9'h107 == _GEN_17702 ? phv_data_263 : _GEN_11027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11029 = 9'h108 == _GEN_17702 ? phv_data_264 : _GEN_11028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11030 = 9'h109 == _GEN_17702 ? phv_data_265 : _GEN_11029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11031 = 9'h10a == _GEN_17702 ? phv_data_266 : _GEN_11030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11032 = 9'h10b == _GEN_17702 ? phv_data_267 : _GEN_11031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11033 = 9'h10c == _GEN_17702 ? phv_data_268 : _GEN_11032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11034 = 9'h10d == _GEN_17702 ? phv_data_269 : _GEN_11033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11035 = 9'h10e == _GEN_17702 ? phv_data_270 : _GEN_11034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11036 = 9'h10f == _GEN_17702 ? phv_data_271 : _GEN_11035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11037 = 9'h110 == _GEN_17702 ? phv_data_272 : _GEN_11036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11038 = 9'h111 == _GEN_17702 ? phv_data_273 : _GEN_11037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11039 = 9'h112 == _GEN_17702 ? phv_data_274 : _GEN_11038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11040 = 9'h113 == _GEN_17702 ? phv_data_275 : _GEN_11039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11041 = 9'h114 == _GEN_17702 ? phv_data_276 : _GEN_11040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11042 = 9'h115 == _GEN_17702 ? phv_data_277 : _GEN_11041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11043 = 9'h116 == _GEN_17702 ? phv_data_278 : _GEN_11042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11044 = 9'h117 == _GEN_17702 ? phv_data_279 : _GEN_11043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11045 = 9'h118 == _GEN_17702 ? phv_data_280 : _GEN_11044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11046 = 9'h119 == _GEN_17702 ? phv_data_281 : _GEN_11045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11047 = 9'h11a == _GEN_17702 ? phv_data_282 : _GEN_11046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11048 = 9'h11b == _GEN_17702 ? phv_data_283 : _GEN_11047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11049 = 9'h11c == _GEN_17702 ? phv_data_284 : _GEN_11048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11050 = 9'h11d == _GEN_17702 ? phv_data_285 : _GEN_11049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11051 = 9'h11e == _GEN_17702 ? phv_data_286 : _GEN_11050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11052 = 9'h11f == _GEN_17702 ? phv_data_287 : _GEN_11051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11053 = 9'h120 == _GEN_17702 ? phv_data_288 : _GEN_11052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11054 = 9'h121 == _GEN_17702 ? phv_data_289 : _GEN_11053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11055 = 9'h122 == _GEN_17702 ? phv_data_290 : _GEN_11054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11056 = 9'h123 == _GEN_17702 ? phv_data_291 : _GEN_11055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11057 = 9'h124 == _GEN_17702 ? phv_data_292 : _GEN_11056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11058 = 9'h125 == _GEN_17702 ? phv_data_293 : _GEN_11057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11059 = 9'h126 == _GEN_17702 ? phv_data_294 : _GEN_11058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11060 = 9'h127 == _GEN_17702 ? phv_data_295 : _GEN_11059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11061 = 9'h128 == _GEN_17702 ? phv_data_296 : _GEN_11060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11062 = 9'h129 == _GEN_17702 ? phv_data_297 : _GEN_11061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11063 = 9'h12a == _GEN_17702 ? phv_data_298 : _GEN_11062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11064 = 9'h12b == _GEN_17702 ? phv_data_299 : _GEN_11063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11065 = 9'h12c == _GEN_17702 ? phv_data_300 : _GEN_11064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11066 = 9'h12d == _GEN_17702 ? phv_data_301 : _GEN_11065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11067 = 9'h12e == _GEN_17702 ? phv_data_302 : _GEN_11066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11068 = 9'h12f == _GEN_17702 ? phv_data_303 : _GEN_11067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11069 = 9'h130 == _GEN_17702 ? phv_data_304 : _GEN_11068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11070 = 9'h131 == _GEN_17702 ? phv_data_305 : _GEN_11069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11071 = 9'h132 == _GEN_17702 ? phv_data_306 : _GEN_11070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11072 = 9'h133 == _GEN_17702 ? phv_data_307 : _GEN_11071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11073 = 9'h134 == _GEN_17702 ? phv_data_308 : _GEN_11072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11074 = 9'h135 == _GEN_17702 ? phv_data_309 : _GEN_11073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11075 = 9'h136 == _GEN_17702 ? phv_data_310 : _GEN_11074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11076 = 9'h137 == _GEN_17702 ? phv_data_311 : _GEN_11075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11077 = 9'h138 == _GEN_17702 ? phv_data_312 : _GEN_11076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11078 = 9'h139 == _GEN_17702 ? phv_data_313 : _GEN_11077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11079 = 9'h13a == _GEN_17702 ? phv_data_314 : _GEN_11078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11080 = 9'h13b == _GEN_17702 ? phv_data_315 : _GEN_11079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11081 = 9'h13c == _GEN_17702 ? phv_data_316 : _GEN_11080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11082 = 9'h13d == _GEN_17702 ? phv_data_317 : _GEN_11081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11083 = 9'h13e == _GEN_17702 ? phv_data_318 : _GEN_11082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11084 = 9'h13f == _GEN_17702 ? phv_data_319 : _GEN_11083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11085 = 9'h140 == _GEN_17702 ? phv_data_320 : _GEN_11084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11086 = 9'h141 == _GEN_17702 ? phv_data_321 : _GEN_11085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11087 = 9'h142 == _GEN_17702 ? phv_data_322 : _GEN_11086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11088 = 9'h143 == _GEN_17702 ? phv_data_323 : _GEN_11087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11089 = 9'h144 == _GEN_17702 ? phv_data_324 : _GEN_11088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11090 = 9'h145 == _GEN_17702 ? phv_data_325 : _GEN_11089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11091 = 9'h146 == _GEN_17702 ? phv_data_326 : _GEN_11090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11092 = 9'h147 == _GEN_17702 ? phv_data_327 : _GEN_11091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11093 = 9'h148 == _GEN_17702 ? phv_data_328 : _GEN_11092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11094 = 9'h149 == _GEN_17702 ? phv_data_329 : _GEN_11093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11095 = 9'h14a == _GEN_17702 ? phv_data_330 : _GEN_11094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11096 = 9'h14b == _GEN_17702 ? phv_data_331 : _GEN_11095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11097 = 9'h14c == _GEN_17702 ? phv_data_332 : _GEN_11096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11098 = 9'h14d == _GEN_17702 ? phv_data_333 : _GEN_11097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11099 = 9'h14e == _GEN_17702 ? phv_data_334 : _GEN_11098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11100 = 9'h14f == _GEN_17702 ? phv_data_335 : _GEN_11099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11101 = 9'h150 == _GEN_17702 ? phv_data_336 : _GEN_11100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11102 = 9'h151 == _GEN_17702 ? phv_data_337 : _GEN_11101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11103 = 9'h152 == _GEN_17702 ? phv_data_338 : _GEN_11102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11104 = 9'h153 == _GEN_17702 ? phv_data_339 : _GEN_11103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11105 = 9'h154 == _GEN_17702 ? phv_data_340 : _GEN_11104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11106 = 9'h155 == _GEN_17702 ? phv_data_341 : _GEN_11105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11107 = 9'h156 == _GEN_17702 ? phv_data_342 : _GEN_11106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11108 = 9'h157 == _GEN_17702 ? phv_data_343 : _GEN_11107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11109 = 9'h158 == _GEN_17702 ? phv_data_344 : _GEN_11108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11110 = 9'h159 == _GEN_17702 ? phv_data_345 : _GEN_11109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11111 = 9'h15a == _GEN_17702 ? phv_data_346 : _GEN_11110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11112 = 9'h15b == _GEN_17702 ? phv_data_347 : _GEN_11111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11113 = 9'h15c == _GEN_17702 ? phv_data_348 : _GEN_11112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11114 = 9'h15d == _GEN_17702 ? phv_data_349 : _GEN_11113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11115 = 9'h15e == _GEN_17702 ? phv_data_350 : _GEN_11114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11116 = 9'h15f == _GEN_17702 ? phv_data_351 : _GEN_11115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11117 = 9'h160 == _GEN_17702 ? phv_data_352 : _GEN_11116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11118 = 9'h161 == _GEN_17702 ? phv_data_353 : _GEN_11117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11119 = 9'h162 == _GEN_17702 ? phv_data_354 : _GEN_11118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11120 = 9'h163 == _GEN_17702 ? phv_data_355 : _GEN_11119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11121 = 9'h164 == _GEN_17702 ? phv_data_356 : _GEN_11120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11122 = 9'h165 == _GEN_17702 ? phv_data_357 : _GEN_11121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11123 = 9'h166 == _GEN_17702 ? phv_data_358 : _GEN_11122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11124 = 9'h167 == _GEN_17702 ? phv_data_359 : _GEN_11123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11125 = 9'h168 == _GEN_17702 ? phv_data_360 : _GEN_11124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11126 = 9'h169 == _GEN_17702 ? phv_data_361 : _GEN_11125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11127 = 9'h16a == _GEN_17702 ? phv_data_362 : _GEN_11126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11128 = 9'h16b == _GEN_17702 ? phv_data_363 : _GEN_11127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11129 = 9'h16c == _GEN_17702 ? phv_data_364 : _GEN_11128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11130 = 9'h16d == _GEN_17702 ? phv_data_365 : _GEN_11129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11131 = 9'h16e == _GEN_17702 ? phv_data_366 : _GEN_11130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11132 = 9'h16f == _GEN_17702 ? phv_data_367 : _GEN_11131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11133 = 9'h170 == _GEN_17702 ? phv_data_368 : _GEN_11132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11134 = 9'h171 == _GEN_17702 ? phv_data_369 : _GEN_11133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11135 = 9'h172 == _GEN_17702 ? phv_data_370 : _GEN_11134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11136 = 9'h173 == _GEN_17702 ? phv_data_371 : _GEN_11135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11137 = 9'h174 == _GEN_17702 ? phv_data_372 : _GEN_11136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11138 = 9'h175 == _GEN_17702 ? phv_data_373 : _GEN_11137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11139 = 9'h176 == _GEN_17702 ? phv_data_374 : _GEN_11138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11140 = 9'h177 == _GEN_17702 ? phv_data_375 : _GEN_11139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11141 = 9'h178 == _GEN_17702 ? phv_data_376 : _GEN_11140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11142 = 9'h179 == _GEN_17702 ? phv_data_377 : _GEN_11141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11143 = 9'h17a == _GEN_17702 ? phv_data_378 : _GEN_11142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11144 = 9'h17b == _GEN_17702 ? phv_data_379 : _GEN_11143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11145 = 9'h17c == _GEN_17702 ? phv_data_380 : _GEN_11144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11146 = 9'h17d == _GEN_17702 ? phv_data_381 : _GEN_11145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11147 = 9'h17e == _GEN_17702 ? phv_data_382 : _GEN_11146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11148 = 9'h17f == _GEN_17702 ? phv_data_383 : _GEN_11147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11149 = 9'h180 == _GEN_17702 ? phv_data_384 : _GEN_11148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11150 = 9'h181 == _GEN_17702 ? phv_data_385 : _GEN_11149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11151 = 9'h182 == _GEN_17702 ? phv_data_386 : _GEN_11150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11152 = 9'h183 == _GEN_17702 ? phv_data_387 : _GEN_11151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11153 = 9'h184 == _GEN_17702 ? phv_data_388 : _GEN_11152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11154 = 9'h185 == _GEN_17702 ? phv_data_389 : _GEN_11153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11155 = 9'h186 == _GEN_17702 ? phv_data_390 : _GEN_11154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11156 = 9'h187 == _GEN_17702 ? phv_data_391 : _GEN_11155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11157 = 9'h188 == _GEN_17702 ? phv_data_392 : _GEN_11156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11158 = 9'h189 == _GEN_17702 ? phv_data_393 : _GEN_11157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11159 = 9'h18a == _GEN_17702 ? phv_data_394 : _GEN_11158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11160 = 9'h18b == _GEN_17702 ? phv_data_395 : _GEN_11159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11161 = 9'h18c == _GEN_17702 ? phv_data_396 : _GEN_11160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11162 = 9'h18d == _GEN_17702 ? phv_data_397 : _GEN_11161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11163 = 9'h18e == _GEN_17702 ? phv_data_398 : _GEN_11162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11164 = 9'h18f == _GEN_17702 ? phv_data_399 : _GEN_11163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11165 = 9'h190 == _GEN_17702 ? phv_data_400 : _GEN_11164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11166 = 9'h191 == _GEN_17702 ? phv_data_401 : _GEN_11165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11167 = 9'h192 == _GEN_17702 ? phv_data_402 : _GEN_11166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11168 = 9'h193 == _GEN_17702 ? phv_data_403 : _GEN_11167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11169 = 9'h194 == _GEN_17702 ? phv_data_404 : _GEN_11168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11170 = 9'h195 == _GEN_17702 ? phv_data_405 : _GEN_11169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11171 = 9'h196 == _GEN_17702 ? phv_data_406 : _GEN_11170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11172 = 9'h197 == _GEN_17702 ? phv_data_407 : _GEN_11171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11173 = 9'h198 == _GEN_17702 ? phv_data_408 : _GEN_11172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11174 = 9'h199 == _GEN_17702 ? phv_data_409 : _GEN_11173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11175 = 9'h19a == _GEN_17702 ? phv_data_410 : _GEN_11174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11176 = 9'h19b == _GEN_17702 ? phv_data_411 : _GEN_11175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11177 = 9'h19c == _GEN_17702 ? phv_data_412 : _GEN_11176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11178 = 9'h19d == _GEN_17702 ? phv_data_413 : _GEN_11177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11179 = 9'h19e == _GEN_17702 ? phv_data_414 : _GEN_11178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11180 = 9'h19f == _GEN_17702 ? phv_data_415 : _GEN_11179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11181 = 9'h1a0 == _GEN_17702 ? phv_data_416 : _GEN_11180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11182 = 9'h1a1 == _GEN_17702 ? phv_data_417 : _GEN_11181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11183 = 9'h1a2 == _GEN_17702 ? phv_data_418 : _GEN_11182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11184 = 9'h1a3 == _GEN_17702 ? phv_data_419 : _GEN_11183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11185 = 9'h1a4 == _GEN_17702 ? phv_data_420 : _GEN_11184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11186 = 9'h1a5 == _GEN_17702 ? phv_data_421 : _GEN_11185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11187 = 9'h1a6 == _GEN_17702 ? phv_data_422 : _GEN_11186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11188 = 9'h1a7 == _GEN_17702 ? phv_data_423 : _GEN_11187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11189 = 9'h1a8 == _GEN_17702 ? phv_data_424 : _GEN_11188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11190 = 9'h1a9 == _GEN_17702 ? phv_data_425 : _GEN_11189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11191 = 9'h1aa == _GEN_17702 ? phv_data_426 : _GEN_11190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11192 = 9'h1ab == _GEN_17702 ? phv_data_427 : _GEN_11191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11193 = 9'h1ac == _GEN_17702 ? phv_data_428 : _GEN_11192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11194 = 9'h1ad == _GEN_17702 ? phv_data_429 : _GEN_11193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11195 = 9'h1ae == _GEN_17702 ? phv_data_430 : _GEN_11194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11196 = 9'h1af == _GEN_17702 ? phv_data_431 : _GEN_11195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11197 = 9'h1b0 == _GEN_17702 ? phv_data_432 : _GEN_11196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11198 = 9'h1b1 == _GEN_17702 ? phv_data_433 : _GEN_11197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11199 = 9'h1b2 == _GEN_17702 ? phv_data_434 : _GEN_11198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11200 = 9'h1b3 == _GEN_17702 ? phv_data_435 : _GEN_11199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11201 = 9'h1b4 == _GEN_17702 ? phv_data_436 : _GEN_11200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11202 = 9'h1b5 == _GEN_17702 ? phv_data_437 : _GEN_11201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11203 = 9'h1b6 == _GEN_17702 ? phv_data_438 : _GEN_11202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11204 = 9'h1b7 == _GEN_17702 ? phv_data_439 : _GEN_11203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11205 = 9'h1b8 == _GEN_17702 ? phv_data_440 : _GEN_11204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11206 = 9'h1b9 == _GEN_17702 ? phv_data_441 : _GEN_11205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11207 = 9'h1ba == _GEN_17702 ? phv_data_442 : _GEN_11206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11208 = 9'h1bb == _GEN_17702 ? phv_data_443 : _GEN_11207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11209 = 9'h1bc == _GEN_17702 ? phv_data_444 : _GEN_11208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11210 = 9'h1bd == _GEN_17702 ? phv_data_445 : _GEN_11209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11211 = 9'h1be == _GEN_17702 ? phv_data_446 : _GEN_11210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11212 = 9'h1bf == _GEN_17702 ? phv_data_447 : _GEN_11211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11213 = 9'h1c0 == _GEN_17702 ? phv_data_448 : _GEN_11212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11214 = 9'h1c1 == _GEN_17702 ? phv_data_449 : _GEN_11213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11215 = 9'h1c2 == _GEN_17702 ? phv_data_450 : _GEN_11214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11216 = 9'h1c3 == _GEN_17702 ? phv_data_451 : _GEN_11215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11217 = 9'h1c4 == _GEN_17702 ? phv_data_452 : _GEN_11216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11218 = 9'h1c5 == _GEN_17702 ? phv_data_453 : _GEN_11217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11219 = 9'h1c6 == _GEN_17702 ? phv_data_454 : _GEN_11218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11220 = 9'h1c7 == _GEN_17702 ? phv_data_455 : _GEN_11219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11221 = 9'h1c8 == _GEN_17702 ? phv_data_456 : _GEN_11220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11222 = 9'h1c9 == _GEN_17702 ? phv_data_457 : _GEN_11221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11223 = 9'h1ca == _GEN_17702 ? phv_data_458 : _GEN_11222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11224 = 9'h1cb == _GEN_17702 ? phv_data_459 : _GEN_11223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11225 = 9'h1cc == _GEN_17702 ? phv_data_460 : _GEN_11224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11226 = 9'h1cd == _GEN_17702 ? phv_data_461 : _GEN_11225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11227 = 9'h1ce == _GEN_17702 ? phv_data_462 : _GEN_11226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11228 = 9'h1cf == _GEN_17702 ? phv_data_463 : _GEN_11227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11229 = 9'h1d0 == _GEN_17702 ? phv_data_464 : _GEN_11228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11230 = 9'h1d1 == _GEN_17702 ? phv_data_465 : _GEN_11229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11231 = 9'h1d2 == _GEN_17702 ? phv_data_466 : _GEN_11230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11232 = 9'h1d3 == _GEN_17702 ? phv_data_467 : _GEN_11231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11233 = 9'h1d4 == _GEN_17702 ? phv_data_468 : _GEN_11232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11234 = 9'h1d5 == _GEN_17702 ? phv_data_469 : _GEN_11233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11235 = 9'h1d6 == _GEN_17702 ? phv_data_470 : _GEN_11234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11236 = 9'h1d7 == _GEN_17702 ? phv_data_471 : _GEN_11235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11237 = 9'h1d8 == _GEN_17702 ? phv_data_472 : _GEN_11236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11238 = 9'h1d9 == _GEN_17702 ? phv_data_473 : _GEN_11237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11239 = 9'h1da == _GEN_17702 ? phv_data_474 : _GEN_11238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11240 = 9'h1db == _GEN_17702 ? phv_data_475 : _GEN_11239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11241 = 9'h1dc == _GEN_17702 ? phv_data_476 : _GEN_11240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11242 = 9'h1dd == _GEN_17702 ? phv_data_477 : _GEN_11241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11243 = 9'h1de == _GEN_17702 ? phv_data_478 : _GEN_11242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11244 = 9'h1df == _GEN_17702 ? phv_data_479 : _GEN_11243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11245 = 9'h1e0 == _GEN_17702 ? phv_data_480 : _GEN_11244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11246 = 9'h1e1 == _GEN_17702 ? phv_data_481 : _GEN_11245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11247 = 9'h1e2 == _GEN_17702 ? phv_data_482 : _GEN_11246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11248 = 9'h1e3 == _GEN_17702 ? phv_data_483 : _GEN_11247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11249 = 9'h1e4 == _GEN_17702 ? phv_data_484 : _GEN_11248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11250 = 9'h1e5 == _GEN_17702 ? phv_data_485 : _GEN_11249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11251 = 9'h1e6 == _GEN_17702 ? phv_data_486 : _GEN_11250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11252 = 9'h1e7 == _GEN_17702 ? phv_data_487 : _GEN_11251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11253 = 9'h1e8 == _GEN_17702 ? phv_data_488 : _GEN_11252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11254 = 9'h1e9 == _GEN_17702 ? phv_data_489 : _GEN_11253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11255 = 9'h1ea == _GEN_17702 ? phv_data_490 : _GEN_11254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11256 = 9'h1eb == _GEN_17702 ? phv_data_491 : _GEN_11255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11257 = 9'h1ec == _GEN_17702 ? phv_data_492 : _GEN_11256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11258 = 9'h1ed == _GEN_17702 ? phv_data_493 : _GEN_11257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11259 = 9'h1ee == _GEN_17702 ? phv_data_494 : _GEN_11258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11260 = 9'h1ef == _GEN_17702 ? phv_data_495 : _GEN_11259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11261 = 9'h1f0 == _GEN_17702 ? phv_data_496 : _GEN_11260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11262 = 9'h1f1 == _GEN_17702 ? phv_data_497 : _GEN_11261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11263 = 9'h1f2 == _GEN_17702 ? phv_data_498 : _GEN_11262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11264 = 9'h1f3 == _GEN_17702 ? phv_data_499 : _GEN_11263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11265 = 9'h1f4 == _GEN_17702 ? phv_data_500 : _GEN_11264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11266 = 9'h1f5 == _GEN_17702 ? phv_data_501 : _GEN_11265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11267 = 9'h1f6 == _GEN_17702 ? phv_data_502 : _GEN_11266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11268 = 9'h1f7 == _GEN_17702 ? phv_data_503 : _GEN_11267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11269 = 9'h1f8 == _GEN_17702 ? phv_data_504 : _GEN_11268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11270 = 9'h1f9 == _GEN_17702 ? phv_data_505 : _GEN_11269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11271 = 9'h1fa == _GEN_17702 ? phv_data_506 : _GEN_11270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11272 = 9'h1fb == _GEN_17702 ? phv_data_507 : _GEN_11271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11273 = 9'h1fc == _GEN_17702 ? phv_data_508 : _GEN_11272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11274 = 9'h1fd == _GEN_17702 ? phv_data_509 : _GEN_11273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11275 = 9'h1fe == _GEN_17702 ? phv_data_510 : _GEN_11274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11276 = 9'h1ff == _GEN_17702 ? phv_data_511 : _GEN_11275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11278 = 8'h1 == _match_key_qbytes_5_T ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11279 = 8'h2 == _match_key_qbytes_5_T ? phv_data_2 : _GEN_11278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11280 = 8'h3 == _match_key_qbytes_5_T ? phv_data_3 : _GEN_11279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11281 = 8'h4 == _match_key_qbytes_5_T ? phv_data_4 : _GEN_11280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11282 = 8'h5 == _match_key_qbytes_5_T ? phv_data_5 : _GEN_11281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11283 = 8'h6 == _match_key_qbytes_5_T ? phv_data_6 : _GEN_11282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11284 = 8'h7 == _match_key_qbytes_5_T ? phv_data_7 : _GEN_11283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11285 = 8'h8 == _match_key_qbytes_5_T ? phv_data_8 : _GEN_11284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11286 = 8'h9 == _match_key_qbytes_5_T ? phv_data_9 : _GEN_11285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11287 = 8'ha == _match_key_qbytes_5_T ? phv_data_10 : _GEN_11286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11288 = 8'hb == _match_key_qbytes_5_T ? phv_data_11 : _GEN_11287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11289 = 8'hc == _match_key_qbytes_5_T ? phv_data_12 : _GEN_11288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11290 = 8'hd == _match_key_qbytes_5_T ? phv_data_13 : _GEN_11289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11291 = 8'he == _match_key_qbytes_5_T ? phv_data_14 : _GEN_11290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11292 = 8'hf == _match_key_qbytes_5_T ? phv_data_15 : _GEN_11291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11293 = 8'h10 == _match_key_qbytes_5_T ? phv_data_16 : _GEN_11292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11294 = 8'h11 == _match_key_qbytes_5_T ? phv_data_17 : _GEN_11293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11295 = 8'h12 == _match_key_qbytes_5_T ? phv_data_18 : _GEN_11294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11296 = 8'h13 == _match_key_qbytes_5_T ? phv_data_19 : _GEN_11295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11297 = 8'h14 == _match_key_qbytes_5_T ? phv_data_20 : _GEN_11296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11298 = 8'h15 == _match_key_qbytes_5_T ? phv_data_21 : _GEN_11297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11299 = 8'h16 == _match_key_qbytes_5_T ? phv_data_22 : _GEN_11298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11300 = 8'h17 == _match_key_qbytes_5_T ? phv_data_23 : _GEN_11299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11301 = 8'h18 == _match_key_qbytes_5_T ? phv_data_24 : _GEN_11300; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11302 = 8'h19 == _match_key_qbytes_5_T ? phv_data_25 : _GEN_11301; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11303 = 8'h1a == _match_key_qbytes_5_T ? phv_data_26 : _GEN_11302; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11304 = 8'h1b == _match_key_qbytes_5_T ? phv_data_27 : _GEN_11303; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11305 = 8'h1c == _match_key_qbytes_5_T ? phv_data_28 : _GEN_11304; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11306 = 8'h1d == _match_key_qbytes_5_T ? phv_data_29 : _GEN_11305; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11307 = 8'h1e == _match_key_qbytes_5_T ? phv_data_30 : _GEN_11306; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11308 = 8'h1f == _match_key_qbytes_5_T ? phv_data_31 : _GEN_11307; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11309 = 8'h20 == _match_key_qbytes_5_T ? phv_data_32 : _GEN_11308; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11310 = 8'h21 == _match_key_qbytes_5_T ? phv_data_33 : _GEN_11309; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11311 = 8'h22 == _match_key_qbytes_5_T ? phv_data_34 : _GEN_11310; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11312 = 8'h23 == _match_key_qbytes_5_T ? phv_data_35 : _GEN_11311; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11313 = 8'h24 == _match_key_qbytes_5_T ? phv_data_36 : _GEN_11312; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11314 = 8'h25 == _match_key_qbytes_5_T ? phv_data_37 : _GEN_11313; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11315 = 8'h26 == _match_key_qbytes_5_T ? phv_data_38 : _GEN_11314; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11316 = 8'h27 == _match_key_qbytes_5_T ? phv_data_39 : _GEN_11315; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11317 = 8'h28 == _match_key_qbytes_5_T ? phv_data_40 : _GEN_11316; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11318 = 8'h29 == _match_key_qbytes_5_T ? phv_data_41 : _GEN_11317; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11319 = 8'h2a == _match_key_qbytes_5_T ? phv_data_42 : _GEN_11318; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11320 = 8'h2b == _match_key_qbytes_5_T ? phv_data_43 : _GEN_11319; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11321 = 8'h2c == _match_key_qbytes_5_T ? phv_data_44 : _GEN_11320; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11322 = 8'h2d == _match_key_qbytes_5_T ? phv_data_45 : _GEN_11321; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11323 = 8'h2e == _match_key_qbytes_5_T ? phv_data_46 : _GEN_11322; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11324 = 8'h2f == _match_key_qbytes_5_T ? phv_data_47 : _GEN_11323; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11325 = 8'h30 == _match_key_qbytes_5_T ? phv_data_48 : _GEN_11324; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11326 = 8'h31 == _match_key_qbytes_5_T ? phv_data_49 : _GEN_11325; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11327 = 8'h32 == _match_key_qbytes_5_T ? phv_data_50 : _GEN_11326; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11328 = 8'h33 == _match_key_qbytes_5_T ? phv_data_51 : _GEN_11327; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11329 = 8'h34 == _match_key_qbytes_5_T ? phv_data_52 : _GEN_11328; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11330 = 8'h35 == _match_key_qbytes_5_T ? phv_data_53 : _GEN_11329; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11331 = 8'h36 == _match_key_qbytes_5_T ? phv_data_54 : _GEN_11330; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11332 = 8'h37 == _match_key_qbytes_5_T ? phv_data_55 : _GEN_11331; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11333 = 8'h38 == _match_key_qbytes_5_T ? phv_data_56 : _GEN_11332; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11334 = 8'h39 == _match_key_qbytes_5_T ? phv_data_57 : _GEN_11333; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11335 = 8'h3a == _match_key_qbytes_5_T ? phv_data_58 : _GEN_11334; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11336 = 8'h3b == _match_key_qbytes_5_T ? phv_data_59 : _GEN_11335; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11337 = 8'h3c == _match_key_qbytes_5_T ? phv_data_60 : _GEN_11336; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11338 = 8'h3d == _match_key_qbytes_5_T ? phv_data_61 : _GEN_11337; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11339 = 8'h3e == _match_key_qbytes_5_T ? phv_data_62 : _GEN_11338; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11340 = 8'h3f == _match_key_qbytes_5_T ? phv_data_63 : _GEN_11339; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11341 = 8'h40 == _match_key_qbytes_5_T ? phv_data_64 : _GEN_11340; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11342 = 8'h41 == _match_key_qbytes_5_T ? phv_data_65 : _GEN_11341; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11343 = 8'h42 == _match_key_qbytes_5_T ? phv_data_66 : _GEN_11342; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11344 = 8'h43 == _match_key_qbytes_5_T ? phv_data_67 : _GEN_11343; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11345 = 8'h44 == _match_key_qbytes_5_T ? phv_data_68 : _GEN_11344; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11346 = 8'h45 == _match_key_qbytes_5_T ? phv_data_69 : _GEN_11345; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11347 = 8'h46 == _match_key_qbytes_5_T ? phv_data_70 : _GEN_11346; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11348 = 8'h47 == _match_key_qbytes_5_T ? phv_data_71 : _GEN_11347; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11349 = 8'h48 == _match_key_qbytes_5_T ? phv_data_72 : _GEN_11348; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11350 = 8'h49 == _match_key_qbytes_5_T ? phv_data_73 : _GEN_11349; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11351 = 8'h4a == _match_key_qbytes_5_T ? phv_data_74 : _GEN_11350; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11352 = 8'h4b == _match_key_qbytes_5_T ? phv_data_75 : _GEN_11351; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11353 = 8'h4c == _match_key_qbytes_5_T ? phv_data_76 : _GEN_11352; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11354 = 8'h4d == _match_key_qbytes_5_T ? phv_data_77 : _GEN_11353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11355 = 8'h4e == _match_key_qbytes_5_T ? phv_data_78 : _GEN_11354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11356 = 8'h4f == _match_key_qbytes_5_T ? phv_data_79 : _GEN_11355; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11357 = 8'h50 == _match_key_qbytes_5_T ? phv_data_80 : _GEN_11356; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11358 = 8'h51 == _match_key_qbytes_5_T ? phv_data_81 : _GEN_11357; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11359 = 8'h52 == _match_key_qbytes_5_T ? phv_data_82 : _GEN_11358; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11360 = 8'h53 == _match_key_qbytes_5_T ? phv_data_83 : _GEN_11359; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11361 = 8'h54 == _match_key_qbytes_5_T ? phv_data_84 : _GEN_11360; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11362 = 8'h55 == _match_key_qbytes_5_T ? phv_data_85 : _GEN_11361; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11363 = 8'h56 == _match_key_qbytes_5_T ? phv_data_86 : _GEN_11362; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11364 = 8'h57 == _match_key_qbytes_5_T ? phv_data_87 : _GEN_11363; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11365 = 8'h58 == _match_key_qbytes_5_T ? phv_data_88 : _GEN_11364; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11366 = 8'h59 == _match_key_qbytes_5_T ? phv_data_89 : _GEN_11365; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11367 = 8'h5a == _match_key_qbytes_5_T ? phv_data_90 : _GEN_11366; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11368 = 8'h5b == _match_key_qbytes_5_T ? phv_data_91 : _GEN_11367; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11369 = 8'h5c == _match_key_qbytes_5_T ? phv_data_92 : _GEN_11368; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11370 = 8'h5d == _match_key_qbytes_5_T ? phv_data_93 : _GEN_11369; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11371 = 8'h5e == _match_key_qbytes_5_T ? phv_data_94 : _GEN_11370; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11372 = 8'h5f == _match_key_qbytes_5_T ? phv_data_95 : _GEN_11371; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11373 = 8'h60 == _match_key_qbytes_5_T ? phv_data_96 : _GEN_11372; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11374 = 8'h61 == _match_key_qbytes_5_T ? phv_data_97 : _GEN_11373; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11375 = 8'h62 == _match_key_qbytes_5_T ? phv_data_98 : _GEN_11374; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11376 = 8'h63 == _match_key_qbytes_5_T ? phv_data_99 : _GEN_11375; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11377 = 8'h64 == _match_key_qbytes_5_T ? phv_data_100 : _GEN_11376; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11378 = 8'h65 == _match_key_qbytes_5_T ? phv_data_101 : _GEN_11377; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11379 = 8'h66 == _match_key_qbytes_5_T ? phv_data_102 : _GEN_11378; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11380 = 8'h67 == _match_key_qbytes_5_T ? phv_data_103 : _GEN_11379; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11381 = 8'h68 == _match_key_qbytes_5_T ? phv_data_104 : _GEN_11380; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11382 = 8'h69 == _match_key_qbytes_5_T ? phv_data_105 : _GEN_11381; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11383 = 8'h6a == _match_key_qbytes_5_T ? phv_data_106 : _GEN_11382; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11384 = 8'h6b == _match_key_qbytes_5_T ? phv_data_107 : _GEN_11383; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11385 = 8'h6c == _match_key_qbytes_5_T ? phv_data_108 : _GEN_11384; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11386 = 8'h6d == _match_key_qbytes_5_T ? phv_data_109 : _GEN_11385; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11387 = 8'h6e == _match_key_qbytes_5_T ? phv_data_110 : _GEN_11386; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11388 = 8'h6f == _match_key_qbytes_5_T ? phv_data_111 : _GEN_11387; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11389 = 8'h70 == _match_key_qbytes_5_T ? phv_data_112 : _GEN_11388; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11390 = 8'h71 == _match_key_qbytes_5_T ? phv_data_113 : _GEN_11389; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11391 = 8'h72 == _match_key_qbytes_5_T ? phv_data_114 : _GEN_11390; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11392 = 8'h73 == _match_key_qbytes_5_T ? phv_data_115 : _GEN_11391; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11393 = 8'h74 == _match_key_qbytes_5_T ? phv_data_116 : _GEN_11392; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11394 = 8'h75 == _match_key_qbytes_5_T ? phv_data_117 : _GEN_11393; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11395 = 8'h76 == _match_key_qbytes_5_T ? phv_data_118 : _GEN_11394; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11396 = 8'h77 == _match_key_qbytes_5_T ? phv_data_119 : _GEN_11395; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11397 = 8'h78 == _match_key_qbytes_5_T ? phv_data_120 : _GEN_11396; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11398 = 8'h79 == _match_key_qbytes_5_T ? phv_data_121 : _GEN_11397; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11399 = 8'h7a == _match_key_qbytes_5_T ? phv_data_122 : _GEN_11398; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11400 = 8'h7b == _match_key_qbytes_5_T ? phv_data_123 : _GEN_11399; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11401 = 8'h7c == _match_key_qbytes_5_T ? phv_data_124 : _GEN_11400; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11402 = 8'h7d == _match_key_qbytes_5_T ? phv_data_125 : _GEN_11401; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11403 = 8'h7e == _match_key_qbytes_5_T ? phv_data_126 : _GEN_11402; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11404 = 8'h7f == _match_key_qbytes_5_T ? phv_data_127 : _GEN_11403; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11405 = 8'h80 == _match_key_qbytes_5_T ? phv_data_128 : _GEN_11404; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11406 = 8'h81 == _match_key_qbytes_5_T ? phv_data_129 : _GEN_11405; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11407 = 8'h82 == _match_key_qbytes_5_T ? phv_data_130 : _GEN_11406; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11408 = 8'h83 == _match_key_qbytes_5_T ? phv_data_131 : _GEN_11407; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11409 = 8'h84 == _match_key_qbytes_5_T ? phv_data_132 : _GEN_11408; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11410 = 8'h85 == _match_key_qbytes_5_T ? phv_data_133 : _GEN_11409; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11411 = 8'h86 == _match_key_qbytes_5_T ? phv_data_134 : _GEN_11410; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11412 = 8'h87 == _match_key_qbytes_5_T ? phv_data_135 : _GEN_11411; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11413 = 8'h88 == _match_key_qbytes_5_T ? phv_data_136 : _GEN_11412; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11414 = 8'h89 == _match_key_qbytes_5_T ? phv_data_137 : _GEN_11413; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11415 = 8'h8a == _match_key_qbytes_5_T ? phv_data_138 : _GEN_11414; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11416 = 8'h8b == _match_key_qbytes_5_T ? phv_data_139 : _GEN_11415; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11417 = 8'h8c == _match_key_qbytes_5_T ? phv_data_140 : _GEN_11416; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11418 = 8'h8d == _match_key_qbytes_5_T ? phv_data_141 : _GEN_11417; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11419 = 8'h8e == _match_key_qbytes_5_T ? phv_data_142 : _GEN_11418; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11420 = 8'h8f == _match_key_qbytes_5_T ? phv_data_143 : _GEN_11419; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11421 = 8'h90 == _match_key_qbytes_5_T ? phv_data_144 : _GEN_11420; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11422 = 8'h91 == _match_key_qbytes_5_T ? phv_data_145 : _GEN_11421; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11423 = 8'h92 == _match_key_qbytes_5_T ? phv_data_146 : _GEN_11422; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11424 = 8'h93 == _match_key_qbytes_5_T ? phv_data_147 : _GEN_11423; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11425 = 8'h94 == _match_key_qbytes_5_T ? phv_data_148 : _GEN_11424; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11426 = 8'h95 == _match_key_qbytes_5_T ? phv_data_149 : _GEN_11425; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11427 = 8'h96 == _match_key_qbytes_5_T ? phv_data_150 : _GEN_11426; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11428 = 8'h97 == _match_key_qbytes_5_T ? phv_data_151 : _GEN_11427; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11429 = 8'h98 == _match_key_qbytes_5_T ? phv_data_152 : _GEN_11428; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11430 = 8'h99 == _match_key_qbytes_5_T ? phv_data_153 : _GEN_11429; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11431 = 8'h9a == _match_key_qbytes_5_T ? phv_data_154 : _GEN_11430; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11432 = 8'h9b == _match_key_qbytes_5_T ? phv_data_155 : _GEN_11431; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11433 = 8'h9c == _match_key_qbytes_5_T ? phv_data_156 : _GEN_11432; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11434 = 8'h9d == _match_key_qbytes_5_T ? phv_data_157 : _GEN_11433; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11435 = 8'h9e == _match_key_qbytes_5_T ? phv_data_158 : _GEN_11434; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11436 = 8'h9f == _match_key_qbytes_5_T ? phv_data_159 : _GEN_11435; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11437 = 8'ha0 == _match_key_qbytes_5_T ? phv_data_160 : _GEN_11436; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11438 = 8'ha1 == _match_key_qbytes_5_T ? phv_data_161 : _GEN_11437; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11439 = 8'ha2 == _match_key_qbytes_5_T ? phv_data_162 : _GEN_11438; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11440 = 8'ha3 == _match_key_qbytes_5_T ? phv_data_163 : _GEN_11439; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11441 = 8'ha4 == _match_key_qbytes_5_T ? phv_data_164 : _GEN_11440; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11442 = 8'ha5 == _match_key_qbytes_5_T ? phv_data_165 : _GEN_11441; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11443 = 8'ha6 == _match_key_qbytes_5_T ? phv_data_166 : _GEN_11442; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11444 = 8'ha7 == _match_key_qbytes_5_T ? phv_data_167 : _GEN_11443; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11445 = 8'ha8 == _match_key_qbytes_5_T ? phv_data_168 : _GEN_11444; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11446 = 8'ha9 == _match_key_qbytes_5_T ? phv_data_169 : _GEN_11445; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11447 = 8'haa == _match_key_qbytes_5_T ? phv_data_170 : _GEN_11446; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11448 = 8'hab == _match_key_qbytes_5_T ? phv_data_171 : _GEN_11447; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11449 = 8'hac == _match_key_qbytes_5_T ? phv_data_172 : _GEN_11448; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11450 = 8'had == _match_key_qbytes_5_T ? phv_data_173 : _GEN_11449; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11451 = 8'hae == _match_key_qbytes_5_T ? phv_data_174 : _GEN_11450; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11452 = 8'haf == _match_key_qbytes_5_T ? phv_data_175 : _GEN_11451; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11453 = 8'hb0 == _match_key_qbytes_5_T ? phv_data_176 : _GEN_11452; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11454 = 8'hb1 == _match_key_qbytes_5_T ? phv_data_177 : _GEN_11453; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11455 = 8'hb2 == _match_key_qbytes_5_T ? phv_data_178 : _GEN_11454; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11456 = 8'hb3 == _match_key_qbytes_5_T ? phv_data_179 : _GEN_11455; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11457 = 8'hb4 == _match_key_qbytes_5_T ? phv_data_180 : _GEN_11456; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11458 = 8'hb5 == _match_key_qbytes_5_T ? phv_data_181 : _GEN_11457; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11459 = 8'hb6 == _match_key_qbytes_5_T ? phv_data_182 : _GEN_11458; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11460 = 8'hb7 == _match_key_qbytes_5_T ? phv_data_183 : _GEN_11459; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11461 = 8'hb8 == _match_key_qbytes_5_T ? phv_data_184 : _GEN_11460; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11462 = 8'hb9 == _match_key_qbytes_5_T ? phv_data_185 : _GEN_11461; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11463 = 8'hba == _match_key_qbytes_5_T ? phv_data_186 : _GEN_11462; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11464 = 8'hbb == _match_key_qbytes_5_T ? phv_data_187 : _GEN_11463; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11465 = 8'hbc == _match_key_qbytes_5_T ? phv_data_188 : _GEN_11464; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11466 = 8'hbd == _match_key_qbytes_5_T ? phv_data_189 : _GEN_11465; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11467 = 8'hbe == _match_key_qbytes_5_T ? phv_data_190 : _GEN_11466; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11468 = 8'hbf == _match_key_qbytes_5_T ? phv_data_191 : _GEN_11467; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11469 = 8'hc0 == _match_key_qbytes_5_T ? phv_data_192 : _GEN_11468; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11470 = 8'hc1 == _match_key_qbytes_5_T ? phv_data_193 : _GEN_11469; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11471 = 8'hc2 == _match_key_qbytes_5_T ? phv_data_194 : _GEN_11470; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11472 = 8'hc3 == _match_key_qbytes_5_T ? phv_data_195 : _GEN_11471; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11473 = 8'hc4 == _match_key_qbytes_5_T ? phv_data_196 : _GEN_11472; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11474 = 8'hc5 == _match_key_qbytes_5_T ? phv_data_197 : _GEN_11473; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11475 = 8'hc6 == _match_key_qbytes_5_T ? phv_data_198 : _GEN_11474; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11476 = 8'hc7 == _match_key_qbytes_5_T ? phv_data_199 : _GEN_11475; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11477 = 8'hc8 == _match_key_qbytes_5_T ? phv_data_200 : _GEN_11476; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11478 = 8'hc9 == _match_key_qbytes_5_T ? phv_data_201 : _GEN_11477; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11479 = 8'hca == _match_key_qbytes_5_T ? phv_data_202 : _GEN_11478; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11480 = 8'hcb == _match_key_qbytes_5_T ? phv_data_203 : _GEN_11479; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11481 = 8'hcc == _match_key_qbytes_5_T ? phv_data_204 : _GEN_11480; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11482 = 8'hcd == _match_key_qbytes_5_T ? phv_data_205 : _GEN_11481; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11483 = 8'hce == _match_key_qbytes_5_T ? phv_data_206 : _GEN_11482; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11484 = 8'hcf == _match_key_qbytes_5_T ? phv_data_207 : _GEN_11483; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11485 = 8'hd0 == _match_key_qbytes_5_T ? phv_data_208 : _GEN_11484; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11486 = 8'hd1 == _match_key_qbytes_5_T ? phv_data_209 : _GEN_11485; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11487 = 8'hd2 == _match_key_qbytes_5_T ? phv_data_210 : _GEN_11486; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11488 = 8'hd3 == _match_key_qbytes_5_T ? phv_data_211 : _GEN_11487; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11489 = 8'hd4 == _match_key_qbytes_5_T ? phv_data_212 : _GEN_11488; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11490 = 8'hd5 == _match_key_qbytes_5_T ? phv_data_213 : _GEN_11489; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11491 = 8'hd6 == _match_key_qbytes_5_T ? phv_data_214 : _GEN_11490; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11492 = 8'hd7 == _match_key_qbytes_5_T ? phv_data_215 : _GEN_11491; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11493 = 8'hd8 == _match_key_qbytes_5_T ? phv_data_216 : _GEN_11492; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11494 = 8'hd9 == _match_key_qbytes_5_T ? phv_data_217 : _GEN_11493; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11495 = 8'hda == _match_key_qbytes_5_T ? phv_data_218 : _GEN_11494; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11496 = 8'hdb == _match_key_qbytes_5_T ? phv_data_219 : _GEN_11495; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11497 = 8'hdc == _match_key_qbytes_5_T ? phv_data_220 : _GEN_11496; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11498 = 8'hdd == _match_key_qbytes_5_T ? phv_data_221 : _GEN_11497; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11499 = 8'hde == _match_key_qbytes_5_T ? phv_data_222 : _GEN_11498; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11500 = 8'hdf == _match_key_qbytes_5_T ? phv_data_223 : _GEN_11499; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11501 = 8'he0 == _match_key_qbytes_5_T ? phv_data_224 : _GEN_11500; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11502 = 8'he1 == _match_key_qbytes_5_T ? phv_data_225 : _GEN_11501; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11503 = 8'he2 == _match_key_qbytes_5_T ? phv_data_226 : _GEN_11502; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11504 = 8'he3 == _match_key_qbytes_5_T ? phv_data_227 : _GEN_11503; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11505 = 8'he4 == _match_key_qbytes_5_T ? phv_data_228 : _GEN_11504; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11506 = 8'he5 == _match_key_qbytes_5_T ? phv_data_229 : _GEN_11505; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11507 = 8'he6 == _match_key_qbytes_5_T ? phv_data_230 : _GEN_11506; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11508 = 8'he7 == _match_key_qbytes_5_T ? phv_data_231 : _GEN_11507; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11509 = 8'he8 == _match_key_qbytes_5_T ? phv_data_232 : _GEN_11508; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11510 = 8'he9 == _match_key_qbytes_5_T ? phv_data_233 : _GEN_11509; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11511 = 8'hea == _match_key_qbytes_5_T ? phv_data_234 : _GEN_11510; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11512 = 8'heb == _match_key_qbytes_5_T ? phv_data_235 : _GEN_11511; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11513 = 8'hec == _match_key_qbytes_5_T ? phv_data_236 : _GEN_11512; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11514 = 8'hed == _match_key_qbytes_5_T ? phv_data_237 : _GEN_11513; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11515 = 8'hee == _match_key_qbytes_5_T ? phv_data_238 : _GEN_11514; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11516 = 8'hef == _match_key_qbytes_5_T ? phv_data_239 : _GEN_11515; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11517 = 8'hf0 == _match_key_qbytes_5_T ? phv_data_240 : _GEN_11516; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11518 = 8'hf1 == _match_key_qbytes_5_T ? phv_data_241 : _GEN_11517; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11519 = 8'hf2 == _match_key_qbytes_5_T ? phv_data_242 : _GEN_11518; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11520 = 8'hf3 == _match_key_qbytes_5_T ? phv_data_243 : _GEN_11519; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11521 = 8'hf4 == _match_key_qbytes_5_T ? phv_data_244 : _GEN_11520; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11522 = 8'hf5 == _match_key_qbytes_5_T ? phv_data_245 : _GEN_11521; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11523 = 8'hf6 == _match_key_qbytes_5_T ? phv_data_246 : _GEN_11522; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11524 = 8'hf7 == _match_key_qbytes_5_T ? phv_data_247 : _GEN_11523; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11525 = 8'hf8 == _match_key_qbytes_5_T ? phv_data_248 : _GEN_11524; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11526 = 8'hf9 == _match_key_qbytes_5_T ? phv_data_249 : _GEN_11525; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11527 = 8'hfa == _match_key_qbytes_5_T ? phv_data_250 : _GEN_11526; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11528 = 8'hfb == _match_key_qbytes_5_T ? phv_data_251 : _GEN_11527; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11529 = 8'hfc == _match_key_qbytes_5_T ? phv_data_252 : _GEN_11528; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11530 = 8'hfd == _match_key_qbytes_5_T ? phv_data_253 : _GEN_11529; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11531 = 8'hfe == _match_key_qbytes_5_T ? phv_data_254 : _GEN_11530; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11532 = 8'hff == _match_key_qbytes_5_T ? phv_data_255 : _GEN_11531; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_17958 = {{1'd0}, _match_key_qbytes_5_T}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11533 = 9'h100 == _GEN_17958 ? phv_data_256 : _GEN_11532; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11534 = 9'h101 == _GEN_17958 ? phv_data_257 : _GEN_11533; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11535 = 9'h102 == _GEN_17958 ? phv_data_258 : _GEN_11534; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11536 = 9'h103 == _GEN_17958 ? phv_data_259 : _GEN_11535; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11537 = 9'h104 == _GEN_17958 ? phv_data_260 : _GEN_11536; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11538 = 9'h105 == _GEN_17958 ? phv_data_261 : _GEN_11537; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11539 = 9'h106 == _GEN_17958 ? phv_data_262 : _GEN_11538; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11540 = 9'h107 == _GEN_17958 ? phv_data_263 : _GEN_11539; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11541 = 9'h108 == _GEN_17958 ? phv_data_264 : _GEN_11540; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11542 = 9'h109 == _GEN_17958 ? phv_data_265 : _GEN_11541; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11543 = 9'h10a == _GEN_17958 ? phv_data_266 : _GEN_11542; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11544 = 9'h10b == _GEN_17958 ? phv_data_267 : _GEN_11543; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11545 = 9'h10c == _GEN_17958 ? phv_data_268 : _GEN_11544; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11546 = 9'h10d == _GEN_17958 ? phv_data_269 : _GEN_11545; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11547 = 9'h10e == _GEN_17958 ? phv_data_270 : _GEN_11546; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11548 = 9'h10f == _GEN_17958 ? phv_data_271 : _GEN_11547; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11549 = 9'h110 == _GEN_17958 ? phv_data_272 : _GEN_11548; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11550 = 9'h111 == _GEN_17958 ? phv_data_273 : _GEN_11549; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11551 = 9'h112 == _GEN_17958 ? phv_data_274 : _GEN_11550; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11552 = 9'h113 == _GEN_17958 ? phv_data_275 : _GEN_11551; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11553 = 9'h114 == _GEN_17958 ? phv_data_276 : _GEN_11552; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11554 = 9'h115 == _GEN_17958 ? phv_data_277 : _GEN_11553; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11555 = 9'h116 == _GEN_17958 ? phv_data_278 : _GEN_11554; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11556 = 9'h117 == _GEN_17958 ? phv_data_279 : _GEN_11555; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11557 = 9'h118 == _GEN_17958 ? phv_data_280 : _GEN_11556; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11558 = 9'h119 == _GEN_17958 ? phv_data_281 : _GEN_11557; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11559 = 9'h11a == _GEN_17958 ? phv_data_282 : _GEN_11558; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11560 = 9'h11b == _GEN_17958 ? phv_data_283 : _GEN_11559; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11561 = 9'h11c == _GEN_17958 ? phv_data_284 : _GEN_11560; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11562 = 9'h11d == _GEN_17958 ? phv_data_285 : _GEN_11561; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11563 = 9'h11e == _GEN_17958 ? phv_data_286 : _GEN_11562; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11564 = 9'h11f == _GEN_17958 ? phv_data_287 : _GEN_11563; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11565 = 9'h120 == _GEN_17958 ? phv_data_288 : _GEN_11564; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11566 = 9'h121 == _GEN_17958 ? phv_data_289 : _GEN_11565; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11567 = 9'h122 == _GEN_17958 ? phv_data_290 : _GEN_11566; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11568 = 9'h123 == _GEN_17958 ? phv_data_291 : _GEN_11567; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11569 = 9'h124 == _GEN_17958 ? phv_data_292 : _GEN_11568; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11570 = 9'h125 == _GEN_17958 ? phv_data_293 : _GEN_11569; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11571 = 9'h126 == _GEN_17958 ? phv_data_294 : _GEN_11570; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11572 = 9'h127 == _GEN_17958 ? phv_data_295 : _GEN_11571; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11573 = 9'h128 == _GEN_17958 ? phv_data_296 : _GEN_11572; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11574 = 9'h129 == _GEN_17958 ? phv_data_297 : _GEN_11573; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11575 = 9'h12a == _GEN_17958 ? phv_data_298 : _GEN_11574; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11576 = 9'h12b == _GEN_17958 ? phv_data_299 : _GEN_11575; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11577 = 9'h12c == _GEN_17958 ? phv_data_300 : _GEN_11576; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11578 = 9'h12d == _GEN_17958 ? phv_data_301 : _GEN_11577; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11579 = 9'h12e == _GEN_17958 ? phv_data_302 : _GEN_11578; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11580 = 9'h12f == _GEN_17958 ? phv_data_303 : _GEN_11579; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11581 = 9'h130 == _GEN_17958 ? phv_data_304 : _GEN_11580; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11582 = 9'h131 == _GEN_17958 ? phv_data_305 : _GEN_11581; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11583 = 9'h132 == _GEN_17958 ? phv_data_306 : _GEN_11582; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11584 = 9'h133 == _GEN_17958 ? phv_data_307 : _GEN_11583; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11585 = 9'h134 == _GEN_17958 ? phv_data_308 : _GEN_11584; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11586 = 9'h135 == _GEN_17958 ? phv_data_309 : _GEN_11585; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11587 = 9'h136 == _GEN_17958 ? phv_data_310 : _GEN_11586; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11588 = 9'h137 == _GEN_17958 ? phv_data_311 : _GEN_11587; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11589 = 9'h138 == _GEN_17958 ? phv_data_312 : _GEN_11588; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11590 = 9'h139 == _GEN_17958 ? phv_data_313 : _GEN_11589; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11591 = 9'h13a == _GEN_17958 ? phv_data_314 : _GEN_11590; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11592 = 9'h13b == _GEN_17958 ? phv_data_315 : _GEN_11591; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11593 = 9'h13c == _GEN_17958 ? phv_data_316 : _GEN_11592; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11594 = 9'h13d == _GEN_17958 ? phv_data_317 : _GEN_11593; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11595 = 9'h13e == _GEN_17958 ? phv_data_318 : _GEN_11594; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11596 = 9'h13f == _GEN_17958 ? phv_data_319 : _GEN_11595; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11597 = 9'h140 == _GEN_17958 ? phv_data_320 : _GEN_11596; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11598 = 9'h141 == _GEN_17958 ? phv_data_321 : _GEN_11597; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11599 = 9'h142 == _GEN_17958 ? phv_data_322 : _GEN_11598; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11600 = 9'h143 == _GEN_17958 ? phv_data_323 : _GEN_11599; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11601 = 9'h144 == _GEN_17958 ? phv_data_324 : _GEN_11600; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11602 = 9'h145 == _GEN_17958 ? phv_data_325 : _GEN_11601; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11603 = 9'h146 == _GEN_17958 ? phv_data_326 : _GEN_11602; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11604 = 9'h147 == _GEN_17958 ? phv_data_327 : _GEN_11603; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11605 = 9'h148 == _GEN_17958 ? phv_data_328 : _GEN_11604; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11606 = 9'h149 == _GEN_17958 ? phv_data_329 : _GEN_11605; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11607 = 9'h14a == _GEN_17958 ? phv_data_330 : _GEN_11606; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11608 = 9'h14b == _GEN_17958 ? phv_data_331 : _GEN_11607; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11609 = 9'h14c == _GEN_17958 ? phv_data_332 : _GEN_11608; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11610 = 9'h14d == _GEN_17958 ? phv_data_333 : _GEN_11609; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11611 = 9'h14e == _GEN_17958 ? phv_data_334 : _GEN_11610; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11612 = 9'h14f == _GEN_17958 ? phv_data_335 : _GEN_11611; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11613 = 9'h150 == _GEN_17958 ? phv_data_336 : _GEN_11612; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11614 = 9'h151 == _GEN_17958 ? phv_data_337 : _GEN_11613; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11615 = 9'h152 == _GEN_17958 ? phv_data_338 : _GEN_11614; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11616 = 9'h153 == _GEN_17958 ? phv_data_339 : _GEN_11615; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11617 = 9'h154 == _GEN_17958 ? phv_data_340 : _GEN_11616; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11618 = 9'h155 == _GEN_17958 ? phv_data_341 : _GEN_11617; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11619 = 9'h156 == _GEN_17958 ? phv_data_342 : _GEN_11618; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11620 = 9'h157 == _GEN_17958 ? phv_data_343 : _GEN_11619; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11621 = 9'h158 == _GEN_17958 ? phv_data_344 : _GEN_11620; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11622 = 9'h159 == _GEN_17958 ? phv_data_345 : _GEN_11621; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11623 = 9'h15a == _GEN_17958 ? phv_data_346 : _GEN_11622; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11624 = 9'h15b == _GEN_17958 ? phv_data_347 : _GEN_11623; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11625 = 9'h15c == _GEN_17958 ? phv_data_348 : _GEN_11624; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11626 = 9'h15d == _GEN_17958 ? phv_data_349 : _GEN_11625; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11627 = 9'h15e == _GEN_17958 ? phv_data_350 : _GEN_11626; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11628 = 9'h15f == _GEN_17958 ? phv_data_351 : _GEN_11627; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11629 = 9'h160 == _GEN_17958 ? phv_data_352 : _GEN_11628; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11630 = 9'h161 == _GEN_17958 ? phv_data_353 : _GEN_11629; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11631 = 9'h162 == _GEN_17958 ? phv_data_354 : _GEN_11630; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11632 = 9'h163 == _GEN_17958 ? phv_data_355 : _GEN_11631; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11633 = 9'h164 == _GEN_17958 ? phv_data_356 : _GEN_11632; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11634 = 9'h165 == _GEN_17958 ? phv_data_357 : _GEN_11633; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11635 = 9'h166 == _GEN_17958 ? phv_data_358 : _GEN_11634; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11636 = 9'h167 == _GEN_17958 ? phv_data_359 : _GEN_11635; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11637 = 9'h168 == _GEN_17958 ? phv_data_360 : _GEN_11636; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11638 = 9'h169 == _GEN_17958 ? phv_data_361 : _GEN_11637; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11639 = 9'h16a == _GEN_17958 ? phv_data_362 : _GEN_11638; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11640 = 9'h16b == _GEN_17958 ? phv_data_363 : _GEN_11639; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11641 = 9'h16c == _GEN_17958 ? phv_data_364 : _GEN_11640; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11642 = 9'h16d == _GEN_17958 ? phv_data_365 : _GEN_11641; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11643 = 9'h16e == _GEN_17958 ? phv_data_366 : _GEN_11642; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11644 = 9'h16f == _GEN_17958 ? phv_data_367 : _GEN_11643; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11645 = 9'h170 == _GEN_17958 ? phv_data_368 : _GEN_11644; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11646 = 9'h171 == _GEN_17958 ? phv_data_369 : _GEN_11645; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11647 = 9'h172 == _GEN_17958 ? phv_data_370 : _GEN_11646; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11648 = 9'h173 == _GEN_17958 ? phv_data_371 : _GEN_11647; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11649 = 9'h174 == _GEN_17958 ? phv_data_372 : _GEN_11648; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11650 = 9'h175 == _GEN_17958 ? phv_data_373 : _GEN_11649; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11651 = 9'h176 == _GEN_17958 ? phv_data_374 : _GEN_11650; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11652 = 9'h177 == _GEN_17958 ? phv_data_375 : _GEN_11651; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11653 = 9'h178 == _GEN_17958 ? phv_data_376 : _GEN_11652; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11654 = 9'h179 == _GEN_17958 ? phv_data_377 : _GEN_11653; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11655 = 9'h17a == _GEN_17958 ? phv_data_378 : _GEN_11654; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11656 = 9'h17b == _GEN_17958 ? phv_data_379 : _GEN_11655; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11657 = 9'h17c == _GEN_17958 ? phv_data_380 : _GEN_11656; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11658 = 9'h17d == _GEN_17958 ? phv_data_381 : _GEN_11657; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11659 = 9'h17e == _GEN_17958 ? phv_data_382 : _GEN_11658; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11660 = 9'h17f == _GEN_17958 ? phv_data_383 : _GEN_11659; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11661 = 9'h180 == _GEN_17958 ? phv_data_384 : _GEN_11660; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11662 = 9'h181 == _GEN_17958 ? phv_data_385 : _GEN_11661; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11663 = 9'h182 == _GEN_17958 ? phv_data_386 : _GEN_11662; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11664 = 9'h183 == _GEN_17958 ? phv_data_387 : _GEN_11663; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11665 = 9'h184 == _GEN_17958 ? phv_data_388 : _GEN_11664; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11666 = 9'h185 == _GEN_17958 ? phv_data_389 : _GEN_11665; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11667 = 9'h186 == _GEN_17958 ? phv_data_390 : _GEN_11666; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11668 = 9'h187 == _GEN_17958 ? phv_data_391 : _GEN_11667; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11669 = 9'h188 == _GEN_17958 ? phv_data_392 : _GEN_11668; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11670 = 9'h189 == _GEN_17958 ? phv_data_393 : _GEN_11669; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11671 = 9'h18a == _GEN_17958 ? phv_data_394 : _GEN_11670; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11672 = 9'h18b == _GEN_17958 ? phv_data_395 : _GEN_11671; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11673 = 9'h18c == _GEN_17958 ? phv_data_396 : _GEN_11672; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11674 = 9'h18d == _GEN_17958 ? phv_data_397 : _GEN_11673; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11675 = 9'h18e == _GEN_17958 ? phv_data_398 : _GEN_11674; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11676 = 9'h18f == _GEN_17958 ? phv_data_399 : _GEN_11675; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11677 = 9'h190 == _GEN_17958 ? phv_data_400 : _GEN_11676; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11678 = 9'h191 == _GEN_17958 ? phv_data_401 : _GEN_11677; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11679 = 9'h192 == _GEN_17958 ? phv_data_402 : _GEN_11678; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11680 = 9'h193 == _GEN_17958 ? phv_data_403 : _GEN_11679; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11681 = 9'h194 == _GEN_17958 ? phv_data_404 : _GEN_11680; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11682 = 9'h195 == _GEN_17958 ? phv_data_405 : _GEN_11681; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11683 = 9'h196 == _GEN_17958 ? phv_data_406 : _GEN_11682; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11684 = 9'h197 == _GEN_17958 ? phv_data_407 : _GEN_11683; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11685 = 9'h198 == _GEN_17958 ? phv_data_408 : _GEN_11684; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11686 = 9'h199 == _GEN_17958 ? phv_data_409 : _GEN_11685; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11687 = 9'h19a == _GEN_17958 ? phv_data_410 : _GEN_11686; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11688 = 9'h19b == _GEN_17958 ? phv_data_411 : _GEN_11687; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11689 = 9'h19c == _GEN_17958 ? phv_data_412 : _GEN_11688; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11690 = 9'h19d == _GEN_17958 ? phv_data_413 : _GEN_11689; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11691 = 9'h19e == _GEN_17958 ? phv_data_414 : _GEN_11690; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11692 = 9'h19f == _GEN_17958 ? phv_data_415 : _GEN_11691; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11693 = 9'h1a0 == _GEN_17958 ? phv_data_416 : _GEN_11692; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11694 = 9'h1a1 == _GEN_17958 ? phv_data_417 : _GEN_11693; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11695 = 9'h1a2 == _GEN_17958 ? phv_data_418 : _GEN_11694; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11696 = 9'h1a3 == _GEN_17958 ? phv_data_419 : _GEN_11695; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11697 = 9'h1a4 == _GEN_17958 ? phv_data_420 : _GEN_11696; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11698 = 9'h1a5 == _GEN_17958 ? phv_data_421 : _GEN_11697; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11699 = 9'h1a6 == _GEN_17958 ? phv_data_422 : _GEN_11698; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11700 = 9'h1a7 == _GEN_17958 ? phv_data_423 : _GEN_11699; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11701 = 9'h1a8 == _GEN_17958 ? phv_data_424 : _GEN_11700; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11702 = 9'h1a9 == _GEN_17958 ? phv_data_425 : _GEN_11701; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11703 = 9'h1aa == _GEN_17958 ? phv_data_426 : _GEN_11702; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11704 = 9'h1ab == _GEN_17958 ? phv_data_427 : _GEN_11703; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11705 = 9'h1ac == _GEN_17958 ? phv_data_428 : _GEN_11704; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11706 = 9'h1ad == _GEN_17958 ? phv_data_429 : _GEN_11705; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11707 = 9'h1ae == _GEN_17958 ? phv_data_430 : _GEN_11706; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11708 = 9'h1af == _GEN_17958 ? phv_data_431 : _GEN_11707; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11709 = 9'h1b0 == _GEN_17958 ? phv_data_432 : _GEN_11708; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11710 = 9'h1b1 == _GEN_17958 ? phv_data_433 : _GEN_11709; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11711 = 9'h1b2 == _GEN_17958 ? phv_data_434 : _GEN_11710; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11712 = 9'h1b3 == _GEN_17958 ? phv_data_435 : _GEN_11711; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11713 = 9'h1b4 == _GEN_17958 ? phv_data_436 : _GEN_11712; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11714 = 9'h1b5 == _GEN_17958 ? phv_data_437 : _GEN_11713; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11715 = 9'h1b6 == _GEN_17958 ? phv_data_438 : _GEN_11714; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11716 = 9'h1b7 == _GEN_17958 ? phv_data_439 : _GEN_11715; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11717 = 9'h1b8 == _GEN_17958 ? phv_data_440 : _GEN_11716; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11718 = 9'h1b9 == _GEN_17958 ? phv_data_441 : _GEN_11717; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11719 = 9'h1ba == _GEN_17958 ? phv_data_442 : _GEN_11718; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11720 = 9'h1bb == _GEN_17958 ? phv_data_443 : _GEN_11719; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11721 = 9'h1bc == _GEN_17958 ? phv_data_444 : _GEN_11720; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11722 = 9'h1bd == _GEN_17958 ? phv_data_445 : _GEN_11721; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11723 = 9'h1be == _GEN_17958 ? phv_data_446 : _GEN_11722; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11724 = 9'h1bf == _GEN_17958 ? phv_data_447 : _GEN_11723; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11725 = 9'h1c0 == _GEN_17958 ? phv_data_448 : _GEN_11724; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11726 = 9'h1c1 == _GEN_17958 ? phv_data_449 : _GEN_11725; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11727 = 9'h1c2 == _GEN_17958 ? phv_data_450 : _GEN_11726; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11728 = 9'h1c3 == _GEN_17958 ? phv_data_451 : _GEN_11727; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11729 = 9'h1c4 == _GEN_17958 ? phv_data_452 : _GEN_11728; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11730 = 9'h1c5 == _GEN_17958 ? phv_data_453 : _GEN_11729; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11731 = 9'h1c6 == _GEN_17958 ? phv_data_454 : _GEN_11730; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11732 = 9'h1c7 == _GEN_17958 ? phv_data_455 : _GEN_11731; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11733 = 9'h1c8 == _GEN_17958 ? phv_data_456 : _GEN_11732; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11734 = 9'h1c9 == _GEN_17958 ? phv_data_457 : _GEN_11733; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11735 = 9'h1ca == _GEN_17958 ? phv_data_458 : _GEN_11734; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11736 = 9'h1cb == _GEN_17958 ? phv_data_459 : _GEN_11735; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11737 = 9'h1cc == _GEN_17958 ? phv_data_460 : _GEN_11736; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11738 = 9'h1cd == _GEN_17958 ? phv_data_461 : _GEN_11737; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11739 = 9'h1ce == _GEN_17958 ? phv_data_462 : _GEN_11738; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11740 = 9'h1cf == _GEN_17958 ? phv_data_463 : _GEN_11739; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11741 = 9'h1d0 == _GEN_17958 ? phv_data_464 : _GEN_11740; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11742 = 9'h1d1 == _GEN_17958 ? phv_data_465 : _GEN_11741; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11743 = 9'h1d2 == _GEN_17958 ? phv_data_466 : _GEN_11742; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11744 = 9'h1d3 == _GEN_17958 ? phv_data_467 : _GEN_11743; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11745 = 9'h1d4 == _GEN_17958 ? phv_data_468 : _GEN_11744; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11746 = 9'h1d5 == _GEN_17958 ? phv_data_469 : _GEN_11745; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11747 = 9'h1d6 == _GEN_17958 ? phv_data_470 : _GEN_11746; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11748 = 9'h1d7 == _GEN_17958 ? phv_data_471 : _GEN_11747; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11749 = 9'h1d8 == _GEN_17958 ? phv_data_472 : _GEN_11748; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11750 = 9'h1d9 == _GEN_17958 ? phv_data_473 : _GEN_11749; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11751 = 9'h1da == _GEN_17958 ? phv_data_474 : _GEN_11750; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11752 = 9'h1db == _GEN_17958 ? phv_data_475 : _GEN_11751; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11753 = 9'h1dc == _GEN_17958 ? phv_data_476 : _GEN_11752; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11754 = 9'h1dd == _GEN_17958 ? phv_data_477 : _GEN_11753; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11755 = 9'h1de == _GEN_17958 ? phv_data_478 : _GEN_11754; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11756 = 9'h1df == _GEN_17958 ? phv_data_479 : _GEN_11755; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11757 = 9'h1e0 == _GEN_17958 ? phv_data_480 : _GEN_11756; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11758 = 9'h1e1 == _GEN_17958 ? phv_data_481 : _GEN_11757; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11759 = 9'h1e2 == _GEN_17958 ? phv_data_482 : _GEN_11758; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11760 = 9'h1e3 == _GEN_17958 ? phv_data_483 : _GEN_11759; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11761 = 9'h1e4 == _GEN_17958 ? phv_data_484 : _GEN_11760; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11762 = 9'h1e5 == _GEN_17958 ? phv_data_485 : _GEN_11761; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11763 = 9'h1e6 == _GEN_17958 ? phv_data_486 : _GEN_11762; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11764 = 9'h1e7 == _GEN_17958 ? phv_data_487 : _GEN_11763; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11765 = 9'h1e8 == _GEN_17958 ? phv_data_488 : _GEN_11764; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11766 = 9'h1e9 == _GEN_17958 ? phv_data_489 : _GEN_11765; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11767 = 9'h1ea == _GEN_17958 ? phv_data_490 : _GEN_11766; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11768 = 9'h1eb == _GEN_17958 ? phv_data_491 : _GEN_11767; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11769 = 9'h1ec == _GEN_17958 ? phv_data_492 : _GEN_11768; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11770 = 9'h1ed == _GEN_17958 ? phv_data_493 : _GEN_11769; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11771 = 9'h1ee == _GEN_17958 ? phv_data_494 : _GEN_11770; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11772 = 9'h1ef == _GEN_17958 ? phv_data_495 : _GEN_11771; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11773 = 9'h1f0 == _GEN_17958 ? phv_data_496 : _GEN_11772; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11774 = 9'h1f1 == _GEN_17958 ? phv_data_497 : _GEN_11773; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11775 = 9'h1f2 == _GEN_17958 ? phv_data_498 : _GEN_11774; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11776 = 9'h1f3 == _GEN_17958 ? phv_data_499 : _GEN_11775; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11777 = 9'h1f4 == _GEN_17958 ? phv_data_500 : _GEN_11776; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11778 = 9'h1f5 == _GEN_17958 ? phv_data_501 : _GEN_11777; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11779 = 9'h1f6 == _GEN_17958 ? phv_data_502 : _GEN_11778; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11780 = 9'h1f7 == _GEN_17958 ? phv_data_503 : _GEN_11779; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11781 = 9'h1f8 == _GEN_17958 ? phv_data_504 : _GEN_11780; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11782 = 9'h1f9 == _GEN_17958 ? phv_data_505 : _GEN_11781; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11783 = 9'h1fa == _GEN_17958 ? phv_data_506 : _GEN_11782; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11784 = 9'h1fb == _GEN_17958 ? phv_data_507 : _GEN_11783; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11785 = 9'h1fc == _GEN_17958 ? phv_data_508 : _GEN_11784; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11786 = 9'h1fd == _GEN_17958 ? phv_data_509 : _GEN_11785; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11787 = 9'h1fe == _GEN_17958 ? phv_data_510 : _GEN_11786; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11788 = 9'h1ff == _GEN_17958 ? phv_data_511 : _GEN_11787; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11790 = 8'h1 == _match_key_qbytes_5_T_1 ? phv_data_1 : phv_data_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11791 = 8'h2 == _match_key_qbytes_5_T_1 ? phv_data_2 : _GEN_11790; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11792 = 8'h3 == _match_key_qbytes_5_T_1 ? phv_data_3 : _GEN_11791; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11793 = 8'h4 == _match_key_qbytes_5_T_1 ? phv_data_4 : _GEN_11792; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11794 = 8'h5 == _match_key_qbytes_5_T_1 ? phv_data_5 : _GEN_11793; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11795 = 8'h6 == _match_key_qbytes_5_T_1 ? phv_data_6 : _GEN_11794; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11796 = 8'h7 == _match_key_qbytes_5_T_1 ? phv_data_7 : _GEN_11795; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11797 = 8'h8 == _match_key_qbytes_5_T_1 ? phv_data_8 : _GEN_11796; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11798 = 8'h9 == _match_key_qbytes_5_T_1 ? phv_data_9 : _GEN_11797; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11799 = 8'ha == _match_key_qbytes_5_T_1 ? phv_data_10 : _GEN_11798; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11800 = 8'hb == _match_key_qbytes_5_T_1 ? phv_data_11 : _GEN_11799; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11801 = 8'hc == _match_key_qbytes_5_T_1 ? phv_data_12 : _GEN_11800; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11802 = 8'hd == _match_key_qbytes_5_T_1 ? phv_data_13 : _GEN_11801; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11803 = 8'he == _match_key_qbytes_5_T_1 ? phv_data_14 : _GEN_11802; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11804 = 8'hf == _match_key_qbytes_5_T_1 ? phv_data_15 : _GEN_11803; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11805 = 8'h10 == _match_key_qbytes_5_T_1 ? phv_data_16 : _GEN_11804; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11806 = 8'h11 == _match_key_qbytes_5_T_1 ? phv_data_17 : _GEN_11805; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11807 = 8'h12 == _match_key_qbytes_5_T_1 ? phv_data_18 : _GEN_11806; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11808 = 8'h13 == _match_key_qbytes_5_T_1 ? phv_data_19 : _GEN_11807; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11809 = 8'h14 == _match_key_qbytes_5_T_1 ? phv_data_20 : _GEN_11808; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11810 = 8'h15 == _match_key_qbytes_5_T_1 ? phv_data_21 : _GEN_11809; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11811 = 8'h16 == _match_key_qbytes_5_T_1 ? phv_data_22 : _GEN_11810; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11812 = 8'h17 == _match_key_qbytes_5_T_1 ? phv_data_23 : _GEN_11811; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11813 = 8'h18 == _match_key_qbytes_5_T_1 ? phv_data_24 : _GEN_11812; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11814 = 8'h19 == _match_key_qbytes_5_T_1 ? phv_data_25 : _GEN_11813; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11815 = 8'h1a == _match_key_qbytes_5_T_1 ? phv_data_26 : _GEN_11814; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11816 = 8'h1b == _match_key_qbytes_5_T_1 ? phv_data_27 : _GEN_11815; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11817 = 8'h1c == _match_key_qbytes_5_T_1 ? phv_data_28 : _GEN_11816; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11818 = 8'h1d == _match_key_qbytes_5_T_1 ? phv_data_29 : _GEN_11817; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11819 = 8'h1e == _match_key_qbytes_5_T_1 ? phv_data_30 : _GEN_11818; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11820 = 8'h1f == _match_key_qbytes_5_T_1 ? phv_data_31 : _GEN_11819; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11821 = 8'h20 == _match_key_qbytes_5_T_1 ? phv_data_32 : _GEN_11820; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11822 = 8'h21 == _match_key_qbytes_5_T_1 ? phv_data_33 : _GEN_11821; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11823 = 8'h22 == _match_key_qbytes_5_T_1 ? phv_data_34 : _GEN_11822; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11824 = 8'h23 == _match_key_qbytes_5_T_1 ? phv_data_35 : _GEN_11823; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11825 = 8'h24 == _match_key_qbytes_5_T_1 ? phv_data_36 : _GEN_11824; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11826 = 8'h25 == _match_key_qbytes_5_T_1 ? phv_data_37 : _GEN_11825; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11827 = 8'h26 == _match_key_qbytes_5_T_1 ? phv_data_38 : _GEN_11826; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11828 = 8'h27 == _match_key_qbytes_5_T_1 ? phv_data_39 : _GEN_11827; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11829 = 8'h28 == _match_key_qbytes_5_T_1 ? phv_data_40 : _GEN_11828; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11830 = 8'h29 == _match_key_qbytes_5_T_1 ? phv_data_41 : _GEN_11829; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11831 = 8'h2a == _match_key_qbytes_5_T_1 ? phv_data_42 : _GEN_11830; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11832 = 8'h2b == _match_key_qbytes_5_T_1 ? phv_data_43 : _GEN_11831; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11833 = 8'h2c == _match_key_qbytes_5_T_1 ? phv_data_44 : _GEN_11832; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11834 = 8'h2d == _match_key_qbytes_5_T_1 ? phv_data_45 : _GEN_11833; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11835 = 8'h2e == _match_key_qbytes_5_T_1 ? phv_data_46 : _GEN_11834; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11836 = 8'h2f == _match_key_qbytes_5_T_1 ? phv_data_47 : _GEN_11835; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11837 = 8'h30 == _match_key_qbytes_5_T_1 ? phv_data_48 : _GEN_11836; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11838 = 8'h31 == _match_key_qbytes_5_T_1 ? phv_data_49 : _GEN_11837; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11839 = 8'h32 == _match_key_qbytes_5_T_1 ? phv_data_50 : _GEN_11838; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11840 = 8'h33 == _match_key_qbytes_5_T_1 ? phv_data_51 : _GEN_11839; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11841 = 8'h34 == _match_key_qbytes_5_T_1 ? phv_data_52 : _GEN_11840; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11842 = 8'h35 == _match_key_qbytes_5_T_1 ? phv_data_53 : _GEN_11841; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11843 = 8'h36 == _match_key_qbytes_5_T_1 ? phv_data_54 : _GEN_11842; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11844 = 8'h37 == _match_key_qbytes_5_T_1 ? phv_data_55 : _GEN_11843; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11845 = 8'h38 == _match_key_qbytes_5_T_1 ? phv_data_56 : _GEN_11844; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11846 = 8'h39 == _match_key_qbytes_5_T_1 ? phv_data_57 : _GEN_11845; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11847 = 8'h3a == _match_key_qbytes_5_T_1 ? phv_data_58 : _GEN_11846; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11848 = 8'h3b == _match_key_qbytes_5_T_1 ? phv_data_59 : _GEN_11847; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11849 = 8'h3c == _match_key_qbytes_5_T_1 ? phv_data_60 : _GEN_11848; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11850 = 8'h3d == _match_key_qbytes_5_T_1 ? phv_data_61 : _GEN_11849; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11851 = 8'h3e == _match_key_qbytes_5_T_1 ? phv_data_62 : _GEN_11850; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11852 = 8'h3f == _match_key_qbytes_5_T_1 ? phv_data_63 : _GEN_11851; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11853 = 8'h40 == _match_key_qbytes_5_T_1 ? phv_data_64 : _GEN_11852; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11854 = 8'h41 == _match_key_qbytes_5_T_1 ? phv_data_65 : _GEN_11853; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11855 = 8'h42 == _match_key_qbytes_5_T_1 ? phv_data_66 : _GEN_11854; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11856 = 8'h43 == _match_key_qbytes_5_T_1 ? phv_data_67 : _GEN_11855; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11857 = 8'h44 == _match_key_qbytes_5_T_1 ? phv_data_68 : _GEN_11856; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11858 = 8'h45 == _match_key_qbytes_5_T_1 ? phv_data_69 : _GEN_11857; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11859 = 8'h46 == _match_key_qbytes_5_T_1 ? phv_data_70 : _GEN_11858; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11860 = 8'h47 == _match_key_qbytes_5_T_1 ? phv_data_71 : _GEN_11859; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11861 = 8'h48 == _match_key_qbytes_5_T_1 ? phv_data_72 : _GEN_11860; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11862 = 8'h49 == _match_key_qbytes_5_T_1 ? phv_data_73 : _GEN_11861; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11863 = 8'h4a == _match_key_qbytes_5_T_1 ? phv_data_74 : _GEN_11862; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11864 = 8'h4b == _match_key_qbytes_5_T_1 ? phv_data_75 : _GEN_11863; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11865 = 8'h4c == _match_key_qbytes_5_T_1 ? phv_data_76 : _GEN_11864; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11866 = 8'h4d == _match_key_qbytes_5_T_1 ? phv_data_77 : _GEN_11865; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11867 = 8'h4e == _match_key_qbytes_5_T_1 ? phv_data_78 : _GEN_11866; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11868 = 8'h4f == _match_key_qbytes_5_T_1 ? phv_data_79 : _GEN_11867; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11869 = 8'h50 == _match_key_qbytes_5_T_1 ? phv_data_80 : _GEN_11868; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11870 = 8'h51 == _match_key_qbytes_5_T_1 ? phv_data_81 : _GEN_11869; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11871 = 8'h52 == _match_key_qbytes_5_T_1 ? phv_data_82 : _GEN_11870; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11872 = 8'h53 == _match_key_qbytes_5_T_1 ? phv_data_83 : _GEN_11871; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11873 = 8'h54 == _match_key_qbytes_5_T_1 ? phv_data_84 : _GEN_11872; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11874 = 8'h55 == _match_key_qbytes_5_T_1 ? phv_data_85 : _GEN_11873; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11875 = 8'h56 == _match_key_qbytes_5_T_1 ? phv_data_86 : _GEN_11874; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11876 = 8'h57 == _match_key_qbytes_5_T_1 ? phv_data_87 : _GEN_11875; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11877 = 8'h58 == _match_key_qbytes_5_T_1 ? phv_data_88 : _GEN_11876; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11878 = 8'h59 == _match_key_qbytes_5_T_1 ? phv_data_89 : _GEN_11877; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11879 = 8'h5a == _match_key_qbytes_5_T_1 ? phv_data_90 : _GEN_11878; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11880 = 8'h5b == _match_key_qbytes_5_T_1 ? phv_data_91 : _GEN_11879; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11881 = 8'h5c == _match_key_qbytes_5_T_1 ? phv_data_92 : _GEN_11880; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11882 = 8'h5d == _match_key_qbytes_5_T_1 ? phv_data_93 : _GEN_11881; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11883 = 8'h5e == _match_key_qbytes_5_T_1 ? phv_data_94 : _GEN_11882; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11884 = 8'h5f == _match_key_qbytes_5_T_1 ? phv_data_95 : _GEN_11883; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11885 = 8'h60 == _match_key_qbytes_5_T_1 ? phv_data_96 : _GEN_11884; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11886 = 8'h61 == _match_key_qbytes_5_T_1 ? phv_data_97 : _GEN_11885; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11887 = 8'h62 == _match_key_qbytes_5_T_1 ? phv_data_98 : _GEN_11886; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11888 = 8'h63 == _match_key_qbytes_5_T_1 ? phv_data_99 : _GEN_11887; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11889 = 8'h64 == _match_key_qbytes_5_T_1 ? phv_data_100 : _GEN_11888; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11890 = 8'h65 == _match_key_qbytes_5_T_1 ? phv_data_101 : _GEN_11889; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11891 = 8'h66 == _match_key_qbytes_5_T_1 ? phv_data_102 : _GEN_11890; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11892 = 8'h67 == _match_key_qbytes_5_T_1 ? phv_data_103 : _GEN_11891; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11893 = 8'h68 == _match_key_qbytes_5_T_1 ? phv_data_104 : _GEN_11892; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11894 = 8'h69 == _match_key_qbytes_5_T_1 ? phv_data_105 : _GEN_11893; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11895 = 8'h6a == _match_key_qbytes_5_T_1 ? phv_data_106 : _GEN_11894; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11896 = 8'h6b == _match_key_qbytes_5_T_1 ? phv_data_107 : _GEN_11895; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11897 = 8'h6c == _match_key_qbytes_5_T_1 ? phv_data_108 : _GEN_11896; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11898 = 8'h6d == _match_key_qbytes_5_T_1 ? phv_data_109 : _GEN_11897; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11899 = 8'h6e == _match_key_qbytes_5_T_1 ? phv_data_110 : _GEN_11898; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11900 = 8'h6f == _match_key_qbytes_5_T_1 ? phv_data_111 : _GEN_11899; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11901 = 8'h70 == _match_key_qbytes_5_T_1 ? phv_data_112 : _GEN_11900; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11902 = 8'h71 == _match_key_qbytes_5_T_1 ? phv_data_113 : _GEN_11901; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11903 = 8'h72 == _match_key_qbytes_5_T_1 ? phv_data_114 : _GEN_11902; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11904 = 8'h73 == _match_key_qbytes_5_T_1 ? phv_data_115 : _GEN_11903; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11905 = 8'h74 == _match_key_qbytes_5_T_1 ? phv_data_116 : _GEN_11904; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11906 = 8'h75 == _match_key_qbytes_5_T_1 ? phv_data_117 : _GEN_11905; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11907 = 8'h76 == _match_key_qbytes_5_T_1 ? phv_data_118 : _GEN_11906; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11908 = 8'h77 == _match_key_qbytes_5_T_1 ? phv_data_119 : _GEN_11907; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11909 = 8'h78 == _match_key_qbytes_5_T_1 ? phv_data_120 : _GEN_11908; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11910 = 8'h79 == _match_key_qbytes_5_T_1 ? phv_data_121 : _GEN_11909; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11911 = 8'h7a == _match_key_qbytes_5_T_1 ? phv_data_122 : _GEN_11910; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11912 = 8'h7b == _match_key_qbytes_5_T_1 ? phv_data_123 : _GEN_11911; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11913 = 8'h7c == _match_key_qbytes_5_T_1 ? phv_data_124 : _GEN_11912; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11914 = 8'h7d == _match_key_qbytes_5_T_1 ? phv_data_125 : _GEN_11913; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11915 = 8'h7e == _match_key_qbytes_5_T_1 ? phv_data_126 : _GEN_11914; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11916 = 8'h7f == _match_key_qbytes_5_T_1 ? phv_data_127 : _GEN_11915; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11917 = 8'h80 == _match_key_qbytes_5_T_1 ? phv_data_128 : _GEN_11916; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11918 = 8'h81 == _match_key_qbytes_5_T_1 ? phv_data_129 : _GEN_11917; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11919 = 8'h82 == _match_key_qbytes_5_T_1 ? phv_data_130 : _GEN_11918; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11920 = 8'h83 == _match_key_qbytes_5_T_1 ? phv_data_131 : _GEN_11919; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11921 = 8'h84 == _match_key_qbytes_5_T_1 ? phv_data_132 : _GEN_11920; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11922 = 8'h85 == _match_key_qbytes_5_T_1 ? phv_data_133 : _GEN_11921; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11923 = 8'h86 == _match_key_qbytes_5_T_1 ? phv_data_134 : _GEN_11922; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11924 = 8'h87 == _match_key_qbytes_5_T_1 ? phv_data_135 : _GEN_11923; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11925 = 8'h88 == _match_key_qbytes_5_T_1 ? phv_data_136 : _GEN_11924; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11926 = 8'h89 == _match_key_qbytes_5_T_1 ? phv_data_137 : _GEN_11925; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11927 = 8'h8a == _match_key_qbytes_5_T_1 ? phv_data_138 : _GEN_11926; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11928 = 8'h8b == _match_key_qbytes_5_T_1 ? phv_data_139 : _GEN_11927; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11929 = 8'h8c == _match_key_qbytes_5_T_1 ? phv_data_140 : _GEN_11928; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11930 = 8'h8d == _match_key_qbytes_5_T_1 ? phv_data_141 : _GEN_11929; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11931 = 8'h8e == _match_key_qbytes_5_T_1 ? phv_data_142 : _GEN_11930; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11932 = 8'h8f == _match_key_qbytes_5_T_1 ? phv_data_143 : _GEN_11931; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11933 = 8'h90 == _match_key_qbytes_5_T_1 ? phv_data_144 : _GEN_11932; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11934 = 8'h91 == _match_key_qbytes_5_T_1 ? phv_data_145 : _GEN_11933; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11935 = 8'h92 == _match_key_qbytes_5_T_1 ? phv_data_146 : _GEN_11934; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11936 = 8'h93 == _match_key_qbytes_5_T_1 ? phv_data_147 : _GEN_11935; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11937 = 8'h94 == _match_key_qbytes_5_T_1 ? phv_data_148 : _GEN_11936; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11938 = 8'h95 == _match_key_qbytes_5_T_1 ? phv_data_149 : _GEN_11937; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11939 = 8'h96 == _match_key_qbytes_5_T_1 ? phv_data_150 : _GEN_11938; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11940 = 8'h97 == _match_key_qbytes_5_T_1 ? phv_data_151 : _GEN_11939; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11941 = 8'h98 == _match_key_qbytes_5_T_1 ? phv_data_152 : _GEN_11940; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11942 = 8'h99 == _match_key_qbytes_5_T_1 ? phv_data_153 : _GEN_11941; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11943 = 8'h9a == _match_key_qbytes_5_T_1 ? phv_data_154 : _GEN_11942; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11944 = 8'h9b == _match_key_qbytes_5_T_1 ? phv_data_155 : _GEN_11943; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11945 = 8'h9c == _match_key_qbytes_5_T_1 ? phv_data_156 : _GEN_11944; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11946 = 8'h9d == _match_key_qbytes_5_T_1 ? phv_data_157 : _GEN_11945; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11947 = 8'h9e == _match_key_qbytes_5_T_1 ? phv_data_158 : _GEN_11946; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11948 = 8'h9f == _match_key_qbytes_5_T_1 ? phv_data_159 : _GEN_11947; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11949 = 8'ha0 == _match_key_qbytes_5_T_1 ? phv_data_160 : _GEN_11948; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11950 = 8'ha1 == _match_key_qbytes_5_T_1 ? phv_data_161 : _GEN_11949; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11951 = 8'ha2 == _match_key_qbytes_5_T_1 ? phv_data_162 : _GEN_11950; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11952 = 8'ha3 == _match_key_qbytes_5_T_1 ? phv_data_163 : _GEN_11951; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11953 = 8'ha4 == _match_key_qbytes_5_T_1 ? phv_data_164 : _GEN_11952; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11954 = 8'ha5 == _match_key_qbytes_5_T_1 ? phv_data_165 : _GEN_11953; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11955 = 8'ha6 == _match_key_qbytes_5_T_1 ? phv_data_166 : _GEN_11954; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11956 = 8'ha7 == _match_key_qbytes_5_T_1 ? phv_data_167 : _GEN_11955; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11957 = 8'ha8 == _match_key_qbytes_5_T_1 ? phv_data_168 : _GEN_11956; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11958 = 8'ha9 == _match_key_qbytes_5_T_1 ? phv_data_169 : _GEN_11957; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11959 = 8'haa == _match_key_qbytes_5_T_1 ? phv_data_170 : _GEN_11958; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11960 = 8'hab == _match_key_qbytes_5_T_1 ? phv_data_171 : _GEN_11959; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11961 = 8'hac == _match_key_qbytes_5_T_1 ? phv_data_172 : _GEN_11960; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11962 = 8'had == _match_key_qbytes_5_T_1 ? phv_data_173 : _GEN_11961; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11963 = 8'hae == _match_key_qbytes_5_T_1 ? phv_data_174 : _GEN_11962; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11964 = 8'haf == _match_key_qbytes_5_T_1 ? phv_data_175 : _GEN_11963; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11965 = 8'hb0 == _match_key_qbytes_5_T_1 ? phv_data_176 : _GEN_11964; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11966 = 8'hb1 == _match_key_qbytes_5_T_1 ? phv_data_177 : _GEN_11965; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11967 = 8'hb2 == _match_key_qbytes_5_T_1 ? phv_data_178 : _GEN_11966; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11968 = 8'hb3 == _match_key_qbytes_5_T_1 ? phv_data_179 : _GEN_11967; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11969 = 8'hb4 == _match_key_qbytes_5_T_1 ? phv_data_180 : _GEN_11968; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11970 = 8'hb5 == _match_key_qbytes_5_T_1 ? phv_data_181 : _GEN_11969; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11971 = 8'hb6 == _match_key_qbytes_5_T_1 ? phv_data_182 : _GEN_11970; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11972 = 8'hb7 == _match_key_qbytes_5_T_1 ? phv_data_183 : _GEN_11971; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11973 = 8'hb8 == _match_key_qbytes_5_T_1 ? phv_data_184 : _GEN_11972; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11974 = 8'hb9 == _match_key_qbytes_5_T_1 ? phv_data_185 : _GEN_11973; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11975 = 8'hba == _match_key_qbytes_5_T_1 ? phv_data_186 : _GEN_11974; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11976 = 8'hbb == _match_key_qbytes_5_T_1 ? phv_data_187 : _GEN_11975; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11977 = 8'hbc == _match_key_qbytes_5_T_1 ? phv_data_188 : _GEN_11976; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11978 = 8'hbd == _match_key_qbytes_5_T_1 ? phv_data_189 : _GEN_11977; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11979 = 8'hbe == _match_key_qbytes_5_T_1 ? phv_data_190 : _GEN_11978; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11980 = 8'hbf == _match_key_qbytes_5_T_1 ? phv_data_191 : _GEN_11979; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11981 = 8'hc0 == _match_key_qbytes_5_T_1 ? phv_data_192 : _GEN_11980; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11982 = 8'hc1 == _match_key_qbytes_5_T_1 ? phv_data_193 : _GEN_11981; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11983 = 8'hc2 == _match_key_qbytes_5_T_1 ? phv_data_194 : _GEN_11982; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11984 = 8'hc3 == _match_key_qbytes_5_T_1 ? phv_data_195 : _GEN_11983; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11985 = 8'hc4 == _match_key_qbytes_5_T_1 ? phv_data_196 : _GEN_11984; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11986 = 8'hc5 == _match_key_qbytes_5_T_1 ? phv_data_197 : _GEN_11985; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11987 = 8'hc6 == _match_key_qbytes_5_T_1 ? phv_data_198 : _GEN_11986; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11988 = 8'hc7 == _match_key_qbytes_5_T_1 ? phv_data_199 : _GEN_11987; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11989 = 8'hc8 == _match_key_qbytes_5_T_1 ? phv_data_200 : _GEN_11988; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11990 = 8'hc9 == _match_key_qbytes_5_T_1 ? phv_data_201 : _GEN_11989; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11991 = 8'hca == _match_key_qbytes_5_T_1 ? phv_data_202 : _GEN_11990; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11992 = 8'hcb == _match_key_qbytes_5_T_1 ? phv_data_203 : _GEN_11991; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11993 = 8'hcc == _match_key_qbytes_5_T_1 ? phv_data_204 : _GEN_11992; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11994 = 8'hcd == _match_key_qbytes_5_T_1 ? phv_data_205 : _GEN_11993; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11995 = 8'hce == _match_key_qbytes_5_T_1 ? phv_data_206 : _GEN_11994; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11996 = 8'hcf == _match_key_qbytes_5_T_1 ? phv_data_207 : _GEN_11995; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11997 = 8'hd0 == _match_key_qbytes_5_T_1 ? phv_data_208 : _GEN_11996; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11998 = 8'hd1 == _match_key_qbytes_5_T_1 ? phv_data_209 : _GEN_11997; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11999 = 8'hd2 == _match_key_qbytes_5_T_1 ? phv_data_210 : _GEN_11998; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12000 = 8'hd3 == _match_key_qbytes_5_T_1 ? phv_data_211 : _GEN_11999; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12001 = 8'hd4 == _match_key_qbytes_5_T_1 ? phv_data_212 : _GEN_12000; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12002 = 8'hd5 == _match_key_qbytes_5_T_1 ? phv_data_213 : _GEN_12001; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12003 = 8'hd6 == _match_key_qbytes_5_T_1 ? phv_data_214 : _GEN_12002; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12004 = 8'hd7 == _match_key_qbytes_5_T_1 ? phv_data_215 : _GEN_12003; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12005 = 8'hd8 == _match_key_qbytes_5_T_1 ? phv_data_216 : _GEN_12004; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12006 = 8'hd9 == _match_key_qbytes_5_T_1 ? phv_data_217 : _GEN_12005; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12007 = 8'hda == _match_key_qbytes_5_T_1 ? phv_data_218 : _GEN_12006; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12008 = 8'hdb == _match_key_qbytes_5_T_1 ? phv_data_219 : _GEN_12007; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12009 = 8'hdc == _match_key_qbytes_5_T_1 ? phv_data_220 : _GEN_12008; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12010 = 8'hdd == _match_key_qbytes_5_T_1 ? phv_data_221 : _GEN_12009; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12011 = 8'hde == _match_key_qbytes_5_T_1 ? phv_data_222 : _GEN_12010; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12012 = 8'hdf == _match_key_qbytes_5_T_1 ? phv_data_223 : _GEN_12011; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12013 = 8'he0 == _match_key_qbytes_5_T_1 ? phv_data_224 : _GEN_12012; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12014 = 8'he1 == _match_key_qbytes_5_T_1 ? phv_data_225 : _GEN_12013; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12015 = 8'he2 == _match_key_qbytes_5_T_1 ? phv_data_226 : _GEN_12014; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12016 = 8'he3 == _match_key_qbytes_5_T_1 ? phv_data_227 : _GEN_12015; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12017 = 8'he4 == _match_key_qbytes_5_T_1 ? phv_data_228 : _GEN_12016; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12018 = 8'he5 == _match_key_qbytes_5_T_1 ? phv_data_229 : _GEN_12017; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12019 = 8'he6 == _match_key_qbytes_5_T_1 ? phv_data_230 : _GEN_12018; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12020 = 8'he7 == _match_key_qbytes_5_T_1 ? phv_data_231 : _GEN_12019; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12021 = 8'he8 == _match_key_qbytes_5_T_1 ? phv_data_232 : _GEN_12020; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12022 = 8'he9 == _match_key_qbytes_5_T_1 ? phv_data_233 : _GEN_12021; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12023 = 8'hea == _match_key_qbytes_5_T_1 ? phv_data_234 : _GEN_12022; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12024 = 8'heb == _match_key_qbytes_5_T_1 ? phv_data_235 : _GEN_12023; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12025 = 8'hec == _match_key_qbytes_5_T_1 ? phv_data_236 : _GEN_12024; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12026 = 8'hed == _match_key_qbytes_5_T_1 ? phv_data_237 : _GEN_12025; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12027 = 8'hee == _match_key_qbytes_5_T_1 ? phv_data_238 : _GEN_12026; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12028 = 8'hef == _match_key_qbytes_5_T_1 ? phv_data_239 : _GEN_12027; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12029 = 8'hf0 == _match_key_qbytes_5_T_1 ? phv_data_240 : _GEN_12028; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12030 = 8'hf1 == _match_key_qbytes_5_T_1 ? phv_data_241 : _GEN_12029; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12031 = 8'hf2 == _match_key_qbytes_5_T_1 ? phv_data_242 : _GEN_12030; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12032 = 8'hf3 == _match_key_qbytes_5_T_1 ? phv_data_243 : _GEN_12031; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12033 = 8'hf4 == _match_key_qbytes_5_T_1 ? phv_data_244 : _GEN_12032; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12034 = 8'hf5 == _match_key_qbytes_5_T_1 ? phv_data_245 : _GEN_12033; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12035 = 8'hf6 == _match_key_qbytes_5_T_1 ? phv_data_246 : _GEN_12034; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12036 = 8'hf7 == _match_key_qbytes_5_T_1 ? phv_data_247 : _GEN_12035; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12037 = 8'hf8 == _match_key_qbytes_5_T_1 ? phv_data_248 : _GEN_12036; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12038 = 8'hf9 == _match_key_qbytes_5_T_1 ? phv_data_249 : _GEN_12037; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12039 = 8'hfa == _match_key_qbytes_5_T_1 ? phv_data_250 : _GEN_12038; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12040 = 8'hfb == _match_key_qbytes_5_T_1 ? phv_data_251 : _GEN_12039; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12041 = 8'hfc == _match_key_qbytes_5_T_1 ? phv_data_252 : _GEN_12040; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12042 = 8'hfd == _match_key_qbytes_5_T_1 ? phv_data_253 : _GEN_12041; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12043 = 8'hfe == _match_key_qbytes_5_T_1 ? phv_data_254 : _GEN_12042; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12044 = 8'hff == _match_key_qbytes_5_T_1 ? phv_data_255 : _GEN_12043; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [8:0] _GEN_18214 = {{1'd0}, _match_key_qbytes_5_T_1}; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12045 = 9'h100 == _GEN_18214 ? phv_data_256 : _GEN_12044; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12046 = 9'h101 == _GEN_18214 ? phv_data_257 : _GEN_12045; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12047 = 9'h102 == _GEN_18214 ? phv_data_258 : _GEN_12046; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12048 = 9'h103 == _GEN_18214 ? phv_data_259 : _GEN_12047; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12049 = 9'h104 == _GEN_18214 ? phv_data_260 : _GEN_12048; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12050 = 9'h105 == _GEN_18214 ? phv_data_261 : _GEN_12049; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12051 = 9'h106 == _GEN_18214 ? phv_data_262 : _GEN_12050; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12052 = 9'h107 == _GEN_18214 ? phv_data_263 : _GEN_12051; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12053 = 9'h108 == _GEN_18214 ? phv_data_264 : _GEN_12052; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12054 = 9'h109 == _GEN_18214 ? phv_data_265 : _GEN_12053; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12055 = 9'h10a == _GEN_18214 ? phv_data_266 : _GEN_12054; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12056 = 9'h10b == _GEN_18214 ? phv_data_267 : _GEN_12055; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12057 = 9'h10c == _GEN_18214 ? phv_data_268 : _GEN_12056; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12058 = 9'h10d == _GEN_18214 ? phv_data_269 : _GEN_12057; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12059 = 9'h10e == _GEN_18214 ? phv_data_270 : _GEN_12058; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12060 = 9'h10f == _GEN_18214 ? phv_data_271 : _GEN_12059; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12061 = 9'h110 == _GEN_18214 ? phv_data_272 : _GEN_12060; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12062 = 9'h111 == _GEN_18214 ? phv_data_273 : _GEN_12061; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12063 = 9'h112 == _GEN_18214 ? phv_data_274 : _GEN_12062; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12064 = 9'h113 == _GEN_18214 ? phv_data_275 : _GEN_12063; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12065 = 9'h114 == _GEN_18214 ? phv_data_276 : _GEN_12064; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12066 = 9'h115 == _GEN_18214 ? phv_data_277 : _GEN_12065; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12067 = 9'h116 == _GEN_18214 ? phv_data_278 : _GEN_12066; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12068 = 9'h117 == _GEN_18214 ? phv_data_279 : _GEN_12067; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12069 = 9'h118 == _GEN_18214 ? phv_data_280 : _GEN_12068; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12070 = 9'h119 == _GEN_18214 ? phv_data_281 : _GEN_12069; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12071 = 9'h11a == _GEN_18214 ? phv_data_282 : _GEN_12070; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12072 = 9'h11b == _GEN_18214 ? phv_data_283 : _GEN_12071; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12073 = 9'h11c == _GEN_18214 ? phv_data_284 : _GEN_12072; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12074 = 9'h11d == _GEN_18214 ? phv_data_285 : _GEN_12073; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12075 = 9'h11e == _GEN_18214 ? phv_data_286 : _GEN_12074; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12076 = 9'h11f == _GEN_18214 ? phv_data_287 : _GEN_12075; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12077 = 9'h120 == _GEN_18214 ? phv_data_288 : _GEN_12076; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12078 = 9'h121 == _GEN_18214 ? phv_data_289 : _GEN_12077; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12079 = 9'h122 == _GEN_18214 ? phv_data_290 : _GEN_12078; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12080 = 9'h123 == _GEN_18214 ? phv_data_291 : _GEN_12079; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12081 = 9'h124 == _GEN_18214 ? phv_data_292 : _GEN_12080; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12082 = 9'h125 == _GEN_18214 ? phv_data_293 : _GEN_12081; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12083 = 9'h126 == _GEN_18214 ? phv_data_294 : _GEN_12082; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12084 = 9'h127 == _GEN_18214 ? phv_data_295 : _GEN_12083; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12085 = 9'h128 == _GEN_18214 ? phv_data_296 : _GEN_12084; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12086 = 9'h129 == _GEN_18214 ? phv_data_297 : _GEN_12085; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12087 = 9'h12a == _GEN_18214 ? phv_data_298 : _GEN_12086; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12088 = 9'h12b == _GEN_18214 ? phv_data_299 : _GEN_12087; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12089 = 9'h12c == _GEN_18214 ? phv_data_300 : _GEN_12088; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12090 = 9'h12d == _GEN_18214 ? phv_data_301 : _GEN_12089; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12091 = 9'h12e == _GEN_18214 ? phv_data_302 : _GEN_12090; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12092 = 9'h12f == _GEN_18214 ? phv_data_303 : _GEN_12091; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12093 = 9'h130 == _GEN_18214 ? phv_data_304 : _GEN_12092; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12094 = 9'h131 == _GEN_18214 ? phv_data_305 : _GEN_12093; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12095 = 9'h132 == _GEN_18214 ? phv_data_306 : _GEN_12094; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12096 = 9'h133 == _GEN_18214 ? phv_data_307 : _GEN_12095; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12097 = 9'h134 == _GEN_18214 ? phv_data_308 : _GEN_12096; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12098 = 9'h135 == _GEN_18214 ? phv_data_309 : _GEN_12097; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12099 = 9'h136 == _GEN_18214 ? phv_data_310 : _GEN_12098; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12100 = 9'h137 == _GEN_18214 ? phv_data_311 : _GEN_12099; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12101 = 9'h138 == _GEN_18214 ? phv_data_312 : _GEN_12100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12102 = 9'h139 == _GEN_18214 ? phv_data_313 : _GEN_12101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12103 = 9'h13a == _GEN_18214 ? phv_data_314 : _GEN_12102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12104 = 9'h13b == _GEN_18214 ? phv_data_315 : _GEN_12103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12105 = 9'h13c == _GEN_18214 ? phv_data_316 : _GEN_12104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12106 = 9'h13d == _GEN_18214 ? phv_data_317 : _GEN_12105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12107 = 9'h13e == _GEN_18214 ? phv_data_318 : _GEN_12106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12108 = 9'h13f == _GEN_18214 ? phv_data_319 : _GEN_12107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12109 = 9'h140 == _GEN_18214 ? phv_data_320 : _GEN_12108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12110 = 9'h141 == _GEN_18214 ? phv_data_321 : _GEN_12109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12111 = 9'h142 == _GEN_18214 ? phv_data_322 : _GEN_12110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12112 = 9'h143 == _GEN_18214 ? phv_data_323 : _GEN_12111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12113 = 9'h144 == _GEN_18214 ? phv_data_324 : _GEN_12112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12114 = 9'h145 == _GEN_18214 ? phv_data_325 : _GEN_12113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12115 = 9'h146 == _GEN_18214 ? phv_data_326 : _GEN_12114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12116 = 9'h147 == _GEN_18214 ? phv_data_327 : _GEN_12115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12117 = 9'h148 == _GEN_18214 ? phv_data_328 : _GEN_12116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12118 = 9'h149 == _GEN_18214 ? phv_data_329 : _GEN_12117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12119 = 9'h14a == _GEN_18214 ? phv_data_330 : _GEN_12118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12120 = 9'h14b == _GEN_18214 ? phv_data_331 : _GEN_12119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12121 = 9'h14c == _GEN_18214 ? phv_data_332 : _GEN_12120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12122 = 9'h14d == _GEN_18214 ? phv_data_333 : _GEN_12121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12123 = 9'h14e == _GEN_18214 ? phv_data_334 : _GEN_12122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12124 = 9'h14f == _GEN_18214 ? phv_data_335 : _GEN_12123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12125 = 9'h150 == _GEN_18214 ? phv_data_336 : _GEN_12124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12126 = 9'h151 == _GEN_18214 ? phv_data_337 : _GEN_12125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12127 = 9'h152 == _GEN_18214 ? phv_data_338 : _GEN_12126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12128 = 9'h153 == _GEN_18214 ? phv_data_339 : _GEN_12127; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12129 = 9'h154 == _GEN_18214 ? phv_data_340 : _GEN_12128; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12130 = 9'h155 == _GEN_18214 ? phv_data_341 : _GEN_12129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12131 = 9'h156 == _GEN_18214 ? phv_data_342 : _GEN_12130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12132 = 9'h157 == _GEN_18214 ? phv_data_343 : _GEN_12131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12133 = 9'h158 == _GEN_18214 ? phv_data_344 : _GEN_12132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12134 = 9'h159 == _GEN_18214 ? phv_data_345 : _GEN_12133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12135 = 9'h15a == _GEN_18214 ? phv_data_346 : _GEN_12134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12136 = 9'h15b == _GEN_18214 ? phv_data_347 : _GEN_12135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12137 = 9'h15c == _GEN_18214 ? phv_data_348 : _GEN_12136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12138 = 9'h15d == _GEN_18214 ? phv_data_349 : _GEN_12137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12139 = 9'h15e == _GEN_18214 ? phv_data_350 : _GEN_12138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12140 = 9'h15f == _GEN_18214 ? phv_data_351 : _GEN_12139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12141 = 9'h160 == _GEN_18214 ? phv_data_352 : _GEN_12140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12142 = 9'h161 == _GEN_18214 ? phv_data_353 : _GEN_12141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12143 = 9'h162 == _GEN_18214 ? phv_data_354 : _GEN_12142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12144 = 9'h163 == _GEN_18214 ? phv_data_355 : _GEN_12143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12145 = 9'h164 == _GEN_18214 ? phv_data_356 : _GEN_12144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12146 = 9'h165 == _GEN_18214 ? phv_data_357 : _GEN_12145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12147 = 9'h166 == _GEN_18214 ? phv_data_358 : _GEN_12146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12148 = 9'h167 == _GEN_18214 ? phv_data_359 : _GEN_12147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12149 = 9'h168 == _GEN_18214 ? phv_data_360 : _GEN_12148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12150 = 9'h169 == _GEN_18214 ? phv_data_361 : _GEN_12149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12151 = 9'h16a == _GEN_18214 ? phv_data_362 : _GEN_12150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12152 = 9'h16b == _GEN_18214 ? phv_data_363 : _GEN_12151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12153 = 9'h16c == _GEN_18214 ? phv_data_364 : _GEN_12152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12154 = 9'h16d == _GEN_18214 ? phv_data_365 : _GEN_12153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12155 = 9'h16e == _GEN_18214 ? phv_data_366 : _GEN_12154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12156 = 9'h16f == _GEN_18214 ? phv_data_367 : _GEN_12155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12157 = 9'h170 == _GEN_18214 ? phv_data_368 : _GEN_12156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12158 = 9'h171 == _GEN_18214 ? phv_data_369 : _GEN_12157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12159 = 9'h172 == _GEN_18214 ? phv_data_370 : _GEN_12158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12160 = 9'h173 == _GEN_18214 ? phv_data_371 : _GEN_12159; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12161 = 9'h174 == _GEN_18214 ? phv_data_372 : _GEN_12160; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12162 = 9'h175 == _GEN_18214 ? phv_data_373 : _GEN_12161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12163 = 9'h176 == _GEN_18214 ? phv_data_374 : _GEN_12162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12164 = 9'h177 == _GEN_18214 ? phv_data_375 : _GEN_12163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12165 = 9'h178 == _GEN_18214 ? phv_data_376 : _GEN_12164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12166 = 9'h179 == _GEN_18214 ? phv_data_377 : _GEN_12165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12167 = 9'h17a == _GEN_18214 ? phv_data_378 : _GEN_12166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12168 = 9'h17b == _GEN_18214 ? phv_data_379 : _GEN_12167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12169 = 9'h17c == _GEN_18214 ? phv_data_380 : _GEN_12168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12170 = 9'h17d == _GEN_18214 ? phv_data_381 : _GEN_12169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12171 = 9'h17e == _GEN_18214 ? phv_data_382 : _GEN_12170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12172 = 9'h17f == _GEN_18214 ? phv_data_383 : _GEN_12171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12173 = 9'h180 == _GEN_18214 ? phv_data_384 : _GEN_12172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12174 = 9'h181 == _GEN_18214 ? phv_data_385 : _GEN_12173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12175 = 9'h182 == _GEN_18214 ? phv_data_386 : _GEN_12174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12176 = 9'h183 == _GEN_18214 ? phv_data_387 : _GEN_12175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12177 = 9'h184 == _GEN_18214 ? phv_data_388 : _GEN_12176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12178 = 9'h185 == _GEN_18214 ? phv_data_389 : _GEN_12177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12179 = 9'h186 == _GEN_18214 ? phv_data_390 : _GEN_12178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12180 = 9'h187 == _GEN_18214 ? phv_data_391 : _GEN_12179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12181 = 9'h188 == _GEN_18214 ? phv_data_392 : _GEN_12180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12182 = 9'h189 == _GEN_18214 ? phv_data_393 : _GEN_12181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12183 = 9'h18a == _GEN_18214 ? phv_data_394 : _GEN_12182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12184 = 9'h18b == _GEN_18214 ? phv_data_395 : _GEN_12183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12185 = 9'h18c == _GEN_18214 ? phv_data_396 : _GEN_12184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12186 = 9'h18d == _GEN_18214 ? phv_data_397 : _GEN_12185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12187 = 9'h18e == _GEN_18214 ? phv_data_398 : _GEN_12186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12188 = 9'h18f == _GEN_18214 ? phv_data_399 : _GEN_12187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12189 = 9'h190 == _GEN_18214 ? phv_data_400 : _GEN_12188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12190 = 9'h191 == _GEN_18214 ? phv_data_401 : _GEN_12189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12191 = 9'h192 == _GEN_18214 ? phv_data_402 : _GEN_12190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12192 = 9'h193 == _GEN_18214 ? phv_data_403 : _GEN_12191; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12193 = 9'h194 == _GEN_18214 ? phv_data_404 : _GEN_12192; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12194 = 9'h195 == _GEN_18214 ? phv_data_405 : _GEN_12193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12195 = 9'h196 == _GEN_18214 ? phv_data_406 : _GEN_12194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12196 = 9'h197 == _GEN_18214 ? phv_data_407 : _GEN_12195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12197 = 9'h198 == _GEN_18214 ? phv_data_408 : _GEN_12196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12198 = 9'h199 == _GEN_18214 ? phv_data_409 : _GEN_12197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12199 = 9'h19a == _GEN_18214 ? phv_data_410 : _GEN_12198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12200 = 9'h19b == _GEN_18214 ? phv_data_411 : _GEN_12199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12201 = 9'h19c == _GEN_18214 ? phv_data_412 : _GEN_12200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12202 = 9'h19d == _GEN_18214 ? phv_data_413 : _GEN_12201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12203 = 9'h19e == _GEN_18214 ? phv_data_414 : _GEN_12202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12204 = 9'h19f == _GEN_18214 ? phv_data_415 : _GEN_12203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12205 = 9'h1a0 == _GEN_18214 ? phv_data_416 : _GEN_12204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12206 = 9'h1a1 == _GEN_18214 ? phv_data_417 : _GEN_12205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12207 = 9'h1a2 == _GEN_18214 ? phv_data_418 : _GEN_12206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12208 = 9'h1a3 == _GEN_18214 ? phv_data_419 : _GEN_12207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12209 = 9'h1a4 == _GEN_18214 ? phv_data_420 : _GEN_12208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12210 = 9'h1a5 == _GEN_18214 ? phv_data_421 : _GEN_12209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12211 = 9'h1a6 == _GEN_18214 ? phv_data_422 : _GEN_12210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12212 = 9'h1a7 == _GEN_18214 ? phv_data_423 : _GEN_12211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12213 = 9'h1a8 == _GEN_18214 ? phv_data_424 : _GEN_12212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12214 = 9'h1a9 == _GEN_18214 ? phv_data_425 : _GEN_12213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12215 = 9'h1aa == _GEN_18214 ? phv_data_426 : _GEN_12214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12216 = 9'h1ab == _GEN_18214 ? phv_data_427 : _GEN_12215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12217 = 9'h1ac == _GEN_18214 ? phv_data_428 : _GEN_12216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12218 = 9'h1ad == _GEN_18214 ? phv_data_429 : _GEN_12217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12219 = 9'h1ae == _GEN_18214 ? phv_data_430 : _GEN_12218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12220 = 9'h1af == _GEN_18214 ? phv_data_431 : _GEN_12219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12221 = 9'h1b0 == _GEN_18214 ? phv_data_432 : _GEN_12220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12222 = 9'h1b1 == _GEN_18214 ? phv_data_433 : _GEN_12221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12223 = 9'h1b2 == _GEN_18214 ? phv_data_434 : _GEN_12222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12224 = 9'h1b3 == _GEN_18214 ? phv_data_435 : _GEN_12223; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12225 = 9'h1b4 == _GEN_18214 ? phv_data_436 : _GEN_12224; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12226 = 9'h1b5 == _GEN_18214 ? phv_data_437 : _GEN_12225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12227 = 9'h1b6 == _GEN_18214 ? phv_data_438 : _GEN_12226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12228 = 9'h1b7 == _GEN_18214 ? phv_data_439 : _GEN_12227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12229 = 9'h1b8 == _GEN_18214 ? phv_data_440 : _GEN_12228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12230 = 9'h1b9 == _GEN_18214 ? phv_data_441 : _GEN_12229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12231 = 9'h1ba == _GEN_18214 ? phv_data_442 : _GEN_12230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12232 = 9'h1bb == _GEN_18214 ? phv_data_443 : _GEN_12231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12233 = 9'h1bc == _GEN_18214 ? phv_data_444 : _GEN_12232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12234 = 9'h1bd == _GEN_18214 ? phv_data_445 : _GEN_12233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12235 = 9'h1be == _GEN_18214 ? phv_data_446 : _GEN_12234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12236 = 9'h1bf == _GEN_18214 ? phv_data_447 : _GEN_12235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12237 = 9'h1c0 == _GEN_18214 ? phv_data_448 : _GEN_12236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12238 = 9'h1c1 == _GEN_18214 ? phv_data_449 : _GEN_12237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12239 = 9'h1c2 == _GEN_18214 ? phv_data_450 : _GEN_12238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12240 = 9'h1c3 == _GEN_18214 ? phv_data_451 : _GEN_12239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12241 = 9'h1c4 == _GEN_18214 ? phv_data_452 : _GEN_12240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12242 = 9'h1c5 == _GEN_18214 ? phv_data_453 : _GEN_12241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12243 = 9'h1c6 == _GEN_18214 ? phv_data_454 : _GEN_12242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12244 = 9'h1c7 == _GEN_18214 ? phv_data_455 : _GEN_12243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12245 = 9'h1c8 == _GEN_18214 ? phv_data_456 : _GEN_12244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12246 = 9'h1c9 == _GEN_18214 ? phv_data_457 : _GEN_12245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12247 = 9'h1ca == _GEN_18214 ? phv_data_458 : _GEN_12246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12248 = 9'h1cb == _GEN_18214 ? phv_data_459 : _GEN_12247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12249 = 9'h1cc == _GEN_18214 ? phv_data_460 : _GEN_12248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12250 = 9'h1cd == _GEN_18214 ? phv_data_461 : _GEN_12249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12251 = 9'h1ce == _GEN_18214 ? phv_data_462 : _GEN_12250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12252 = 9'h1cf == _GEN_18214 ? phv_data_463 : _GEN_12251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12253 = 9'h1d0 == _GEN_18214 ? phv_data_464 : _GEN_12252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12254 = 9'h1d1 == _GEN_18214 ? phv_data_465 : _GEN_12253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12255 = 9'h1d2 == _GEN_18214 ? phv_data_466 : _GEN_12254; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12256 = 9'h1d3 == _GEN_18214 ? phv_data_467 : _GEN_12255; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12257 = 9'h1d4 == _GEN_18214 ? phv_data_468 : _GEN_12256; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12258 = 9'h1d5 == _GEN_18214 ? phv_data_469 : _GEN_12257; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12259 = 9'h1d6 == _GEN_18214 ? phv_data_470 : _GEN_12258; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12260 = 9'h1d7 == _GEN_18214 ? phv_data_471 : _GEN_12259; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12261 = 9'h1d8 == _GEN_18214 ? phv_data_472 : _GEN_12260; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12262 = 9'h1d9 == _GEN_18214 ? phv_data_473 : _GEN_12261; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12263 = 9'h1da == _GEN_18214 ? phv_data_474 : _GEN_12262; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12264 = 9'h1db == _GEN_18214 ? phv_data_475 : _GEN_12263; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12265 = 9'h1dc == _GEN_18214 ? phv_data_476 : _GEN_12264; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12266 = 9'h1dd == _GEN_18214 ? phv_data_477 : _GEN_12265; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12267 = 9'h1de == _GEN_18214 ? phv_data_478 : _GEN_12266; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12268 = 9'h1df == _GEN_18214 ? phv_data_479 : _GEN_12267; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12269 = 9'h1e0 == _GEN_18214 ? phv_data_480 : _GEN_12268; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12270 = 9'h1e1 == _GEN_18214 ? phv_data_481 : _GEN_12269; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12271 = 9'h1e2 == _GEN_18214 ? phv_data_482 : _GEN_12270; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12272 = 9'h1e3 == _GEN_18214 ? phv_data_483 : _GEN_12271; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12273 = 9'h1e4 == _GEN_18214 ? phv_data_484 : _GEN_12272; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12274 = 9'h1e5 == _GEN_18214 ? phv_data_485 : _GEN_12273; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12275 = 9'h1e6 == _GEN_18214 ? phv_data_486 : _GEN_12274; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12276 = 9'h1e7 == _GEN_18214 ? phv_data_487 : _GEN_12275; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12277 = 9'h1e8 == _GEN_18214 ? phv_data_488 : _GEN_12276; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12278 = 9'h1e9 == _GEN_18214 ? phv_data_489 : _GEN_12277; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12279 = 9'h1ea == _GEN_18214 ? phv_data_490 : _GEN_12278; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12280 = 9'h1eb == _GEN_18214 ? phv_data_491 : _GEN_12279; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12281 = 9'h1ec == _GEN_18214 ? phv_data_492 : _GEN_12280; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12282 = 9'h1ed == _GEN_18214 ? phv_data_493 : _GEN_12281; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12283 = 9'h1ee == _GEN_18214 ? phv_data_494 : _GEN_12282; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12284 = 9'h1ef == _GEN_18214 ? phv_data_495 : _GEN_12283; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12285 = 9'h1f0 == _GEN_18214 ? phv_data_496 : _GEN_12284; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12286 = 9'h1f1 == _GEN_18214 ? phv_data_497 : _GEN_12285; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12287 = 9'h1f2 == _GEN_18214 ? phv_data_498 : _GEN_12286; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12288 = 9'h1f3 == _GEN_18214 ? phv_data_499 : _GEN_12287; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12289 = 9'h1f4 == _GEN_18214 ? phv_data_500 : _GEN_12288; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12290 = 9'h1f5 == _GEN_18214 ? phv_data_501 : _GEN_12289; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12291 = 9'h1f6 == _GEN_18214 ? phv_data_502 : _GEN_12290; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12292 = 9'h1f7 == _GEN_18214 ? phv_data_503 : _GEN_12291; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12293 = 9'h1f8 == _GEN_18214 ? phv_data_504 : _GEN_12292; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12294 = 9'h1f9 == _GEN_18214 ? phv_data_505 : _GEN_12293; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12295 = 9'h1fa == _GEN_18214 ? phv_data_506 : _GEN_12294; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12296 = 9'h1fb == _GEN_18214 ? phv_data_507 : _GEN_12295; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12297 = 9'h1fc == _GEN_18214 ? phv_data_508 : _GEN_12296; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12298 = 9'h1fd == _GEN_18214 ? phv_data_509 : _GEN_12297; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12299 = 9'h1fe == _GEN_18214 ? phv_data_510 : _GEN_12298; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12300 = 9'h1ff == _GEN_18214 ? phv_data_511 : _GEN_12299; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _match_key_qbytes_5_T_3 = {_GEN_11788,_GEN_12300,_GEN_10764,_GEN_11276}; // @[Cat.scala 30:58]
  wire [31:0] match_key_qbytes_5 = local_offset_5 < end_offset ? _match_key_qbytes_5_T_3 : 32'h0; // @[matcher.scala 88:54 matcher.scala 89:45 matcher.scala 97:45]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_256 = phv_data_256; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_257 = phv_data_257; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_258 = phv_data_258; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_259 = phv_data_259; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_260 = phv_data_260; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_261 = phv_data_261; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_262 = phv_data_262; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_263 = phv_data_263; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_264 = phv_data_264; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_265 = phv_data_265; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_266 = phv_data_266; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_267 = phv_data_267; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_268 = phv_data_268; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_269 = phv_data_269; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_270 = phv_data_270; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_271 = phv_data_271; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_272 = phv_data_272; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_273 = phv_data_273; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_274 = phv_data_274; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_275 = phv_data_275; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_276 = phv_data_276; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_277 = phv_data_277; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_278 = phv_data_278; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_279 = phv_data_279; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_280 = phv_data_280; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_281 = phv_data_281; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_282 = phv_data_282; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_283 = phv_data_283; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_284 = phv_data_284; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_285 = phv_data_285; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_286 = phv_data_286; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_287 = phv_data_287; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_288 = phv_data_288; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_289 = phv_data_289; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_290 = phv_data_290; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_291 = phv_data_291; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_292 = phv_data_292; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_293 = phv_data_293; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_294 = phv_data_294; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_295 = phv_data_295; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_296 = phv_data_296; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_297 = phv_data_297; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_298 = phv_data_298; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_299 = phv_data_299; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_300 = phv_data_300; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_301 = phv_data_301; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_302 = phv_data_302; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_303 = phv_data_303; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_304 = phv_data_304; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_305 = phv_data_305; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_306 = phv_data_306; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_307 = phv_data_307; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_308 = phv_data_308; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_309 = phv_data_309; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_310 = phv_data_310; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_311 = phv_data_311; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_312 = phv_data_312; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_313 = phv_data_313; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_314 = phv_data_314; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_315 = phv_data_315; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_316 = phv_data_316; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_317 = phv_data_317; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_318 = phv_data_318; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_319 = phv_data_319; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_320 = phv_data_320; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_321 = phv_data_321; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_322 = phv_data_322; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_323 = phv_data_323; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_324 = phv_data_324; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_325 = phv_data_325; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_326 = phv_data_326; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_327 = phv_data_327; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_328 = phv_data_328; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_329 = phv_data_329; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_330 = phv_data_330; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_331 = phv_data_331; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_332 = phv_data_332; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_333 = phv_data_333; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_334 = phv_data_334; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_335 = phv_data_335; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_336 = phv_data_336; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_337 = phv_data_337; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_338 = phv_data_338; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_339 = phv_data_339; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_340 = phv_data_340; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_341 = phv_data_341; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_342 = phv_data_342; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_343 = phv_data_343; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_344 = phv_data_344; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_345 = phv_data_345; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_346 = phv_data_346; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_347 = phv_data_347; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_348 = phv_data_348; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_349 = phv_data_349; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_350 = phv_data_350; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_351 = phv_data_351; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_352 = phv_data_352; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_353 = phv_data_353; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_354 = phv_data_354; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_355 = phv_data_355; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_356 = phv_data_356; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_357 = phv_data_357; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_358 = phv_data_358; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_359 = phv_data_359; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_360 = phv_data_360; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_361 = phv_data_361; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_362 = phv_data_362; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_363 = phv_data_363; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_364 = phv_data_364; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_365 = phv_data_365; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_366 = phv_data_366; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_367 = phv_data_367; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_368 = phv_data_368; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_369 = phv_data_369; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_370 = phv_data_370; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_371 = phv_data_371; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_372 = phv_data_372; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_373 = phv_data_373; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_374 = phv_data_374; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_375 = phv_data_375; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_376 = phv_data_376; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_377 = phv_data_377; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_378 = phv_data_378; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_379 = phv_data_379; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_380 = phv_data_380; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_381 = phv_data_381; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_382 = phv_data_382; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_383 = phv_data_383; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_384 = phv_data_384; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_385 = phv_data_385; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_386 = phv_data_386; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_387 = phv_data_387; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_388 = phv_data_388; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_389 = phv_data_389; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_390 = phv_data_390; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_391 = phv_data_391; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_392 = phv_data_392; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_393 = phv_data_393; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_394 = phv_data_394; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_395 = phv_data_395; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_396 = phv_data_396; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_397 = phv_data_397; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_398 = phv_data_398; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_399 = phv_data_399; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_400 = phv_data_400; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_401 = phv_data_401; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_402 = phv_data_402; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_403 = phv_data_403; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_404 = phv_data_404; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_405 = phv_data_405; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_406 = phv_data_406; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_407 = phv_data_407; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_408 = phv_data_408; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_409 = phv_data_409; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_410 = phv_data_410; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_411 = phv_data_411; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_412 = phv_data_412; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_413 = phv_data_413; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_414 = phv_data_414; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_415 = phv_data_415; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_416 = phv_data_416; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_417 = phv_data_417; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_418 = phv_data_418; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_419 = phv_data_419; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_420 = phv_data_420; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_421 = phv_data_421; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_422 = phv_data_422; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_423 = phv_data_423; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_424 = phv_data_424; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_425 = phv_data_425; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_426 = phv_data_426; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_427 = phv_data_427; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_428 = phv_data_428; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_429 = phv_data_429; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_430 = phv_data_430; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_431 = phv_data_431; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_432 = phv_data_432; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_433 = phv_data_433; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_434 = phv_data_434; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_435 = phv_data_435; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_436 = phv_data_436; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_437 = phv_data_437; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_438 = phv_data_438; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_439 = phv_data_439; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_440 = phv_data_440; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_441 = phv_data_441; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_442 = phv_data_442; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_443 = phv_data_443; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_444 = phv_data_444; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_445 = phv_data_445; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_446 = phv_data_446; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_447 = phv_data_447; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_448 = phv_data_448; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_449 = phv_data_449; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_450 = phv_data_450; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_451 = phv_data_451; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_452 = phv_data_452; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_453 = phv_data_453; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_454 = phv_data_454; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_455 = phv_data_455; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_456 = phv_data_456; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_457 = phv_data_457; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_458 = phv_data_458; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_459 = phv_data_459; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_460 = phv_data_460; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_461 = phv_data_461; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_462 = phv_data_462; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_463 = phv_data_463; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_464 = phv_data_464; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_465 = phv_data_465; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_466 = phv_data_466; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_467 = phv_data_467; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_468 = phv_data_468; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_469 = phv_data_469; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_470 = phv_data_470; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_471 = phv_data_471; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_472 = phv_data_472; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_473 = phv_data_473; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_474 = phv_data_474; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_475 = phv_data_475; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_476 = phv_data_476; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_477 = phv_data_477; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_478 = phv_data_478; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_479 = phv_data_479; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_480 = phv_data_480; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_481 = phv_data_481; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_482 = phv_data_482; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_483 = phv_data_483; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_484 = phv_data_484; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_485 = phv_data_485; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_486 = phv_data_486; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_487 = phv_data_487; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_488 = phv_data_488; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_489 = phv_data_489; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_490 = phv_data_490; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_491 = phv_data_491; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_492 = phv_data_492; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_493 = phv_data_493; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_494 = phv_data_494; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_495 = phv_data_495; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_496 = phv_data_496; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_497 = phv_data_497; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_498 = phv_data_498; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_499 = phv_data_499; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_500 = phv_data_500; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_501 = phv_data_501; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_502 = phv_data_502; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_503 = phv_data_503; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_504 = phv_data_504; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_505 = phv_data_505; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_506 = phv_data_506; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_507 = phv_data_507; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_508 = phv_data_508; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_509 = phv_data_509; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_510 = phv_data_510; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_data_511 = phv_data_511; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher.scala 69:29]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher.scala 69:29]
  assign io_bias_out = key_offset[1:0]; // @[matcher.scala 79:38]
  assign io_match_key_bytes_0 = phv_is_valid_processor ? match_key_qbytes_0[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_1 = phv_is_valid_processor ? match_key_qbytes_0[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_2 = phv_is_valid_processor ? match_key_qbytes_0[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_3 = phv_is_valid_processor ? match_key_qbytes_0[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_4 = phv_is_valid_processor ? match_key_qbytes_1[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_5 = phv_is_valid_processor ? match_key_qbytes_1[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_6 = phv_is_valid_processor ? match_key_qbytes_1[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_7 = phv_is_valid_processor ? match_key_qbytes_1[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_8 = phv_is_valid_processor ? match_key_qbytes_2[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_9 = phv_is_valid_processor ? match_key_qbytes_2[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_10 = phv_is_valid_processor ? match_key_qbytes_2[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_11 = phv_is_valid_processor ? match_key_qbytes_2[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_12 = phv_is_valid_processor ? match_key_qbytes_3[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_13 = phv_is_valid_processor ? match_key_qbytes_3[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_14 = phv_is_valid_processor ? match_key_qbytes_3[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_15 = phv_is_valid_processor ? match_key_qbytes_3[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_16 = phv_is_valid_processor ? match_key_qbytes_4[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_17 = phv_is_valid_processor ? match_key_qbytes_4[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_18 = phv_is_valid_processor ? match_key_qbytes_4[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_19 = phv_is_valid_processor ? match_key_qbytes_4[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_20 = phv_is_valid_processor ? match_key_qbytes_5[7:0] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_21 = phv_is_valid_processor ? match_key_qbytes_5[15:8] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_22 = phv_is_valid_processor ? match_key_qbytes_5[23:16] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  assign io_match_key_bytes_23 = phv_is_valid_processor ? match_key_qbytes_5[31:24] : 8'h0; // @[matcher.scala 81:43 matcher.scala 100:51 matcher.scala 105:43]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher.scala 68:17]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher.scala 68:17]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher.scala 68:17]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher.scala 68:17]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher.scala 68:17]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher.scala 68:17]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher.scala 68:17]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher.scala 68:17]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher.scala 68:17]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher.scala 68:17]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher.scala 68:17]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher.scala 68:17]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher.scala 68:17]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher.scala 68:17]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher.scala 68:17]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher.scala 68:17]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher.scala 68:17]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher.scala 68:17]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher.scala 68:17]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher.scala 68:17]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher.scala 68:17]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher.scala 68:17]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher.scala 68:17]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher.scala 68:17]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher.scala 68:17]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher.scala 68:17]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher.scala 68:17]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher.scala 68:17]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher.scala 68:17]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher.scala 68:17]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher.scala 68:17]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher.scala 68:17]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher.scala 68:17]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher.scala 68:17]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher.scala 68:17]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher.scala 68:17]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher.scala 68:17]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher.scala 68:17]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher.scala 68:17]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher.scala 68:17]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher.scala 68:17]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher.scala 68:17]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher.scala 68:17]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher.scala 68:17]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher.scala 68:17]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher.scala 68:17]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher.scala 68:17]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher.scala 68:17]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher.scala 68:17]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher.scala 68:17]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher.scala 68:17]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher.scala 68:17]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher.scala 68:17]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher.scala 68:17]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher.scala 68:17]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher.scala 68:17]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher.scala 68:17]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher.scala 68:17]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher.scala 68:17]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher.scala 68:17]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher.scala 68:17]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher.scala 68:17]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher.scala 68:17]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher.scala 68:17]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher.scala 68:17]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher.scala 68:17]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher.scala 68:17]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher.scala 68:17]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher.scala 68:17]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher.scala 68:17]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher.scala 68:17]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher.scala 68:17]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher.scala 68:17]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher.scala 68:17]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher.scala 68:17]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher.scala 68:17]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher.scala 68:17]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher.scala 68:17]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher.scala 68:17]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher.scala 68:17]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher.scala 68:17]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher.scala 68:17]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher.scala 68:17]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher.scala 68:17]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher.scala 68:17]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher.scala 68:17]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher.scala 68:17]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher.scala 68:17]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher.scala 68:17]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher.scala 68:17]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher.scala 68:17]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher.scala 68:17]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher.scala 68:17]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher.scala 68:17]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher.scala 68:17]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher.scala 68:17]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher.scala 68:17]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher.scala 68:17]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher.scala 68:17]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher.scala 68:17]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher.scala 68:17]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher.scala 68:17]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher.scala 68:17]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher.scala 68:17]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher.scala 68:17]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher.scala 68:17]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher.scala 68:17]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher.scala 68:17]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher.scala 68:17]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher.scala 68:17]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher.scala 68:17]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher.scala 68:17]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher.scala 68:17]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher.scala 68:17]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher.scala 68:17]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher.scala 68:17]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher.scala 68:17]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher.scala 68:17]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher.scala 68:17]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher.scala 68:17]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher.scala 68:17]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher.scala 68:17]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher.scala 68:17]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher.scala 68:17]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher.scala 68:17]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher.scala 68:17]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher.scala 68:17]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher.scala 68:17]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher.scala 68:17]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher.scala 68:17]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher.scala 68:17]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher.scala 68:17]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher.scala 68:17]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher.scala 68:17]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher.scala 68:17]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher.scala 68:17]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher.scala 68:17]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher.scala 68:17]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher.scala 68:17]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher.scala 68:17]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher.scala 68:17]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher.scala 68:17]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher.scala 68:17]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher.scala 68:17]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher.scala 68:17]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher.scala 68:17]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher.scala 68:17]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher.scala 68:17]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher.scala 68:17]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher.scala 68:17]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher.scala 68:17]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher.scala 68:17]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher.scala 68:17]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher.scala 68:17]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher.scala 68:17]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher.scala 68:17]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher.scala 68:17]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher.scala 68:17]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher.scala 68:17]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher.scala 68:17]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[matcher.scala 68:17]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[matcher.scala 68:17]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[matcher.scala 68:17]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[matcher.scala 68:17]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[matcher.scala 68:17]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[matcher.scala 68:17]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[matcher.scala 68:17]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[matcher.scala 68:17]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[matcher.scala 68:17]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[matcher.scala 68:17]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[matcher.scala 68:17]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[matcher.scala 68:17]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[matcher.scala 68:17]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[matcher.scala 68:17]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[matcher.scala 68:17]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[matcher.scala 68:17]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[matcher.scala 68:17]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[matcher.scala 68:17]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[matcher.scala 68:17]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[matcher.scala 68:17]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[matcher.scala 68:17]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[matcher.scala 68:17]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[matcher.scala 68:17]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[matcher.scala 68:17]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[matcher.scala 68:17]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[matcher.scala 68:17]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[matcher.scala 68:17]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[matcher.scala 68:17]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[matcher.scala 68:17]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[matcher.scala 68:17]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[matcher.scala 68:17]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[matcher.scala 68:17]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[matcher.scala 68:17]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[matcher.scala 68:17]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[matcher.scala 68:17]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[matcher.scala 68:17]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[matcher.scala 68:17]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[matcher.scala 68:17]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[matcher.scala 68:17]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[matcher.scala 68:17]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[matcher.scala 68:17]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[matcher.scala 68:17]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[matcher.scala 68:17]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[matcher.scala 68:17]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[matcher.scala 68:17]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[matcher.scala 68:17]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[matcher.scala 68:17]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[matcher.scala 68:17]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[matcher.scala 68:17]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[matcher.scala 68:17]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[matcher.scala 68:17]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[matcher.scala 68:17]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[matcher.scala 68:17]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[matcher.scala 68:17]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[matcher.scala 68:17]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[matcher.scala 68:17]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[matcher.scala 68:17]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[matcher.scala 68:17]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[matcher.scala 68:17]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[matcher.scala 68:17]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[matcher.scala 68:17]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[matcher.scala 68:17]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[matcher.scala 68:17]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[matcher.scala 68:17]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[matcher.scala 68:17]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[matcher.scala 68:17]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[matcher.scala 68:17]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[matcher.scala 68:17]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[matcher.scala 68:17]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[matcher.scala 68:17]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[matcher.scala 68:17]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[matcher.scala 68:17]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[matcher.scala 68:17]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[matcher.scala 68:17]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[matcher.scala 68:17]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[matcher.scala 68:17]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[matcher.scala 68:17]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[matcher.scala 68:17]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[matcher.scala 68:17]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[matcher.scala 68:17]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[matcher.scala 68:17]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[matcher.scala 68:17]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[matcher.scala 68:17]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[matcher.scala 68:17]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[matcher.scala 68:17]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[matcher.scala 68:17]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[matcher.scala 68:17]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[matcher.scala 68:17]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[matcher.scala 68:17]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[matcher.scala 68:17]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[matcher.scala 68:17]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[matcher.scala 68:17]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[matcher.scala 68:17]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[matcher.scala 68:17]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[matcher.scala 68:17]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[matcher.scala 68:17]
    phv_data_256 <= io_pipe_phv_in_data_256; // @[matcher.scala 68:17]
    phv_data_257 <= io_pipe_phv_in_data_257; // @[matcher.scala 68:17]
    phv_data_258 <= io_pipe_phv_in_data_258; // @[matcher.scala 68:17]
    phv_data_259 <= io_pipe_phv_in_data_259; // @[matcher.scala 68:17]
    phv_data_260 <= io_pipe_phv_in_data_260; // @[matcher.scala 68:17]
    phv_data_261 <= io_pipe_phv_in_data_261; // @[matcher.scala 68:17]
    phv_data_262 <= io_pipe_phv_in_data_262; // @[matcher.scala 68:17]
    phv_data_263 <= io_pipe_phv_in_data_263; // @[matcher.scala 68:17]
    phv_data_264 <= io_pipe_phv_in_data_264; // @[matcher.scala 68:17]
    phv_data_265 <= io_pipe_phv_in_data_265; // @[matcher.scala 68:17]
    phv_data_266 <= io_pipe_phv_in_data_266; // @[matcher.scala 68:17]
    phv_data_267 <= io_pipe_phv_in_data_267; // @[matcher.scala 68:17]
    phv_data_268 <= io_pipe_phv_in_data_268; // @[matcher.scala 68:17]
    phv_data_269 <= io_pipe_phv_in_data_269; // @[matcher.scala 68:17]
    phv_data_270 <= io_pipe_phv_in_data_270; // @[matcher.scala 68:17]
    phv_data_271 <= io_pipe_phv_in_data_271; // @[matcher.scala 68:17]
    phv_data_272 <= io_pipe_phv_in_data_272; // @[matcher.scala 68:17]
    phv_data_273 <= io_pipe_phv_in_data_273; // @[matcher.scala 68:17]
    phv_data_274 <= io_pipe_phv_in_data_274; // @[matcher.scala 68:17]
    phv_data_275 <= io_pipe_phv_in_data_275; // @[matcher.scala 68:17]
    phv_data_276 <= io_pipe_phv_in_data_276; // @[matcher.scala 68:17]
    phv_data_277 <= io_pipe_phv_in_data_277; // @[matcher.scala 68:17]
    phv_data_278 <= io_pipe_phv_in_data_278; // @[matcher.scala 68:17]
    phv_data_279 <= io_pipe_phv_in_data_279; // @[matcher.scala 68:17]
    phv_data_280 <= io_pipe_phv_in_data_280; // @[matcher.scala 68:17]
    phv_data_281 <= io_pipe_phv_in_data_281; // @[matcher.scala 68:17]
    phv_data_282 <= io_pipe_phv_in_data_282; // @[matcher.scala 68:17]
    phv_data_283 <= io_pipe_phv_in_data_283; // @[matcher.scala 68:17]
    phv_data_284 <= io_pipe_phv_in_data_284; // @[matcher.scala 68:17]
    phv_data_285 <= io_pipe_phv_in_data_285; // @[matcher.scala 68:17]
    phv_data_286 <= io_pipe_phv_in_data_286; // @[matcher.scala 68:17]
    phv_data_287 <= io_pipe_phv_in_data_287; // @[matcher.scala 68:17]
    phv_data_288 <= io_pipe_phv_in_data_288; // @[matcher.scala 68:17]
    phv_data_289 <= io_pipe_phv_in_data_289; // @[matcher.scala 68:17]
    phv_data_290 <= io_pipe_phv_in_data_290; // @[matcher.scala 68:17]
    phv_data_291 <= io_pipe_phv_in_data_291; // @[matcher.scala 68:17]
    phv_data_292 <= io_pipe_phv_in_data_292; // @[matcher.scala 68:17]
    phv_data_293 <= io_pipe_phv_in_data_293; // @[matcher.scala 68:17]
    phv_data_294 <= io_pipe_phv_in_data_294; // @[matcher.scala 68:17]
    phv_data_295 <= io_pipe_phv_in_data_295; // @[matcher.scala 68:17]
    phv_data_296 <= io_pipe_phv_in_data_296; // @[matcher.scala 68:17]
    phv_data_297 <= io_pipe_phv_in_data_297; // @[matcher.scala 68:17]
    phv_data_298 <= io_pipe_phv_in_data_298; // @[matcher.scala 68:17]
    phv_data_299 <= io_pipe_phv_in_data_299; // @[matcher.scala 68:17]
    phv_data_300 <= io_pipe_phv_in_data_300; // @[matcher.scala 68:17]
    phv_data_301 <= io_pipe_phv_in_data_301; // @[matcher.scala 68:17]
    phv_data_302 <= io_pipe_phv_in_data_302; // @[matcher.scala 68:17]
    phv_data_303 <= io_pipe_phv_in_data_303; // @[matcher.scala 68:17]
    phv_data_304 <= io_pipe_phv_in_data_304; // @[matcher.scala 68:17]
    phv_data_305 <= io_pipe_phv_in_data_305; // @[matcher.scala 68:17]
    phv_data_306 <= io_pipe_phv_in_data_306; // @[matcher.scala 68:17]
    phv_data_307 <= io_pipe_phv_in_data_307; // @[matcher.scala 68:17]
    phv_data_308 <= io_pipe_phv_in_data_308; // @[matcher.scala 68:17]
    phv_data_309 <= io_pipe_phv_in_data_309; // @[matcher.scala 68:17]
    phv_data_310 <= io_pipe_phv_in_data_310; // @[matcher.scala 68:17]
    phv_data_311 <= io_pipe_phv_in_data_311; // @[matcher.scala 68:17]
    phv_data_312 <= io_pipe_phv_in_data_312; // @[matcher.scala 68:17]
    phv_data_313 <= io_pipe_phv_in_data_313; // @[matcher.scala 68:17]
    phv_data_314 <= io_pipe_phv_in_data_314; // @[matcher.scala 68:17]
    phv_data_315 <= io_pipe_phv_in_data_315; // @[matcher.scala 68:17]
    phv_data_316 <= io_pipe_phv_in_data_316; // @[matcher.scala 68:17]
    phv_data_317 <= io_pipe_phv_in_data_317; // @[matcher.scala 68:17]
    phv_data_318 <= io_pipe_phv_in_data_318; // @[matcher.scala 68:17]
    phv_data_319 <= io_pipe_phv_in_data_319; // @[matcher.scala 68:17]
    phv_data_320 <= io_pipe_phv_in_data_320; // @[matcher.scala 68:17]
    phv_data_321 <= io_pipe_phv_in_data_321; // @[matcher.scala 68:17]
    phv_data_322 <= io_pipe_phv_in_data_322; // @[matcher.scala 68:17]
    phv_data_323 <= io_pipe_phv_in_data_323; // @[matcher.scala 68:17]
    phv_data_324 <= io_pipe_phv_in_data_324; // @[matcher.scala 68:17]
    phv_data_325 <= io_pipe_phv_in_data_325; // @[matcher.scala 68:17]
    phv_data_326 <= io_pipe_phv_in_data_326; // @[matcher.scala 68:17]
    phv_data_327 <= io_pipe_phv_in_data_327; // @[matcher.scala 68:17]
    phv_data_328 <= io_pipe_phv_in_data_328; // @[matcher.scala 68:17]
    phv_data_329 <= io_pipe_phv_in_data_329; // @[matcher.scala 68:17]
    phv_data_330 <= io_pipe_phv_in_data_330; // @[matcher.scala 68:17]
    phv_data_331 <= io_pipe_phv_in_data_331; // @[matcher.scala 68:17]
    phv_data_332 <= io_pipe_phv_in_data_332; // @[matcher.scala 68:17]
    phv_data_333 <= io_pipe_phv_in_data_333; // @[matcher.scala 68:17]
    phv_data_334 <= io_pipe_phv_in_data_334; // @[matcher.scala 68:17]
    phv_data_335 <= io_pipe_phv_in_data_335; // @[matcher.scala 68:17]
    phv_data_336 <= io_pipe_phv_in_data_336; // @[matcher.scala 68:17]
    phv_data_337 <= io_pipe_phv_in_data_337; // @[matcher.scala 68:17]
    phv_data_338 <= io_pipe_phv_in_data_338; // @[matcher.scala 68:17]
    phv_data_339 <= io_pipe_phv_in_data_339; // @[matcher.scala 68:17]
    phv_data_340 <= io_pipe_phv_in_data_340; // @[matcher.scala 68:17]
    phv_data_341 <= io_pipe_phv_in_data_341; // @[matcher.scala 68:17]
    phv_data_342 <= io_pipe_phv_in_data_342; // @[matcher.scala 68:17]
    phv_data_343 <= io_pipe_phv_in_data_343; // @[matcher.scala 68:17]
    phv_data_344 <= io_pipe_phv_in_data_344; // @[matcher.scala 68:17]
    phv_data_345 <= io_pipe_phv_in_data_345; // @[matcher.scala 68:17]
    phv_data_346 <= io_pipe_phv_in_data_346; // @[matcher.scala 68:17]
    phv_data_347 <= io_pipe_phv_in_data_347; // @[matcher.scala 68:17]
    phv_data_348 <= io_pipe_phv_in_data_348; // @[matcher.scala 68:17]
    phv_data_349 <= io_pipe_phv_in_data_349; // @[matcher.scala 68:17]
    phv_data_350 <= io_pipe_phv_in_data_350; // @[matcher.scala 68:17]
    phv_data_351 <= io_pipe_phv_in_data_351; // @[matcher.scala 68:17]
    phv_data_352 <= io_pipe_phv_in_data_352; // @[matcher.scala 68:17]
    phv_data_353 <= io_pipe_phv_in_data_353; // @[matcher.scala 68:17]
    phv_data_354 <= io_pipe_phv_in_data_354; // @[matcher.scala 68:17]
    phv_data_355 <= io_pipe_phv_in_data_355; // @[matcher.scala 68:17]
    phv_data_356 <= io_pipe_phv_in_data_356; // @[matcher.scala 68:17]
    phv_data_357 <= io_pipe_phv_in_data_357; // @[matcher.scala 68:17]
    phv_data_358 <= io_pipe_phv_in_data_358; // @[matcher.scala 68:17]
    phv_data_359 <= io_pipe_phv_in_data_359; // @[matcher.scala 68:17]
    phv_data_360 <= io_pipe_phv_in_data_360; // @[matcher.scala 68:17]
    phv_data_361 <= io_pipe_phv_in_data_361; // @[matcher.scala 68:17]
    phv_data_362 <= io_pipe_phv_in_data_362; // @[matcher.scala 68:17]
    phv_data_363 <= io_pipe_phv_in_data_363; // @[matcher.scala 68:17]
    phv_data_364 <= io_pipe_phv_in_data_364; // @[matcher.scala 68:17]
    phv_data_365 <= io_pipe_phv_in_data_365; // @[matcher.scala 68:17]
    phv_data_366 <= io_pipe_phv_in_data_366; // @[matcher.scala 68:17]
    phv_data_367 <= io_pipe_phv_in_data_367; // @[matcher.scala 68:17]
    phv_data_368 <= io_pipe_phv_in_data_368; // @[matcher.scala 68:17]
    phv_data_369 <= io_pipe_phv_in_data_369; // @[matcher.scala 68:17]
    phv_data_370 <= io_pipe_phv_in_data_370; // @[matcher.scala 68:17]
    phv_data_371 <= io_pipe_phv_in_data_371; // @[matcher.scala 68:17]
    phv_data_372 <= io_pipe_phv_in_data_372; // @[matcher.scala 68:17]
    phv_data_373 <= io_pipe_phv_in_data_373; // @[matcher.scala 68:17]
    phv_data_374 <= io_pipe_phv_in_data_374; // @[matcher.scala 68:17]
    phv_data_375 <= io_pipe_phv_in_data_375; // @[matcher.scala 68:17]
    phv_data_376 <= io_pipe_phv_in_data_376; // @[matcher.scala 68:17]
    phv_data_377 <= io_pipe_phv_in_data_377; // @[matcher.scala 68:17]
    phv_data_378 <= io_pipe_phv_in_data_378; // @[matcher.scala 68:17]
    phv_data_379 <= io_pipe_phv_in_data_379; // @[matcher.scala 68:17]
    phv_data_380 <= io_pipe_phv_in_data_380; // @[matcher.scala 68:17]
    phv_data_381 <= io_pipe_phv_in_data_381; // @[matcher.scala 68:17]
    phv_data_382 <= io_pipe_phv_in_data_382; // @[matcher.scala 68:17]
    phv_data_383 <= io_pipe_phv_in_data_383; // @[matcher.scala 68:17]
    phv_data_384 <= io_pipe_phv_in_data_384; // @[matcher.scala 68:17]
    phv_data_385 <= io_pipe_phv_in_data_385; // @[matcher.scala 68:17]
    phv_data_386 <= io_pipe_phv_in_data_386; // @[matcher.scala 68:17]
    phv_data_387 <= io_pipe_phv_in_data_387; // @[matcher.scala 68:17]
    phv_data_388 <= io_pipe_phv_in_data_388; // @[matcher.scala 68:17]
    phv_data_389 <= io_pipe_phv_in_data_389; // @[matcher.scala 68:17]
    phv_data_390 <= io_pipe_phv_in_data_390; // @[matcher.scala 68:17]
    phv_data_391 <= io_pipe_phv_in_data_391; // @[matcher.scala 68:17]
    phv_data_392 <= io_pipe_phv_in_data_392; // @[matcher.scala 68:17]
    phv_data_393 <= io_pipe_phv_in_data_393; // @[matcher.scala 68:17]
    phv_data_394 <= io_pipe_phv_in_data_394; // @[matcher.scala 68:17]
    phv_data_395 <= io_pipe_phv_in_data_395; // @[matcher.scala 68:17]
    phv_data_396 <= io_pipe_phv_in_data_396; // @[matcher.scala 68:17]
    phv_data_397 <= io_pipe_phv_in_data_397; // @[matcher.scala 68:17]
    phv_data_398 <= io_pipe_phv_in_data_398; // @[matcher.scala 68:17]
    phv_data_399 <= io_pipe_phv_in_data_399; // @[matcher.scala 68:17]
    phv_data_400 <= io_pipe_phv_in_data_400; // @[matcher.scala 68:17]
    phv_data_401 <= io_pipe_phv_in_data_401; // @[matcher.scala 68:17]
    phv_data_402 <= io_pipe_phv_in_data_402; // @[matcher.scala 68:17]
    phv_data_403 <= io_pipe_phv_in_data_403; // @[matcher.scala 68:17]
    phv_data_404 <= io_pipe_phv_in_data_404; // @[matcher.scala 68:17]
    phv_data_405 <= io_pipe_phv_in_data_405; // @[matcher.scala 68:17]
    phv_data_406 <= io_pipe_phv_in_data_406; // @[matcher.scala 68:17]
    phv_data_407 <= io_pipe_phv_in_data_407; // @[matcher.scala 68:17]
    phv_data_408 <= io_pipe_phv_in_data_408; // @[matcher.scala 68:17]
    phv_data_409 <= io_pipe_phv_in_data_409; // @[matcher.scala 68:17]
    phv_data_410 <= io_pipe_phv_in_data_410; // @[matcher.scala 68:17]
    phv_data_411 <= io_pipe_phv_in_data_411; // @[matcher.scala 68:17]
    phv_data_412 <= io_pipe_phv_in_data_412; // @[matcher.scala 68:17]
    phv_data_413 <= io_pipe_phv_in_data_413; // @[matcher.scala 68:17]
    phv_data_414 <= io_pipe_phv_in_data_414; // @[matcher.scala 68:17]
    phv_data_415 <= io_pipe_phv_in_data_415; // @[matcher.scala 68:17]
    phv_data_416 <= io_pipe_phv_in_data_416; // @[matcher.scala 68:17]
    phv_data_417 <= io_pipe_phv_in_data_417; // @[matcher.scala 68:17]
    phv_data_418 <= io_pipe_phv_in_data_418; // @[matcher.scala 68:17]
    phv_data_419 <= io_pipe_phv_in_data_419; // @[matcher.scala 68:17]
    phv_data_420 <= io_pipe_phv_in_data_420; // @[matcher.scala 68:17]
    phv_data_421 <= io_pipe_phv_in_data_421; // @[matcher.scala 68:17]
    phv_data_422 <= io_pipe_phv_in_data_422; // @[matcher.scala 68:17]
    phv_data_423 <= io_pipe_phv_in_data_423; // @[matcher.scala 68:17]
    phv_data_424 <= io_pipe_phv_in_data_424; // @[matcher.scala 68:17]
    phv_data_425 <= io_pipe_phv_in_data_425; // @[matcher.scala 68:17]
    phv_data_426 <= io_pipe_phv_in_data_426; // @[matcher.scala 68:17]
    phv_data_427 <= io_pipe_phv_in_data_427; // @[matcher.scala 68:17]
    phv_data_428 <= io_pipe_phv_in_data_428; // @[matcher.scala 68:17]
    phv_data_429 <= io_pipe_phv_in_data_429; // @[matcher.scala 68:17]
    phv_data_430 <= io_pipe_phv_in_data_430; // @[matcher.scala 68:17]
    phv_data_431 <= io_pipe_phv_in_data_431; // @[matcher.scala 68:17]
    phv_data_432 <= io_pipe_phv_in_data_432; // @[matcher.scala 68:17]
    phv_data_433 <= io_pipe_phv_in_data_433; // @[matcher.scala 68:17]
    phv_data_434 <= io_pipe_phv_in_data_434; // @[matcher.scala 68:17]
    phv_data_435 <= io_pipe_phv_in_data_435; // @[matcher.scala 68:17]
    phv_data_436 <= io_pipe_phv_in_data_436; // @[matcher.scala 68:17]
    phv_data_437 <= io_pipe_phv_in_data_437; // @[matcher.scala 68:17]
    phv_data_438 <= io_pipe_phv_in_data_438; // @[matcher.scala 68:17]
    phv_data_439 <= io_pipe_phv_in_data_439; // @[matcher.scala 68:17]
    phv_data_440 <= io_pipe_phv_in_data_440; // @[matcher.scala 68:17]
    phv_data_441 <= io_pipe_phv_in_data_441; // @[matcher.scala 68:17]
    phv_data_442 <= io_pipe_phv_in_data_442; // @[matcher.scala 68:17]
    phv_data_443 <= io_pipe_phv_in_data_443; // @[matcher.scala 68:17]
    phv_data_444 <= io_pipe_phv_in_data_444; // @[matcher.scala 68:17]
    phv_data_445 <= io_pipe_phv_in_data_445; // @[matcher.scala 68:17]
    phv_data_446 <= io_pipe_phv_in_data_446; // @[matcher.scala 68:17]
    phv_data_447 <= io_pipe_phv_in_data_447; // @[matcher.scala 68:17]
    phv_data_448 <= io_pipe_phv_in_data_448; // @[matcher.scala 68:17]
    phv_data_449 <= io_pipe_phv_in_data_449; // @[matcher.scala 68:17]
    phv_data_450 <= io_pipe_phv_in_data_450; // @[matcher.scala 68:17]
    phv_data_451 <= io_pipe_phv_in_data_451; // @[matcher.scala 68:17]
    phv_data_452 <= io_pipe_phv_in_data_452; // @[matcher.scala 68:17]
    phv_data_453 <= io_pipe_phv_in_data_453; // @[matcher.scala 68:17]
    phv_data_454 <= io_pipe_phv_in_data_454; // @[matcher.scala 68:17]
    phv_data_455 <= io_pipe_phv_in_data_455; // @[matcher.scala 68:17]
    phv_data_456 <= io_pipe_phv_in_data_456; // @[matcher.scala 68:17]
    phv_data_457 <= io_pipe_phv_in_data_457; // @[matcher.scala 68:17]
    phv_data_458 <= io_pipe_phv_in_data_458; // @[matcher.scala 68:17]
    phv_data_459 <= io_pipe_phv_in_data_459; // @[matcher.scala 68:17]
    phv_data_460 <= io_pipe_phv_in_data_460; // @[matcher.scala 68:17]
    phv_data_461 <= io_pipe_phv_in_data_461; // @[matcher.scala 68:17]
    phv_data_462 <= io_pipe_phv_in_data_462; // @[matcher.scala 68:17]
    phv_data_463 <= io_pipe_phv_in_data_463; // @[matcher.scala 68:17]
    phv_data_464 <= io_pipe_phv_in_data_464; // @[matcher.scala 68:17]
    phv_data_465 <= io_pipe_phv_in_data_465; // @[matcher.scala 68:17]
    phv_data_466 <= io_pipe_phv_in_data_466; // @[matcher.scala 68:17]
    phv_data_467 <= io_pipe_phv_in_data_467; // @[matcher.scala 68:17]
    phv_data_468 <= io_pipe_phv_in_data_468; // @[matcher.scala 68:17]
    phv_data_469 <= io_pipe_phv_in_data_469; // @[matcher.scala 68:17]
    phv_data_470 <= io_pipe_phv_in_data_470; // @[matcher.scala 68:17]
    phv_data_471 <= io_pipe_phv_in_data_471; // @[matcher.scala 68:17]
    phv_data_472 <= io_pipe_phv_in_data_472; // @[matcher.scala 68:17]
    phv_data_473 <= io_pipe_phv_in_data_473; // @[matcher.scala 68:17]
    phv_data_474 <= io_pipe_phv_in_data_474; // @[matcher.scala 68:17]
    phv_data_475 <= io_pipe_phv_in_data_475; // @[matcher.scala 68:17]
    phv_data_476 <= io_pipe_phv_in_data_476; // @[matcher.scala 68:17]
    phv_data_477 <= io_pipe_phv_in_data_477; // @[matcher.scala 68:17]
    phv_data_478 <= io_pipe_phv_in_data_478; // @[matcher.scala 68:17]
    phv_data_479 <= io_pipe_phv_in_data_479; // @[matcher.scala 68:17]
    phv_data_480 <= io_pipe_phv_in_data_480; // @[matcher.scala 68:17]
    phv_data_481 <= io_pipe_phv_in_data_481; // @[matcher.scala 68:17]
    phv_data_482 <= io_pipe_phv_in_data_482; // @[matcher.scala 68:17]
    phv_data_483 <= io_pipe_phv_in_data_483; // @[matcher.scala 68:17]
    phv_data_484 <= io_pipe_phv_in_data_484; // @[matcher.scala 68:17]
    phv_data_485 <= io_pipe_phv_in_data_485; // @[matcher.scala 68:17]
    phv_data_486 <= io_pipe_phv_in_data_486; // @[matcher.scala 68:17]
    phv_data_487 <= io_pipe_phv_in_data_487; // @[matcher.scala 68:17]
    phv_data_488 <= io_pipe_phv_in_data_488; // @[matcher.scala 68:17]
    phv_data_489 <= io_pipe_phv_in_data_489; // @[matcher.scala 68:17]
    phv_data_490 <= io_pipe_phv_in_data_490; // @[matcher.scala 68:17]
    phv_data_491 <= io_pipe_phv_in_data_491; // @[matcher.scala 68:17]
    phv_data_492 <= io_pipe_phv_in_data_492; // @[matcher.scala 68:17]
    phv_data_493 <= io_pipe_phv_in_data_493; // @[matcher.scala 68:17]
    phv_data_494 <= io_pipe_phv_in_data_494; // @[matcher.scala 68:17]
    phv_data_495 <= io_pipe_phv_in_data_495; // @[matcher.scala 68:17]
    phv_data_496 <= io_pipe_phv_in_data_496; // @[matcher.scala 68:17]
    phv_data_497 <= io_pipe_phv_in_data_497; // @[matcher.scala 68:17]
    phv_data_498 <= io_pipe_phv_in_data_498; // @[matcher.scala 68:17]
    phv_data_499 <= io_pipe_phv_in_data_499; // @[matcher.scala 68:17]
    phv_data_500 <= io_pipe_phv_in_data_500; // @[matcher.scala 68:17]
    phv_data_501 <= io_pipe_phv_in_data_501; // @[matcher.scala 68:17]
    phv_data_502 <= io_pipe_phv_in_data_502; // @[matcher.scala 68:17]
    phv_data_503 <= io_pipe_phv_in_data_503; // @[matcher.scala 68:17]
    phv_data_504 <= io_pipe_phv_in_data_504; // @[matcher.scala 68:17]
    phv_data_505 <= io_pipe_phv_in_data_505; // @[matcher.scala 68:17]
    phv_data_506 <= io_pipe_phv_in_data_506; // @[matcher.scala 68:17]
    phv_data_507 <= io_pipe_phv_in_data_507; // @[matcher.scala 68:17]
    phv_data_508 <= io_pipe_phv_in_data_508; // @[matcher.scala 68:17]
    phv_data_509 <= io_pipe_phv_in_data_509; // @[matcher.scala 68:17]
    phv_data_510 <= io_pipe_phv_in_data_510; // @[matcher.scala 68:17]
    phv_data_511 <= io_pipe_phv_in_data_511; // @[matcher.scala 68:17]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[matcher.scala 68:17]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[matcher.scala 68:17]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[matcher.scala 68:17]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[matcher.scala 68:17]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[matcher.scala 68:17]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[matcher.scala 68:17]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[matcher.scala 68:17]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[matcher.scala 68:17]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[matcher.scala 68:17]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[matcher.scala 68:17]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[matcher.scala 68:17]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[matcher.scala 68:17]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[matcher.scala 68:17]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[matcher.scala 68:17]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[matcher.scala 68:17]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[matcher.scala 68:17]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[matcher.scala 68:17]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[matcher.scala 68:17]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[matcher.scala 68:17]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[matcher.scala 68:17]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher.scala 68:17]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher.scala 68:17]
    key_offset <= io_key_offset_in; // @[matcher.scala 72:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_data_256 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  phv_data_257 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  phv_data_258 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  phv_data_259 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  phv_data_260 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  phv_data_261 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  phv_data_262 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  phv_data_263 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  phv_data_264 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  phv_data_265 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  phv_data_266 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  phv_data_267 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  phv_data_268 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  phv_data_269 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  phv_data_270 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  phv_data_271 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  phv_data_272 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_data_273 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_data_274 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  phv_data_275 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  phv_data_276 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  phv_data_277 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  phv_data_278 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  phv_data_279 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  phv_data_280 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  phv_data_281 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  phv_data_282 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  phv_data_283 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  phv_data_284 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  phv_data_285 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  phv_data_286 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  phv_data_287 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  phv_data_288 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  phv_data_289 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  phv_data_290 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  phv_data_291 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  phv_data_292 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  phv_data_293 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  phv_data_294 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  phv_data_295 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  phv_data_296 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  phv_data_297 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  phv_data_298 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  phv_data_299 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  phv_data_300 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  phv_data_301 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  phv_data_302 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  phv_data_303 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  phv_data_304 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  phv_data_305 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  phv_data_306 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  phv_data_307 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  phv_data_308 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  phv_data_309 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  phv_data_310 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  phv_data_311 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  phv_data_312 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  phv_data_313 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  phv_data_314 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  phv_data_315 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  phv_data_316 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  phv_data_317 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  phv_data_318 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  phv_data_319 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  phv_data_320 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  phv_data_321 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  phv_data_322 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  phv_data_323 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  phv_data_324 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  phv_data_325 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  phv_data_326 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  phv_data_327 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  phv_data_328 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  phv_data_329 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  phv_data_330 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  phv_data_331 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  phv_data_332 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  phv_data_333 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  phv_data_334 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  phv_data_335 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  phv_data_336 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  phv_data_337 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  phv_data_338 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  phv_data_339 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  phv_data_340 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  phv_data_341 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  phv_data_342 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  phv_data_343 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  phv_data_344 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  phv_data_345 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  phv_data_346 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  phv_data_347 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  phv_data_348 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  phv_data_349 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  phv_data_350 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  phv_data_351 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  phv_data_352 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  phv_data_353 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  phv_data_354 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  phv_data_355 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  phv_data_356 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  phv_data_357 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  phv_data_358 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  phv_data_359 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  phv_data_360 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  phv_data_361 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  phv_data_362 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  phv_data_363 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  phv_data_364 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  phv_data_365 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  phv_data_366 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  phv_data_367 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  phv_data_368 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  phv_data_369 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  phv_data_370 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  phv_data_371 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  phv_data_372 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  phv_data_373 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  phv_data_374 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  phv_data_375 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  phv_data_376 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  phv_data_377 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  phv_data_378 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  phv_data_379 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  phv_data_380 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  phv_data_381 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  phv_data_382 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  phv_data_383 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  phv_data_384 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  phv_data_385 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  phv_data_386 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  phv_data_387 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  phv_data_388 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  phv_data_389 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  phv_data_390 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  phv_data_391 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  phv_data_392 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  phv_data_393 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  phv_data_394 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  phv_data_395 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  phv_data_396 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  phv_data_397 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  phv_data_398 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  phv_data_399 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  phv_data_400 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  phv_data_401 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  phv_data_402 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  phv_data_403 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  phv_data_404 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  phv_data_405 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  phv_data_406 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  phv_data_407 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  phv_data_408 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  phv_data_409 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  phv_data_410 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  phv_data_411 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  phv_data_412 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  phv_data_413 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  phv_data_414 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  phv_data_415 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  phv_data_416 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  phv_data_417 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  phv_data_418 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  phv_data_419 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  phv_data_420 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  phv_data_421 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  phv_data_422 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  phv_data_423 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  phv_data_424 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  phv_data_425 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  phv_data_426 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  phv_data_427 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  phv_data_428 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  phv_data_429 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  phv_data_430 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  phv_data_431 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  phv_data_432 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  phv_data_433 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  phv_data_434 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  phv_data_435 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  phv_data_436 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  phv_data_437 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  phv_data_438 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  phv_data_439 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  phv_data_440 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  phv_data_441 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  phv_data_442 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  phv_data_443 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  phv_data_444 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  phv_data_445 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  phv_data_446 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  phv_data_447 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  phv_data_448 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  phv_data_449 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  phv_data_450 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  phv_data_451 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  phv_data_452 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  phv_data_453 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  phv_data_454 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  phv_data_455 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  phv_data_456 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  phv_data_457 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  phv_data_458 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  phv_data_459 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  phv_data_460 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  phv_data_461 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  phv_data_462 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  phv_data_463 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  phv_data_464 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  phv_data_465 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  phv_data_466 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  phv_data_467 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  phv_data_468 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  phv_data_469 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  phv_data_470 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  phv_data_471 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  phv_data_472 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  phv_data_473 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  phv_data_474 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  phv_data_475 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  phv_data_476 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  phv_data_477 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  phv_data_478 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  phv_data_479 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  phv_data_480 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  phv_data_481 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  phv_data_482 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  phv_data_483 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  phv_data_484 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  phv_data_485 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  phv_data_486 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  phv_data_487 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  phv_data_488 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  phv_data_489 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  phv_data_490 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  phv_data_491 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  phv_data_492 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  phv_data_493 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  phv_data_494 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  phv_data_495 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  phv_data_496 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  phv_data_497 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  phv_data_498 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  phv_data_499 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  phv_data_500 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  phv_data_501 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  phv_data_502 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  phv_data_503 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  phv_data_504 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  phv_data_505 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  phv_data_506 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  phv_data_507 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  phv_data_508 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  phv_data_509 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  phv_data_510 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  phv_data_511 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  phv_header_0 = _RAND_512[15:0];
  _RAND_513 = {1{`RANDOM}};
  phv_header_1 = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  phv_header_2 = _RAND_514[15:0];
  _RAND_515 = {1{`RANDOM}};
  phv_header_3 = _RAND_515[15:0];
  _RAND_516 = {1{`RANDOM}};
  phv_header_4 = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  phv_header_5 = _RAND_517[15:0];
  _RAND_518 = {1{`RANDOM}};
  phv_header_6 = _RAND_518[15:0];
  _RAND_519 = {1{`RANDOM}};
  phv_header_7 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  phv_header_8 = _RAND_520[15:0];
  _RAND_521 = {1{`RANDOM}};
  phv_header_9 = _RAND_521[15:0];
  _RAND_522 = {1{`RANDOM}};
  phv_header_10 = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  phv_header_11 = _RAND_523[15:0];
  _RAND_524 = {1{`RANDOM}};
  phv_header_12 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  phv_header_13 = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  phv_header_14 = _RAND_526[15:0];
  _RAND_527 = {1{`RANDOM}};
  phv_header_15 = _RAND_527[15:0];
  _RAND_528 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_530[15:0];
  _RAND_531 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  phv_next_config_id = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  key_offset = _RAND_534[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
