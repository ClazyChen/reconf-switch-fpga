module Matcher(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [2:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [2:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_config_id,
  input  [7:0]  io_mod_key_mod_header_id,
  input  [7:0]  io_mod_key_mod_internal_offset,
  input  [7:0]  io_mod_key_mod_key_length,
  input  [5:0]  io_mod_table_mod_sram_id_table_0,
  input  [5:0]  io_mod_table_mod_sram_id_table_1,
  input  [5:0]  io_mod_table_mod_sram_id_table_2,
  input  [5:0]  io_mod_table_mod_sram_id_table_3,
  input  [5:0]  io_mod_table_mod_sram_id_table_4,
  input  [5:0]  io_mod_table_mod_sram_id_table_5,
  input  [5:0]  io_mod_table_mod_sram_id_table_6,
  input  [5:0]  io_mod_table_mod_sram_id_table_7,
  input  [5:0]  io_mod_table_mod_sram_id_table_8,
  input  [5:0]  io_mod_table_mod_sram_id_table_9,
  input  [5:0]  io_mod_table_mod_sram_id_table_10,
  input  [5:0]  io_mod_table_mod_sram_id_table_11,
  input  [5:0]  io_mod_table_mod_sram_id_table_12,
  input  [5:0]  io_mod_table_mod_sram_id_table_13,
  input  [5:0]  io_mod_table_mod_sram_id_table_14,
  input  [5:0]  io_mod_table_mod_sram_id_table_15,
  input  [5:0]  io_mod_table_mod_sram_id_table_16,
  input  [5:0]  io_mod_table_mod_sram_id_table_17,
  input  [5:0]  io_mod_table_mod_sram_id_table_18,
  input  [5:0]  io_mod_table_mod_sram_id_table_19,
  input  [5:0]  io_mod_table_mod_sram_id_table_20,
  input  [5:0]  io_mod_table_mod_sram_id_table_21,
  input  [5:0]  io_mod_table_mod_sram_id_table_22,
  input  [5:0]  io_mod_table_mod_sram_id_table_23,
  input  [5:0]  io_mod_table_mod_sram_id_table_24,
  input  [5:0]  io_mod_table_mod_sram_id_table_25,
  input  [5:0]  io_mod_table_mod_sram_id_table_26,
  input  [5:0]  io_mod_table_mod_sram_id_table_27,
  input  [5:0]  io_mod_table_mod_sram_id_table_28,
  input  [5:0]  io_mod_table_mod_sram_id_table_29,
  input  [5:0]  io_mod_table_mod_sram_id_table_30,
  input  [5:0]  io_mod_table_mod_sram_id_table_31,
  input  [5:0]  io_mod_table_mod_sram_id_table_32,
  input  [5:0]  io_mod_table_mod_sram_id_table_33,
  input  [5:0]  io_mod_table_mod_sram_id_table_34,
  input  [5:0]  io_mod_table_mod_sram_id_table_35,
  input  [5:0]  io_mod_table_mod_sram_id_table_36,
  input  [5:0]  io_mod_table_mod_sram_id_table_37,
  input  [5:0]  io_mod_table_mod_sram_id_table_38,
  input  [5:0]  io_mod_table_mod_sram_id_table_39,
  input  [5:0]  io_mod_table_mod_sram_id_table_40,
  input  [5:0]  io_mod_table_mod_sram_id_table_41,
  input  [5:0]  io_mod_table_mod_sram_id_table_42,
  input  [5:0]  io_mod_table_mod_sram_id_table_43,
  input  [5:0]  io_mod_table_mod_sram_id_table_44,
  input  [5:0]  io_mod_table_mod_sram_id_table_45,
  input  [5:0]  io_mod_table_mod_sram_id_table_46,
  input  [5:0]  io_mod_table_mod_sram_id_table_47,
  input  [5:0]  io_mod_table_mod_sram_id_table_48,
  input  [5:0]  io_mod_table_mod_sram_id_table_49,
  input  [5:0]  io_mod_table_mod_sram_id_table_50,
  input  [5:0]  io_mod_table_mod_sram_id_table_51,
  input  [5:0]  io_mod_table_mod_sram_id_table_52,
  input  [5:0]  io_mod_table_mod_sram_id_table_53,
  input  [5:0]  io_mod_table_mod_sram_id_table_54,
  input  [5:0]  io_mod_table_mod_sram_id_table_55,
  input  [5:0]  io_mod_table_mod_sram_id_table_56,
  input  [5:0]  io_mod_table_mod_sram_id_table_57,
  input  [5:0]  io_mod_table_mod_sram_id_table_58,
  input  [5:0]  io_mod_table_mod_sram_id_table_59,
  input  [5:0]  io_mod_table_mod_sram_id_table_60,
  input  [5:0]  io_mod_table_mod_sram_id_table_61,
  input  [5:0]  io_mod_table_mod_sram_id_table_62,
  input  [5:0]  io_mod_table_mod_sram_id_table_63,
  input  [6:0]  io_mod_table_mod_table_width,
  input  [6:0]  io_mod_table_mod_table_depth,
  output        io_hit,
  output [63:0] io_match_value,
  output        io_mem_cluster_0_en,
  output [7:0]  io_mem_cluster_0_addr,
  input  [63:0] io_mem_cluster_0_data,
  output        io_mem_cluster_1_en,
  output [7:0]  io_mem_cluster_1_addr,
  input  [63:0] io_mem_cluster_1_data,
  output        io_mem_cluster_2_en,
  output [7:0]  io_mem_cluster_2_addr,
  input  [63:0] io_mem_cluster_2_data,
  output        io_mem_cluster_3_en,
  output [7:0]  io_mem_cluster_3_addr,
  input  [63:0] io_mem_cluster_3_data,
  output        io_mem_cluster_4_en,
  output [7:0]  io_mem_cluster_4_addr,
  input  [63:0] io_mem_cluster_4_data,
  output        io_mem_cluster_5_en,
  output [7:0]  io_mem_cluster_5_addr,
  input  [63:0] io_mem_cluster_5_data,
  output        io_mem_cluster_6_en,
  output [7:0]  io_mem_cluster_6_addr,
  input  [63:0] io_mem_cluster_6_data,
  output        io_mem_cluster_7_en,
  output [7:0]  io_mem_cluster_7_addr,
  input  [63:0] io_mem_cluster_7_data,
  output        io_mem_cluster_8_en,
  output [7:0]  io_mem_cluster_8_addr,
  input  [63:0] io_mem_cluster_8_data,
  output        io_mem_cluster_9_en,
  output [7:0]  io_mem_cluster_9_addr,
  input  [63:0] io_mem_cluster_9_data,
  output        io_mem_cluster_10_en,
  output [7:0]  io_mem_cluster_10_addr,
  input  [63:0] io_mem_cluster_10_data,
  output        io_mem_cluster_11_en,
  output [7:0]  io_mem_cluster_11_addr,
  input  [63:0] io_mem_cluster_11_data,
  output        io_mem_cluster_12_en,
  output [7:0]  io_mem_cluster_12_addr,
  input  [63:0] io_mem_cluster_12_data,
  output        io_mem_cluster_13_en,
  output [7:0]  io_mem_cluster_13_addr,
  input  [63:0] io_mem_cluster_13_data,
  output        io_mem_cluster_14_en,
  output [7:0]  io_mem_cluster_14_addr,
  input  [63:0] io_mem_cluster_14_data,
  output        io_mem_cluster_15_en,
  output [7:0]  io_mem_cluster_15_addr,
  input  [63:0] io_mem_cluster_15_data,
  output        io_mem_cluster_16_en,
  output [7:0]  io_mem_cluster_16_addr,
  input  [63:0] io_mem_cluster_16_data,
  output        io_mem_cluster_17_en,
  output [7:0]  io_mem_cluster_17_addr,
  input  [63:0] io_mem_cluster_17_data,
  output        io_mem_cluster_18_en,
  output [7:0]  io_mem_cluster_18_addr,
  input  [63:0] io_mem_cluster_18_data,
  output        io_mem_cluster_19_en,
  output [7:0]  io_mem_cluster_19_addr,
  input  [63:0] io_mem_cluster_19_data,
  output        io_mem_cluster_20_en,
  output [7:0]  io_mem_cluster_20_addr,
  input  [63:0] io_mem_cluster_20_data,
  output        io_mem_cluster_21_en,
  output [7:0]  io_mem_cluster_21_addr,
  input  [63:0] io_mem_cluster_21_data,
  output        io_mem_cluster_22_en,
  output [7:0]  io_mem_cluster_22_addr,
  input  [63:0] io_mem_cluster_22_data,
  output        io_mem_cluster_23_en,
  output [7:0]  io_mem_cluster_23_addr,
  input  [63:0] io_mem_cluster_23_data,
  output        io_mem_cluster_24_en,
  output [7:0]  io_mem_cluster_24_addr,
  input  [63:0] io_mem_cluster_24_data,
  output        io_mem_cluster_25_en,
  output [7:0]  io_mem_cluster_25_addr,
  input  [63:0] io_mem_cluster_25_data,
  output        io_mem_cluster_26_en,
  output [7:0]  io_mem_cluster_26_addr,
  input  [63:0] io_mem_cluster_26_data,
  output        io_mem_cluster_27_en,
  output [7:0]  io_mem_cluster_27_addr,
  input  [63:0] io_mem_cluster_27_data,
  output        io_mem_cluster_28_en,
  output [7:0]  io_mem_cluster_28_addr,
  input  [63:0] io_mem_cluster_28_data,
  output        io_mem_cluster_29_en,
  output [7:0]  io_mem_cluster_29_addr,
  input  [63:0] io_mem_cluster_29_data,
  output        io_mem_cluster_30_en,
  output [7:0]  io_mem_cluster_30_addr,
  input  [63:0] io_mem_cluster_30_data,
  output        io_mem_cluster_31_en,
  output [7:0]  io_mem_cluster_31_addr,
  input  [63:0] io_mem_cluster_31_data,
  output        io_mem_cluster_32_en,
  output [7:0]  io_mem_cluster_32_addr,
  input  [63:0] io_mem_cluster_32_data,
  output        io_mem_cluster_33_en,
  output [7:0]  io_mem_cluster_33_addr,
  input  [63:0] io_mem_cluster_33_data,
  output        io_mem_cluster_34_en,
  output [7:0]  io_mem_cluster_34_addr,
  input  [63:0] io_mem_cluster_34_data,
  output        io_mem_cluster_35_en,
  output [7:0]  io_mem_cluster_35_addr,
  input  [63:0] io_mem_cluster_35_data,
  output        io_mem_cluster_36_en,
  output [7:0]  io_mem_cluster_36_addr,
  input  [63:0] io_mem_cluster_36_data,
  output        io_mem_cluster_37_en,
  output [7:0]  io_mem_cluster_37_addr,
  input  [63:0] io_mem_cluster_37_data,
  output        io_mem_cluster_38_en,
  output [7:0]  io_mem_cluster_38_addr,
  input  [63:0] io_mem_cluster_38_data,
  output        io_mem_cluster_39_en,
  output [7:0]  io_mem_cluster_39_addr,
  input  [63:0] io_mem_cluster_39_data,
  output        io_mem_cluster_40_en,
  output [7:0]  io_mem_cluster_40_addr,
  input  [63:0] io_mem_cluster_40_data,
  output        io_mem_cluster_41_en,
  output [7:0]  io_mem_cluster_41_addr,
  input  [63:0] io_mem_cluster_41_data,
  output        io_mem_cluster_42_en,
  output [7:0]  io_mem_cluster_42_addr,
  input  [63:0] io_mem_cluster_42_data,
  output        io_mem_cluster_43_en,
  output [7:0]  io_mem_cluster_43_addr,
  input  [63:0] io_mem_cluster_43_data,
  output        io_mem_cluster_44_en,
  output [7:0]  io_mem_cluster_44_addr,
  input  [63:0] io_mem_cluster_44_data,
  output        io_mem_cluster_45_en,
  output [7:0]  io_mem_cluster_45_addr,
  input  [63:0] io_mem_cluster_45_data,
  output        io_mem_cluster_46_en,
  output [7:0]  io_mem_cluster_46_addr,
  input  [63:0] io_mem_cluster_46_data,
  output        io_mem_cluster_47_en,
  output [7:0]  io_mem_cluster_47_addr,
  input  [63:0] io_mem_cluster_47_data,
  output        io_mem_cluster_48_en,
  output [7:0]  io_mem_cluster_48_addr,
  input  [63:0] io_mem_cluster_48_data,
  output        io_mem_cluster_49_en,
  output [7:0]  io_mem_cluster_49_addr,
  input  [63:0] io_mem_cluster_49_data,
  output        io_mem_cluster_50_en,
  output [7:0]  io_mem_cluster_50_addr,
  input  [63:0] io_mem_cluster_50_data,
  output        io_mem_cluster_51_en,
  output [7:0]  io_mem_cluster_51_addr,
  input  [63:0] io_mem_cluster_51_data,
  output        io_mem_cluster_52_en,
  output [7:0]  io_mem_cluster_52_addr,
  input  [63:0] io_mem_cluster_52_data,
  output        io_mem_cluster_53_en,
  output [7:0]  io_mem_cluster_53_addr,
  input  [63:0] io_mem_cluster_53_data,
  output        io_mem_cluster_54_en,
  output [7:0]  io_mem_cluster_54_addr,
  input  [63:0] io_mem_cluster_54_data,
  output        io_mem_cluster_55_en,
  output [7:0]  io_mem_cluster_55_addr,
  input  [63:0] io_mem_cluster_55_data,
  output        io_mem_cluster_56_en,
  output [7:0]  io_mem_cluster_56_addr,
  input  [63:0] io_mem_cluster_56_data,
  output        io_mem_cluster_57_en,
  output [7:0]  io_mem_cluster_57_addr,
  input  [63:0] io_mem_cluster_57_data,
  output        io_mem_cluster_58_en,
  output [7:0]  io_mem_cluster_58_addr,
  input  [63:0] io_mem_cluster_58_data,
  output        io_mem_cluster_59_en,
  output [7:0]  io_mem_cluster_59_addr,
  input  [63:0] io_mem_cluster_59_data,
  output        io_mem_cluster_60_en,
  output [7:0]  io_mem_cluster_60_addr,
  input  [63:0] io_mem_cluster_60_data,
  output        io_mem_cluster_61_en,
  output [7:0]  io_mem_cluster_61_addr,
  input  [63:0] io_mem_cluster_61_data,
  output        io_mem_cluster_62_en,
  output [7:0]  io_mem_cluster_62_addr,
  input  [63:0] io_mem_cluster_62_data,
  output        io_mem_cluster_63_en,
  output [7:0]  io_mem_cluster_63_addr,
  input  [63:0] io_mem_cluster_63_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 343:23]
  wire [2:0] pipe1_io_pipe_phv_in_next_processor_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 343:23]
  wire [2:0] pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_0_header_id; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_0_internal_offset; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_1_header_id; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_config_1_internal_offset; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_key_offset; // @[matcher.scala 343:23]
  wire  pipe2_clock; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 344:23]
  wire [2:0] pipe2_io_pipe_phv_in_next_processor_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 344:23]
  wire [2:0] pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_key_config_0_key_length; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_key_config_1_key_length; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_key_offset; // @[matcher.scala 344:23]
  wire [191:0] pipe2_io_match_key; // @[matcher.scala 344:23]
  wire  pipe3to8_clock; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_0; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_1; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_2; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_3; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_4; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_5; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_6; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_7; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_8; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_9; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_10; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_11; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_12; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_13; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_14; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_16; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_17; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_18; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_19; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_20; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_21; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_22; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_23; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_24; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_25; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_26; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_27; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_28; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_29; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_30; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_31; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_32; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_33; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_34; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_35; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_36; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_37; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_38; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_39; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_40; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_41; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_42; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_43; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_44; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_45; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_46; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_47; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_48; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_49; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_50; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_51; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_52; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_53; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_54; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_55; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_56; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_57; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_58; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_59; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_60; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_61; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_62; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_63; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_64; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_65; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_66; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_67; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_68; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_69; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_70; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_71; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_72; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_73; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_74; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_75; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_76; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_77; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_78; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_79; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_80; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_81; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_82; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_83; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_84; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_85; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_86; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_87; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_88; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_89; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_90; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_91; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_92; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_93; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_94; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_95; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_96; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_97; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_98; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_99; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_100; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_101; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_102; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_103; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_104; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_105; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_106; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_107; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_108; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_109; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_110; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_111; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_112; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_113; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_114; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_115; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_116; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_117; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_118; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_119; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_120; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_121; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_122; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_123; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_124; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_125; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_126; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_127; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_128; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_129; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_130; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_131; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_132; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_133; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_134; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_135; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_136; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_137; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_138; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_139; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_140; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_141; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_142; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_143; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_144; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_145; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_146; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_147; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_148; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_149; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_150; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_151; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_152; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_153; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_154; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_155; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_156; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_157; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_158; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_159; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_160; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_161; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_162; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_163; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_164; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_165; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_166; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_167; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_168; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_169; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_170; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_171; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_172; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_173; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_174; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_175; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_176; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_177; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_178; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_179; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_180; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_181; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_182; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_183; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_184; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_185; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_186; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_187; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_188; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_189; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_190; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_191; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_192; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_193; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_194; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_195; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_196; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_197; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_198; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_199; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_200; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_201; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_202; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_203; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_204; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_205; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_206; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_207; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_208; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_209; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_210; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_211; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_212; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_213; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_214; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_215; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_216; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_217; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_218; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_219; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_220; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_221; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_222; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_223; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_224; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_225; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_226; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_227; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_228; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_229; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_230; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_231; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_232; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_233; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_234; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_235; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_236; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_237; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_238; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_239; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_240; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_241; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_242; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_243; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_244; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_245; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_246; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_247; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_248; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_249; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_250; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_251; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_252; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_253; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_254; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_255; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_0; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_1; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_2; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_3; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_4; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_5; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_6; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_7; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_8; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_9; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_10; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_11; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_12; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_13; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_14; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_state; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 345:26]
  wire [2:0] pipe3to8_io_pipe_phv_in_next_processor_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_next_config_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_96; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_97; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_98; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_99; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_100; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_101; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_102; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_103; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_104; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_105; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_106; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_107; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_108; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_109; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_110; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_111; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_112; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_113; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_114; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_115; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_116; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_117; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_118; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_119; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_120; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_121; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_122; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_123; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_124; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_125; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_126; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_127; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_128; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_129; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_130; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_131; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_132; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_133; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_134; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_135; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_136; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_137; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_138; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_139; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_140; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_141; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_142; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_143; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_144; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_145; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_146; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_147; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_148; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_149; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_150; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_151; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_152; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_153; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_154; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_155; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_156; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_157; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_158; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_159; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_160; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_161; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_162; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_163; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_164; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_165; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_166; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_167; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_168; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_169; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_170; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_171; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_172; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_173; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_174; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_175; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_176; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_177; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_178; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_179; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_180; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_181; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_182; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_183; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_184; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_185; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_186; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_187; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_188; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_189; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_190; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_191; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_192; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_193; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_194; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_195; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_196; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_197; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_198; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_199; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_200; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_201; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_202; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_203; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_204; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_205; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_206; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_207; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_208; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_209; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_210; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_211; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_212; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_213; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_214; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_215; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_216; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_217; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_218; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_219; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_220; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_221; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_222; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_223; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_224; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_225; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_226; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_227; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_228; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_229; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_230; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_231; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_232; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_233; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_234; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_235; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_236; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_237; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_238; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_239; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_240; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_241; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_242; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_243; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_244; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_245; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_246; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_247; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_248; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_249; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_250; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_251; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_252; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_253; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_254; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_255; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 345:26]
  wire [2:0] pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 345:26]
  wire  pipe3to8_io_mod_hash_depth_mod; // @[matcher.scala 345:26]
  wire  pipe3to8_io_mod_config_id; // @[matcher.scala 345:26]
  wire [5:0] pipe3to8_io_mod_hash_depth; // @[matcher.scala 345:26]
  wire [191:0] pipe3to8_io_key_in; // @[matcher.scala 345:26]
  wire [191:0] pipe3to8_io_key_out; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_hash_val; // @[matcher.scala 345:26]
  wire [5:0] pipe3to8_io_hash_val_cs; // @[matcher.scala 345:26]
  wire  pipe9_clock; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_0; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_1; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_2; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_3; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_4; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_5; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_6; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_7; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_8; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_9; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_10; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_11; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_12; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_13; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_14; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_16; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_17; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_18; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_19; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_20; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_21; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_22; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_23; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_24; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_25; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_26; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_27; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_28; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_29; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_30; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_31; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_32; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_33; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_34; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_35; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_36; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_37; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_38; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_39; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_40; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_41; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_42; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_43; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_44; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_45; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_46; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_47; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_48; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_49; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_50; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_51; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_52; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_53; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_54; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_55; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_56; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_57; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_58; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_59; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_60; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_61; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_62; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_63; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_64; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_65; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_66; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_67; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_68; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_69; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_70; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_71; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_72; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_73; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_74; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_75; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_76; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_77; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_78; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_79; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_80; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_81; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_82; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_83; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_84; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_85; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_86; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_87; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_88; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_89; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_90; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_91; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_92; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_93; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_94; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_95; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_96; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_97; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_98; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_99; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_100; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_101; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_102; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_103; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_104; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_105; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_106; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_107; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_108; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_109; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_110; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_111; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_112; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_113; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_114; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_115; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_116; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_117; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_118; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_119; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_120; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_121; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_122; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_123; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_124; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_125; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_126; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_127; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_128; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_129; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_130; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_131; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_132; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_133; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_134; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_135; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_136; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_137; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_138; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_139; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_140; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_141; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_142; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_143; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_144; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_145; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_146; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_147; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_148; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_149; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_150; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_151; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_152; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_153; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_154; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_155; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_156; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_157; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_158; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_159; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_160; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_161; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_162; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_163; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_164; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_165; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_166; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_167; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_168; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_169; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_170; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_171; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_172; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_173; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_174; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_175; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_176; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_177; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_178; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_179; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_180; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_181; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_182; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_183; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_184; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_185; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_186; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_187; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_188; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_189; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_190; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_191; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_192; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_193; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_194; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_195; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_196; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_197; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_198; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_199; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_200; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_201; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_202; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_203; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_204; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_205; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_206; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_207; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_208; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_209; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_210; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_211; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_212; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_213; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_214; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_215; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_216; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_217; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_218; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_219; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_220; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_221; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_222; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_223; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_224; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_225; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_226; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_227; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_228; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_229; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_230; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_231; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_232; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_233; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_234; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_235; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_236; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_237; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_238; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_239; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_240; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_241; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_242; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_243; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_244; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_245; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_246; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_247; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_248; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_249; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_250; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_251; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_252; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_253; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_254; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_255; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_0; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_1; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_2; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_3; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_4; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_5; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_6; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_7; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_8; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_9; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_10; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_11; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_12; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_13; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_14; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_state; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 346:23]
  wire [2:0] pipe9_io_pipe_phv_in_next_processor_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_next_config_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_96; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_97; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_98; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_99; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_100; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_101; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_102; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_103; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_104; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_105; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_106; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_107; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_108; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_109; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_110; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_111; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_112; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_113; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_114; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_115; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_116; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_117; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_118; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_119; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_120; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_121; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_122; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_123; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_124; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_125; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_126; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_127; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_128; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_129; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_130; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_131; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_132; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_133; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_134; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_135; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_136; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_137; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_138; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_139; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_140; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_141; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_142; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_143; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_144; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_145; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_146; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_147; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_148; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_149; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_150; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_151; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_152; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_153; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_154; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_155; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_156; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_157; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_158; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_159; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_160; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_161; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_162; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_163; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_164; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_165; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_166; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_167; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_168; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_169; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_170; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_171; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_172; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_173; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_174; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_175; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_176; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_177; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_178; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_179; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_180; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_181; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_182; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_183; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_184; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_185; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_186; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_187; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_188; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_189; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_190; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_191; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_192; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_193; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_194; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_195; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_196; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_197; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_198; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_199; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_200; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_201; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_202; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_203; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_204; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_205; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_206; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_207; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_208; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_209; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_210; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_211; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_212; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_213; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_214; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_215; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_216; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_217; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_218; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_219; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_220; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_221; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_222; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_223; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_224; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_225; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_226; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_227; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_228; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_229; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_230; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_231; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_232; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_233; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_234; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_235; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_236; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_237; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_238; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_239; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_240; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_241; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_242; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_243; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_244; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_245; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_246; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_247; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_248; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_249; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_250; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_251; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_252; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_253; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_254; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_255; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 346:23]
  wire [2:0] pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_0; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_1; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_2; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_3; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_4; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_5; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_6; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_7; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_8; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_9; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_10; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_11; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_12; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_13; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_14; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_15; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_16; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_17; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_18; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_19; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_20; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_21; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_22; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_23; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_24; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_25; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_26; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_27; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_28; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_29; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_30; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_31; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_32; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_33; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_34; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_35; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_36; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_37; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_38; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_39; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_40; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_41; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_42; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_43; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_44; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_45; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_46; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_47; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_48; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_49; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_50; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_51; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_52; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_53; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_54; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_55; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_56; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_57; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_58; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_59; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_60; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_61; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_62; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_0_sram_id_table_63; // @[matcher.scala 346:23]
  wire [6:0] pipe9_io_table_config_0_table_width; // @[matcher.scala 346:23]
  wire [6:0] pipe9_io_table_config_0_table_depth; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_0; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_1; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_2; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_3; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_4; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_5; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_6; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_7; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_8; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_9; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_10; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_11; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_12; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_13; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_14; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_15; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_16; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_17; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_18; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_19; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_20; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_21; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_22; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_23; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_24; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_25; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_26; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_27; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_28; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_29; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_30; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_31; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_32; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_33; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_34; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_35; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_36; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_37; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_38; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_39; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_40; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_41; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_42; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_43; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_44; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_45; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_46; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_47; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_48; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_49; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_50; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_51; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_52; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_53; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_54; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_55; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_56; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_57; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_58; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_59; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_60; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_61; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_62; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_table_config_1_sram_id_table_63; // @[matcher.scala 346:23]
  wire [6:0] pipe9_io_table_config_1_table_width; // @[matcher.scala 346:23]
  wire [6:0] pipe9_io_table_config_1_table_depth; // @[matcher.scala 346:23]
  wire [191:0] pipe9_io_key_in; // @[matcher.scala 346:23]
  wire [191:0] pipe9_io_key_out; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_addr_in; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_addr_out; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_cs_in; // @[matcher.scala 346:23]
  wire [5:0] pipe9_io_cs_out; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_0; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_1; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_2; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_3; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_4; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_5; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_6; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_7; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_8; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_9; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_10; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_11; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_12; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_13; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_14; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_15; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_16; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_17; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_18; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_19; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_20; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_21; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_22; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_23; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_24; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_25; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_26; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_27; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_28; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_29; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_30; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_31; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_32; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_33; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_34; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_35; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_36; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_37; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_38; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_39; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_40; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_41; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_42; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_43; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_44; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_45; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_46; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_47; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_48; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_49; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_50; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_51; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_52; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_53; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_54; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_55; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_56; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_57; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_58; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_59; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_60; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_61; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_62; // @[matcher.scala 346:23]
  wire  pipe9_io_cs_vec_out_63; // @[matcher.scala 346:23]
  wire  pipe10_clock; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_0; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_1; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_2; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_3; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_4; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_5; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_6; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_7; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_8; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_9; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_10; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_11; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_12; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_13; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_14; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_16; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_17; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_18; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_19; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_20; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_21; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_22; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_23; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_24; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_25; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_26; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_27; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_28; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_29; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_30; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_31; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_32; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_33; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_34; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_35; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_36; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_37; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_38; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_39; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_40; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_41; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_42; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_43; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_44; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_45; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_46; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_47; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_48; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_49; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_50; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_51; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_52; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_53; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_54; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_55; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_56; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_57; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_58; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_59; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_60; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_61; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_62; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_63; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_64; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_65; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_66; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_67; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_68; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_69; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_70; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_71; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_72; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_73; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_74; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_75; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_76; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_77; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_78; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_79; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_80; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_81; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_82; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_83; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_84; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_85; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_86; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_87; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_88; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_89; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_90; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_91; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_92; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_93; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_94; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_95; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_96; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_97; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_98; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_99; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_100; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_101; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_102; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_103; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_104; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_105; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_106; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_107; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_108; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_109; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_110; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_111; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_112; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_113; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_114; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_115; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_116; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_117; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_118; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_119; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_120; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_121; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_122; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_123; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_124; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_125; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_126; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_127; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_128; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_129; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_130; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_131; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_132; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_133; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_134; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_135; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_136; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_137; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_138; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_139; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_140; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_141; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_142; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_143; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_144; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_145; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_146; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_147; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_148; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_149; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_150; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_151; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_152; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_153; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_154; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_155; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_156; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_157; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_158; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_159; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_160; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_161; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_162; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_163; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_164; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_165; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_166; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_167; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_168; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_169; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_170; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_171; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_172; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_173; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_174; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_175; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_176; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_177; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_178; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_179; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_180; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_181; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_182; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_183; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_184; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_185; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_186; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_187; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_188; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_189; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_190; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_191; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_192; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_193; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_194; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_195; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_196; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_197; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_198; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_199; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_200; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_201; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_202; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_203; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_204; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_205; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_206; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_207; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_208; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_209; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_210; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_211; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_212; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_213; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_214; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_215; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_216; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_217; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_218; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_219; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_220; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_221; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_222; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_223; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_224; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_225; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_226; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_227; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_228; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_229; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_230; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_231; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_232; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_233; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_234; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_235; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_236; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_237; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_238; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_239; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_240; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_241; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_242; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_243; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_244; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_245; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_246; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_247; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_248; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_249; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_250; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_251; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_252; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_253; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_254; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_255; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_0; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_1; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_2; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_3; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_4; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_5; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_6; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_7; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_8; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_9; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_10; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_11; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_12; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_13; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_14; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_state; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 347:24]
  wire [2:0] pipe10_io_pipe_phv_in_next_processor_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_next_config_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_96; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_97; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_98; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_99; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_100; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_101; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_102; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_103; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_104; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_105; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_106; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_107; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_108; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_109; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_110; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_111; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_112; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_113; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_114; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_115; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_116; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_117; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_118; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_119; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_120; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_121; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_122; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_123; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_124; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_125; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_126; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_127; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_128; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_129; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_130; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_131; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_132; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_133; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_134; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_135; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_136; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_137; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_138; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_139; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_140; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_141; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_142; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_143; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_144; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_145; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_146; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_147; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_148; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_149; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_150; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_151; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_152; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_153; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_154; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_155; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_156; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_157; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_158; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_159; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_160; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_161; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_162; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_163; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_164; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_165; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_166; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_167; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_168; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_169; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_170; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_171; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_172; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_173; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_174; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_175; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_176; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_177; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_178; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_179; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_180; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_181; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_182; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_183; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_184; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_185; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_186; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_187; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_188; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_189; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_190; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_191; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_192; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_193; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_194; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_195; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_196; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_197; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_198; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_199; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_200; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_201; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_202; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_203; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_204; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_205; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_206; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_207; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_208; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_209; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_210; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_211; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_212; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_213; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_214; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_215; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_216; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_217; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_218; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_219; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_220; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_221; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_222; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_223; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_224; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_225; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_226; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_227; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_228; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_229; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_230; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_231; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_232; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_233; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_234; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_235; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_236; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_237; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_238; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_239; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_240; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_241; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_242; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_243; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_244; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_245; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_246; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_247; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_248; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_249; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_250; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_251; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_252; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_253; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_254; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_255; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 347:24]
  wire [2:0] pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 347:24]
  wire [191:0] pipe10_io_key_in; // @[matcher.scala 347:24]
  wire [191:0] pipe10_io_key_out; // @[matcher.scala 347:24]
  wire [5:0] pipe10_io_cs_in; // @[matcher.scala 347:24]
  wire [5:0] pipe10_io_cs_out; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_addr_in; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_0; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_1; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_2; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_3; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_4; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_5; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_6; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_7; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_8; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_9; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_10; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_11; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_12; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_13; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_14; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_15; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_16; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_17; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_18; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_19; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_20; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_21; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_22; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_23; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_24; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_25; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_26; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_27; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_28; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_29; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_30; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_31; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_32; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_33; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_34; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_35; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_36; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_37; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_38; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_39; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_40; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_41; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_42; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_43; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_44; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_45; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_46; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_47; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_48; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_49; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_50; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_51; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_52; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_53; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_54; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_55; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_56; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_57; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_58; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_59; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_60; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_61; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_62; // @[matcher.scala 347:24]
  wire  pipe10_io_cs_vec_in_63; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_0; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_1; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_2; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_3; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_4; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_5; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_6; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_7; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_8; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_9; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_10; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_11; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_12; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_13; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_14; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_15; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_16; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_17; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_18; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_19; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_20; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_21; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_22; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_23; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_24; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_25; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_26; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_27; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_28; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_29; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_30; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_31; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_32; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_33; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_34; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_35; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_36; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_37; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_38; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_39; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_40; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_41; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_42; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_43; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_44; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_45; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_46; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_47; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_48; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_49; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_50; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_51; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_52; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_53; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_54; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_55; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_56; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_57; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_58; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_59; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_60; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_61; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_62; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_data_out_63; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_0_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_0_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_0_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_1_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_1_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_1_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_2_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_2_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_2_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_3_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_3_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_3_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_4_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_4_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_4_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_5_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_5_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_5_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_6_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_6_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_6_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_7_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_7_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_7_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_8_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_8_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_8_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_9_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_9_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_9_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_10_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_10_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_10_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_11_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_11_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_11_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_12_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_12_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_12_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_13_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_13_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_13_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_14_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_14_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_14_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_15_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_15_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_15_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_16_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_16_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_16_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_17_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_17_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_17_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_18_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_18_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_18_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_19_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_19_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_19_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_20_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_20_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_20_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_21_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_21_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_21_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_22_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_22_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_22_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_23_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_23_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_23_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_24_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_24_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_24_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_25_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_25_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_25_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_26_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_26_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_26_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_27_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_27_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_27_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_28_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_28_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_28_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_29_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_29_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_29_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_30_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_30_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_30_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_31_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_31_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_31_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_32_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_32_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_32_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_33_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_33_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_33_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_34_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_34_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_34_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_35_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_35_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_35_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_36_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_36_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_36_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_37_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_37_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_37_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_38_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_38_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_38_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_39_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_39_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_39_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_40_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_40_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_40_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_41_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_41_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_41_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_42_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_42_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_42_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_43_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_43_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_43_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_44_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_44_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_44_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_45_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_45_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_45_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_46_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_46_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_46_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_47_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_47_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_47_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_48_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_48_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_48_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_49_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_49_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_49_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_50_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_50_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_50_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_51_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_51_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_51_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_52_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_52_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_52_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_53_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_53_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_53_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_54_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_54_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_54_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_55_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_55_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_55_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_56_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_56_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_56_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_57_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_57_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_57_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_58_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_58_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_58_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_59_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_59_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_59_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_60_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_60_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_60_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_61_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_61_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_61_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_62_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_62_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_62_data; // @[matcher.scala 347:24]
  wire  pipe10_io_mem_cluster_63_en; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_mem_cluster_63_addr; // @[matcher.scala 347:24]
  wire [63:0] pipe10_io_mem_cluster_63_data; // @[matcher.scala 347:24]
  wire  pipe11_clock; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_0; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_1; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_2; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_3; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_4; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_5; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_6; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_7; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_8; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_9; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_10; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_11; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_12; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_13; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_14; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_16; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_17; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_18; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_19; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_20; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_21; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_22; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_23; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_24; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_25; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_26; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_27; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_28; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_29; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_30; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_31; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_32; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_33; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_34; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_35; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_36; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_37; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_38; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_39; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_40; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_41; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_42; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_43; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_44; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_45; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_46; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_47; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_48; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_49; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_50; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_51; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_52; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_53; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_54; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_55; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_56; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_57; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_58; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_59; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_60; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_61; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_62; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_63; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_64; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_65; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_66; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_67; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_68; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_69; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_70; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_71; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_72; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_73; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_74; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_75; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_76; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_77; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_78; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_79; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_80; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_81; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_82; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_83; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_84; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_85; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_86; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_87; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_88; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_89; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_90; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_91; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_92; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_93; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_94; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_95; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_96; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_97; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_98; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_99; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_100; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_101; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_102; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_103; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_104; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_105; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_106; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_107; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_108; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_109; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_110; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_111; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_112; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_113; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_114; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_115; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_116; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_117; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_118; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_119; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_120; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_121; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_122; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_123; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_124; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_125; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_126; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_127; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_128; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_129; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_130; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_131; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_132; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_133; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_134; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_135; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_136; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_137; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_138; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_139; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_140; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_141; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_142; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_143; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_144; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_145; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_146; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_147; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_148; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_149; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_150; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_151; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_152; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_153; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_154; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_155; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_156; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_157; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_158; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_159; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_160; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_161; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_162; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_163; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_164; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_165; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_166; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_167; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_168; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_169; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_170; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_171; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_172; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_173; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_174; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_175; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_176; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_177; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_178; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_179; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_180; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_181; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_182; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_183; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_184; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_185; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_186; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_187; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_188; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_189; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_190; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_191; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_192; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_193; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_194; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_195; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_196; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_197; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_198; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_199; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_200; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_201; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_202; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_203; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_204; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_205; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_206; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_207; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_208; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_209; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_210; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_211; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_212; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_213; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_214; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_215; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_216; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_217; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_218; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_219; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_220; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_221; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_222; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_223; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_224; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_225; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_226; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_227; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_228; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_229; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_230; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_231; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_232; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_233; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_234; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_235; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_236; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_237; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_238; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_239; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_240; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_241; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_242; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_243; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_244; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_245; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_246; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_247; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_248; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_249; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_250; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_251; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_252; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_253; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_254; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_255; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_0; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_1; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_2; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_3; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_4; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_5; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_6; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_7; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_8; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_9; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_10; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_11; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_12; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_13; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_14; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_state; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 348:24]
  wire [2:0] pipe11_io_pipe_phv_in_next_processor_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_next_config_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_96; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_97; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_98; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_99; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_100; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_101; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_102; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_103; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_104; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_105; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_106; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_107; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_108; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_109; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_110; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_111; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_112; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_113; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_114; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_115; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_116; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_117; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_118; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_119; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_120; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_121; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_122; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_123; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_124; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_125; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_126; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_127; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_128; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_129; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_130; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_131; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_132; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_133; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_134; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_135; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_136; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_137; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_138; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_139; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_140; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_141; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_142; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_143; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_144; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_145; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_146; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_147; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_148; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_149; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_150; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_151; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_152; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_153; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_154; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_155; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_156; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_157; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_158; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_159; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_160; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_161; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_162; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_163; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_164; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_165; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_166; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_167; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_168; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_169; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_170; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_171; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_172; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_173; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_174; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_175; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_176; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_177; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_178; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_179; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_180; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_181; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_182; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_183; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_184; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_185; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_186; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_187; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_188; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_189; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_190; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_191; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_192; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_193; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_194; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_195; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_196; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_197; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_198; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_199; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_200; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_201; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_202; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_203; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_204; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_205; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_206; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_207; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_208; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_209; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_210; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_211; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_212; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_213; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_214; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_215; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_216; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_217; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_218; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_219; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_220; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_221; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_222; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_223; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_224; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_225; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_226; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_227; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_228; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_229; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_230; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_231; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_232; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_233; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_234; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_235; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_236; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_237; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_238; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_239; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_240; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_241; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_242; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_243; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_244; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_245; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_246; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_247; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_248; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_249; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_250; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_251; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_252; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_253; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_254; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_255; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 348:24]
  wire [2:0] pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 348:24]
  wire [6:0] pipe11_io_table_config_0_table_width; // @[matcher.scala 348:24]
  wire [6:0] pipe11_io_table_config_0_table_depth; // @[matcher.scala 348:24]
  wire [6:0] pipe11_io_table_config_1_table_width; // @[matcher.scala 348:24]
  wire [6:0] pipe11_io_table_config_1_table_depth; // @[matcher.scala 348:24]
  wire [191:0] pipe11_io_key_in; // @[matcher.scala 348:24]
  wire [191:0] pipe11_io_key_out; // @[matcher.scala 348:24]
  wire [5:0] pipe11_io_cs_in; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_0; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_1; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_2; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_3; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_4; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_5; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_6; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_7; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_8; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_9; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_10; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_11; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_12; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_13; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_14; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_15; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_16; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_17; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_18; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_19; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_20; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_21; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_22; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_23; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_24; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_25; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_26; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_27; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_28; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_29; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_30; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_31; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_32; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_33; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_34; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_35; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_36; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_37; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_38; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_39; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_40; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_41; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_42; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_43; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_44; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_45; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_46; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_47; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_48; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_49; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_50; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_51; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_52; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_53; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_54; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_55; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_56; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_57; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_58; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_59; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_60; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_61; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_62; // @[matcher.scala 348:24]
  wire [63:0] pipe11_io_data_in_63; // @[matcher.scala 348:24]
  wire [255:0] pipe11_io_data_out; // @[matcher.scala 348:24]
  wire  pipe12_clock; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_0; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_1; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_2; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_3; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_4; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_5; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_6; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_7; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_8; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_9; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_10; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_11; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_12; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_13; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_14; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_16; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_17; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_18; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_19; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_20; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_21; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_22; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_23; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_24; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_25; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_26; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_27; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_28; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_29; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_30; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_31; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_32; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_33; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_34; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_35; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_36; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_37; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_38; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_39; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_40; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_41; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_42; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_43; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_44; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_45; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_46; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_47; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_48; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_49; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_50; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_51; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_52; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_53; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_54; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_55; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_56; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_57; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_58; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_59; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_60; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_61; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_62; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_63; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_64; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_65; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_66; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_67; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_68; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_69; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_70; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_71; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_72; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_73; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_74; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_75; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_76; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_77; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_78; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_79; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_80; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_81; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_82; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_83; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_84; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_85; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_86; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_87; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_88; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_89; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_90; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_91; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_92; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_93; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_94; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_95; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_96; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_97; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_98; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_99; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_100; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_101; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_102; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_103; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_104; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_105; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_106; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_107; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_108; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_109; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_110; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_111; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_112; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_113; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_114; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_115; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_116; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_117; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_118; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_119; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_120; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_121; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_122; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_123; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_124; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_125; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_126; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_127; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_128; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_129; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_130; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_131; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_132; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_133; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_134; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_135; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_136; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_137; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_138; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_139; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_140; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_141; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_142; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_143; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_144; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_145; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_146; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_147; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_148; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_149; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_150; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_151; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_152; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_153; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_154; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_155; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_156; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_157; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_158; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_159; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_160; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_161; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_162; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_163; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_164; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_165; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_166; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_167; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_168; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_169; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_170; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_171; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_172; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_173; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_174; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_175; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_176; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_177; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_178; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_179; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_180; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_181; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_182; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_183; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_184; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_185; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_186; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_187; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_188; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_189; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_190; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_191; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_192; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_193; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_194; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_195; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_196; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_197; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_198; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_199; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_200; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_201; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_202; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_203; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_204; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_205; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_206; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_207; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_208; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_209; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_210; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_211; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_212; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_213; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_214; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_215; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_216; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_217; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_218; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_219; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_220; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_221; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_222; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_223; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_224; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_225; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_226; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_227; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_228; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_229; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_230; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_231; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_232; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_233; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_234; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_235; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_236; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_237; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_238; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_239; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_240; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_241; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_242; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_243; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_244; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_245; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_246; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_247; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_248; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_249; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_250; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_251; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_252; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_253; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_254; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_255; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_0; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_1; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_2; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_3; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_4; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_5; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_6; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_7; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_8; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_9; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_10; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_11; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_12; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_13; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_14; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_state; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 349:24]
  wire [2:0] pipe12_io_pipe_phv_in_next_processor_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_next_config_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_96; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_97; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_98; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_99; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_100; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_101; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_102; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_103; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_104; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_105; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_106; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_107; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_108; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_109; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_110; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_111; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_112; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_113; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_114; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_115; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_116; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_117; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_118; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_119; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_120; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_121; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_122; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_123; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_124; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_125; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_126; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_127; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_128; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_129; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_130; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_131; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_132; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_133; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_134; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_135; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_136; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_137; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_138; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_139; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_140; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_141; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_142; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_143; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_144; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_145; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_146; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_147; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_148; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_149; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_150; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_151; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_152; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_153; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_154; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_155; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_156; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_157; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_158; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_159; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_160; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_161; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_162; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_163; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_164; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_165; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_166; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_167; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_168; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_169; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_170; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_171; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_172; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_173; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_174; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_175; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_176; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_177; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_178; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_179; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_180; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_181; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_182; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_183; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_184; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_185; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_186; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_187; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_188; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_189; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_190; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_191; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_192; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_193; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_194; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_195; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_196; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_197; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_198; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_199; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_200; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_201; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_202; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_203; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_204; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_205; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_206; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_207; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_208; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_209; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_210; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_211; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_212; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_213; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_214; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_215; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_216; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_217; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_218; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_219; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_220; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_221; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_222; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_223; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_224; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_225; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_226; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_227; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_228; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_229; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_230; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_231; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_232; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_233; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_234; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_235; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_236; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_237; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_238; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_239; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_240; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_241; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_242; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_243; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_244; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_245; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_246; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_247; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_248; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_249; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_250; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_251; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_252; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_253; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_254; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_255; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 349:24]
  wire [2:0] pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_key_config_0_key_length; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_key_config_1_key_length; // @[matcher.scala 349:24]
  wire [191:0] pipe12_io_key_in; // @[matcher.scala 349:24]
  wire [255:0] pipe12_io_data_in; // @[matcher.scala 349:24]
  wire  pipe12_io_hit; // @[matcher.scala 349:24]
  wire [63:0] pipe12_io_match_value; // @[matcher.scala 349:24]
  reg [7:0] key_config_0_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_0_internal_offset; // @[matcher.scala 17:25]
  reg [7:0] key_config_0_key_length; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_header_id; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_internal_offset; // @[matcher.scala 17:25]
  reg [7:0] key_config_1_key_length; // @[matcher.scala 17:25]
  reg [5:0] table_config_0_sram_id_table_0; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_1; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_2; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_3; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_4; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_5; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_6; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_7; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_8; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_9; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_10; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_11; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_12; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_13; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_14; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_15; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_16; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_17; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_18; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_19; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_20; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_21; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_22; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_23; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_24; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_25; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_26; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_27; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_28; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_29; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_30; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_31; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_32; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_33; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_34; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_35; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_36; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_37; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_38; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_39; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_40; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_41; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_42; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_43; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_44; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_45; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_46; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_47; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_48; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_49; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_50; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_51; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_52; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_53; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_54; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_55; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_56; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_57; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_58; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_59; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_60; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_61; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_62; // @[matcher.scala 18:27]
  reg [5:0] table_config_0_sram_id_table_63; // @[matcher.scala 18:27]
  reg [6:0] table_config_0_table_width; // @[matcher.scala 18:27]
  reg [6:0] table_config_0_table_depth; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_0; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_1; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_2; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_3; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_4; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_5; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_6; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_7; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_8; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_9; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_10; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_11; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_12; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_13; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_14; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_15; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_16; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_17; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_18; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_19; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_20; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_21; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_22; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_23; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_24; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_25; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_26; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_27; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_28; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_29; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_30; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_31; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_32; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_33; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_34; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_35; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_36; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_37; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_38; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_39; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_40; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_41; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_42; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_43; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_44; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_45; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_46; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_47; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_48; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_49; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_50; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_51; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_52; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_53; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_54; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_55; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_56; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_57; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_58; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_59; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_60; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_61; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_62; // @[matcher.scala 18:27]
  reg [5:0] table_config_1_sram_id_table_63; // @[matcher.scala 18:27]
  reg [6:0] table_config_1_table_width; // @[matcher.scala 18:27]
  reg [6:0] table_config_1_table_depth; // @[matcher.scala 18:27]
  MatchGetOffset pipe1 ( // @[matcher.scala 343:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_header_id(pipe1_io_key_config_0_header_id),
    .io_key_config_0_internal_offset(pipe1_io_key_config_0_internal_offset),
    .io_key_config_1_header_id(pipe1_io_key_config_1_header_id),
    .io_key_config_1_internal_offset(pipe1_io_key_config_1_internal_offset),
    .io_key_offset(pipe1_io_key_offset)
  );
  MatchGetKey pipe2 ( // @[matcher.scala 344:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe2_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe2_io_key_config_1_key_length),
    .io_key_offset(pipe2_io_key_offset),
    .io_match_key(pipe2_io_match_key)
  );
  Hash pipe3to8 ( // @[matcher.scala 345:26]
    .clock(pipe3to8_clock),
    .io_pipe_phv_in_data_0(pipe3to8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3to8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3to8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3to8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3to8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3to8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3to8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3to8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3to8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3to8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3to8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3to8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3to8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3to8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3to8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3to8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3to8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3to8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3to8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3to8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3to8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3to8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3to8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3to8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3to8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3to8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3to8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3to8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3to8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3to8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3to8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3to8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3to8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3to8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3to8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3to8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3to8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3to8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3to8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3to8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3to8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3to8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3to8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3to8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3to8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3to8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3to8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3to8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3to8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3to8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3to8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3to8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3to8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3to8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3to8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3to8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3to8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3to8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3to8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3to8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3to8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3to8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3to8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3to8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3to8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3to8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3to8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3to8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3to8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3to8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3to8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3to8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3to8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3to8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3to8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3to8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3to8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3to8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3to8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3to8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3to8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3to8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3to8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3to8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3to8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3to8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3to8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3to8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3to8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3to8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3to8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3to8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3to8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3to8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3to8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3to8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3to8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3to8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3to8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3to8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3to8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3to8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3to8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3to8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3to8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3to8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3to8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3to8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3to8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3to8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3to8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3to8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3to8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3to8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3to8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3to8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3to8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3to8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3to8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3to8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3to8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3to8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3to8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3to8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3to8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3to8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3to8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3to8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3to8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3to8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3to8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3to8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3to8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3to8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3to8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3to8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3to8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3to8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3to8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3to8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3to8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3to8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3to8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3to8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3to8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3to8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3to8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3to8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3to8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3to8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3to8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3to8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3to8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3to8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3to8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3to8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3to8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3to8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3to8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3to8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3to8_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3to8_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3to8_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3to8_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3to8_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3to8_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3to8_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3to8_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3to8_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3to8_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3to8_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3to8_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3to8_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3to8_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3to8_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3to8_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3to8_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3to8_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3to8_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3to8_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3to8_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3to8_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3to8_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3to8_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3to8_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3to8_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3to8_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3to8_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3to8_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3to8_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3to8_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3to8_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3to8_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3to8_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3to8_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3to8_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3to8_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3to8_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3to8_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3to8_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3to8_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3to8_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3to8_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3to8_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3to8_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3to8_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3to8_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3to8_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3to8_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3to8_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3to8_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3to8_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3to8_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3to8_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3to8_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3to8_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3to8_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3to8_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3to8_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3to8_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3to8_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3to8_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3to8_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3to8_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3to8_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3to8_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3to8_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3to8_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3to8_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3to8_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3to8_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3to8_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3to8_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3to8_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3to8_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3to8_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3to8_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3to8_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3to8_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3to8_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3to8_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3to8_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3to8_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3to8_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3to8_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3to8_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3to8_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3to8_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3to8_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3to8_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3to8_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3to8_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3to8_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3to8_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3to8_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3to8_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe3to8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3to8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3to8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3to8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3to8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3to8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3to8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3to8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3to8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3to8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3to8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3to8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3to8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3to8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3to8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3to8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3to8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3to8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3to8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3to8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3to8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3to8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3to8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3to8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3to8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3to8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3to8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3to8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3to8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3to8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3to8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3to8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3to8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3to8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3to8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3to8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3to8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3to8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3to8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3to8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3to8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3to8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3to8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3to8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3to8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3to8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3to8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3to8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3to8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3to8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3to8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3to8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3to8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3to8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3to8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3to8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3to8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3to8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3to8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3to8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3to8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3to8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3to8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3to8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3to8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3to8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3to8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3to8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3to8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3to8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3to8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3to8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3to8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3to8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3to8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3to8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3to8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3to8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3to8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3to8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3to8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3to8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3to8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3to8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3to8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3to8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3to8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3to8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3to8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3to8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3to8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3to8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3to8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3to8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3to8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3to8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3to8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3to8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3to8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3to8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3to8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3to8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3to8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3to8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3to8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3to8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3to8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3to8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3to8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3to8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3to8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3to8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3to8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3to8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3to8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3to8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3to8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3to8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3to8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3to8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3to8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3to8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3to8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3to8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3to8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3to8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3to8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3to8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3to8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3to8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3to8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3to8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3to8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3to8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3to8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3to8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3to8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3to8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3to8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3to8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3to8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3to8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3to8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3to8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3to8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3to8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3to8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3to8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3to8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3to8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3to8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3to8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3to8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3to8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3to8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3to8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3to8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3to8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3to8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3to8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3to8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3to8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3to8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3to8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3to8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3to8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3to8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3to8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3to8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3to8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3to8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3to8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3to8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3to8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3to8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3to8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3to8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3to8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3to8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3to8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3to8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3to8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3to8_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3to8_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3to8_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3to8_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3to8_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3to8_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3to8_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3to8_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3to8_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3to8_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3to8_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3to8_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3to8_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3to8_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3to8_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3to8_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3to8_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3to8_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3to8_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3to8_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3to8_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3to8_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3to8_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3to8_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3to8_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3to8_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3to8_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3to8_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3to8_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3to8_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3to8_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3to8_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3to8_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3to8_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3to8_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3to8_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3to8_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3to8_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3to8_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3to8_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3to8_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3to8_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3to8_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3to8_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3to8_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3to8_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3to8_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3to8_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3to8_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3to8_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3to8_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3to8_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3to8_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3to8_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3to8_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3to8_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3to8_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3to8_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3to8_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3to8_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3to8_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3to8_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3to8_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3to8_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3to8_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3to8_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3to8_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3to8_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3to8_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3to8_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3to8_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3to8_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3to8_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3to8_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3to8_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3to8_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3to8_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3to8_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3to8_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3to8_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3to8_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3to8_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3to8_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3to8_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3to8_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3to8_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3to8_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3to8_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3to8_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3to8_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3to8_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3to8_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3to8_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3to8_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3to8_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3to8_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe3to8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3to8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3to8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3to8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3to8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3to8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3to8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3to8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3to8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3to8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3to8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3to8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3to8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3to8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3to8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3to8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3to8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3to8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3to8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3to8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3to8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3to8_io_pipe_phv_out_is_valid_processor),
    .io_mod_hash_depth_mod(pipe3to8_io_mod_hash_depth_mod),
    .io_mod_config_id(pipe3to8_io_mod_config_id),
    .io_mod_hash_depth(pipe3to8_io_mod_hash_depth),
    .io_key_in(pipe3to8_io_key_in),
    .io_key_out(pipe3to8_io_key_out),
    .io_hash_val(pipe3to8_io_hash_val),
    .io_hash_val_cs(pipe3to8_io_hash_val_cs)
  );
  MatchGetCs pipe9 ( // @[matcher.scala 346:23]
    .clock(pipe9_clock),
    .io_pipe_phv_in_data_0(pipe9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe9_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe9_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe9_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe9_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe9_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe9_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe9_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe9_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe9_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe9_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe9_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe9_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe9_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe9_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe9_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe9_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe9_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe9_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe9_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe9_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe9_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe9_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe9_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe9_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe9_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe9_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe9_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe9_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe9_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe9_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe9_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe9_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe9_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe9_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe9_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe9_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe9_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe9_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe9_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe9_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe9_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe9_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe9_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe9_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe9_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe9_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe9_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe9_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe9_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe9_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe9_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe9_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe9_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe9_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe9_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe9_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe9_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe9_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe9_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe9_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe9_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe9_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe9_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe9_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe9_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe9_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe9_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe9_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe9_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe9_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe9_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe9_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe9_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe9_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe9_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe9_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe9_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe9_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe9_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe9_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe9_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe9_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe9_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe9_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe9_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe9_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe9_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe9_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe9_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe9_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe9_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe9_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe9_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe9_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe9_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe9_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe9_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe9_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe9_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe9_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe9_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe9_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe9_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe9_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe9_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe9_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe9_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe9_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe9_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe9_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe9_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe9_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe9_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe9_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe9_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe9_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe9_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe9_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe9_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe9_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe9_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe9_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe9_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe9_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe9_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe9_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe9_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe9_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe9_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe9_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe9_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe9_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe9_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe9_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe9_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe9_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe9_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe9_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe9_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe9_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe9_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe9_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe9_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe9_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe9_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe9_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe9_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe9_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe9_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe9_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe9_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe9_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe9_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe9_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe9_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe9_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe9_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe9_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe9_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe9_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe9_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe9_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe9_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe9_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe9_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe9_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe9_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe9_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe9_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe9_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe9_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe9_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe9_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe9_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe9_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe9_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe9_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe9_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe9_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe9_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe9_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe9_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe9_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe9_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe9_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe9_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe9_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe9_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe9_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe9_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe9_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe9_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe9_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe9_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe9_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe9_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe9_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe9_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe9_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe9_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe9_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe9_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe9_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe9_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe9_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe9_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe9_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe9_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe9_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe9_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe9_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe9_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe9_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe9_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe9_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe9_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe9_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe9_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe9_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe9_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe9_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe9_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe9_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe9_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe9_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe9_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe9_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe9_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe9_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe9_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe9_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe9_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe9_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe9_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe9_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe9_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe9_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe9_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe9_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe9_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe9_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe9_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe9_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe9_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe9_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe9_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe9_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe9_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe9_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe9_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe9_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe9_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe9_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe9_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe9_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe9_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe9_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe9_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe9_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe9_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe9_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe9_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe9_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe9_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe9_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe9_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe9_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe9_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe9_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe9_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe9_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe9_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe9_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe9_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe9_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe9_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe9_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe9_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe9_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe9_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe9_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe9_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe9_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe9_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe9_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe9_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe9_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe9_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe9_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe9_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe9_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe9_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe9_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe9_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe9_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe9_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe9_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe9_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe9_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe9_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe9_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe9_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe9_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe9_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe9_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe9_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe9_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe9_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe9_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe9_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe9_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe9_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe9_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe9_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe9_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe9_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe9_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe9_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe9_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe9_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe9_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe9_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe9_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe9_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe9_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe9_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe9_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe9_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe9_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe9_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe9_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe9_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe9_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe9_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe9_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe9_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe9_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe9_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe9_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe9_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe9_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe9_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe9_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe9_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe9_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe9_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe9_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe9_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe9_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe9_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe9_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe9_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe9_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe9_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe9_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe9_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe9_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe9_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe9_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_sram_id_table_0(pipe9_io_table_config_0_sram_id_table_0),
    .io_table_config_0_sram_id_table_1(pipe9_io_table_config_0_sram_id_table_1),
    .io_table_config_0_sram_id_table_2(pipe9_io_table_config_0_sram_id_table_2),
    .io_table_config_0_sram_id_table_3(pipe9_io_table_config_0_sram_id_table_3),
    .io_table_config_0_sram_id_table_4(pipe9_io_table_config_0_sram_id_table_4),
    .io_table_config_0_sram_id_table_5(pipe9_io_table_config_0_sram_id_table_5),
    .io_table_config_0_sram_id_table_6(pipe9_io_table_config_0_sram_id_table_6),
    .io_table_config_0_sram_id_table_7(pipe9_io_table_config_0_sram_id_table_7),
    .io_table_config_0_sram_id_table_8(pipe9_io_table_config_0_sram_id_table_8),
    .io_table_config_0_sram_id_table_9(pipe9_io_table_config_0_sram_id_table_9),
    .io_table_config_0_sram_id_table_10(pipe9_io_table_config_0_sram_id_table_10),
    .io_table_config_0_sram_id_table_11(pipe9_io_table_config_0_sram_id_table_11),
    .io_table_config_0_sram_id_table_12(pipe9_io_table_config_0_sram_id_table_12),
    .io_table_config_0_sram_id_table_13(pipe9_io_table_config_0_sram_id_table_13),
    .io_table_config_0_sram_id_table_14(pipe9_io_table_config_0_sram_id_table_14),
    .io_table_config_0_sram_id_table_15(pipe9_io_table_config_0_sram_id_table_15),
    .io_table_config_0_sram_id_table_16(pipe9_io_table_config_0_sram_id_table_16),
    .io_table_config_0_sram_id_table_17(pipe9_io_table_config_0_sram_id_table_17),
    .io_table_config_0_sram_id_table_18(pipe9_io_table_config_0_sram_id_table_18),
    .io_table_config_0_sram_id_table_19(pipe9_io_table_config_0_sram_id_table_19),
    .io_table_config_0_sram_id_table_20(pipe9_io_table_config_0_sram_id_table_20),
    .io_table_config_0_sram_id_table_21(pipe9_io_table_config_0_sram_id_table_21),
    .io_table_config_0_sram_id_table_22(pipe9_io_table_config_0_sram_id_table_22),
    .io_table_config_0_sram_id_table_23(pipe9_io_table_config_0_sram_id_table_23),
    .io_table_config_0_sram_id_table_24(pipe9_io_table_config_0_sram_id_table_24),
    .io_table_config_0_sram_id_table_25(pipe9_io_table_config_0_sram_id_table_25),
    .io_table_config_0_sram_id_table_26(pipe9_io_table_config_0_sram_id_table_26),
    .io_table_config_0_sram_id_table_27(pipe9_io_table_config_0_sram_id_table_27),
    .io_table_config_0_sram_id_table_28(pipe9_io_table_config_0_sram_id_table_28),
    .io_table_config_0_sram_id_table_29(pipe9_io_table_config_0_sram_id_table_29),
    .io_table_config_0_sram_id_table_30(pipe9_io_table_config_0_sram_id_table_30),
    .io_table_config_0_sram_id_table_31(pipe9_io_table_config_0_sram_id_table_31),
    .io_table_config_0_sram_id_table_32(pipe9_io_table_config_0_sram_id_table_32),
    .io_table_config_0_sram_id_table_33(pipe9_io_table_config_0_sram_id_table_33),
    .io_table_config_0_sram_id_table_34(pipe9_io_table_config_0_sram_id_table_34),
    .io_table_config_0_sram_id_table_35(pipe9_io_table_config_0_sram_id_table_35),
    .io_table_config_0_sram_id_table_36(pipe9_io_table_config_0_sram_id_table_36),
    .io_table_config_0_sram_id_table_37(pipe9_io_table_config_0_sram_id_table_37),
    .io_table_config_0_sram_id_table_38(pipe9_io_table_config_0_sram_id_table_38),
    .io_table_config_0_sram_id_table_39(pipe9_io_table_config_0_sram_id_table_39),
    .io_table_config_0_sram_id_table_40(pipe9_io_table_config_0_sram_id_table_40),
    .io_table_config_0_sram_id_table_41(pipe9_io_table_config_0_sram_id_table_41),
    .io_table_config_0_sram_id_table_42(pipe9_io_table_config_0_sram_id_table_42),
    .io_table_config_0_sram_id_table_43(pipe9_io_table_config_0_sram_id_table_43),
    .io_table_config_0_sram_id_table_44(pipe9_io_table_config_0_sram_id_table_44),
    .io_table_config_0_sram_id_table_45(pipe9_io_table_config_0_sram_id_table_45),
    .io_table_config_0_sram_id_table_46(pipe9_io_table_config_0_sram_id_table_46),
    .io_table_config_0_sram_id_table_47(pipe9_io_table_config_0_sram_id_table_47),
    .io_table_config_0_sram_id_table_48(pipe9_io_table_config_0_sram_id_table_48),
    .io_table_config_0_sram_id_table_49(pipe9_io_table_config_0_sram_id_table_49),
    .io_table_config_0_sram_id_table_50(pipe9_io_table_config_0_sram_id_table_50),
    .io_table_config_0_sram_id_table_51(pipe9_io_table_config_0_sram_id_table_51),
    .io_table_config_0_sram_id_table_52(pipe9_io_table_config_0_sram_id_table_52),
    .io_table_config_0_sram_id_table_53(pipe9_io_table_config_0_sram_id_table_53),
    .io_table_config_0_sram_id_table_54(pipe9_io_table_config_0_sram_id_table_54),
    .io_table_config_0_sram_id_table_55(pipe9_io_table_config_0_sram_id_table_55),
    .io_table_config_0_sram_id_table_56(pipe9_io_table_config_0_sram_id_table_56),
    .io_table_config_0_sram_id_table_57(pipe9_io_table_config_0_sram_id_table_57),
    .io_table_config_0_sram_id_table_58(pipe9_io_table_config_0_sram_id_table_58),
    .io_table_config_0_sram_id_table_59(pipe9_io_table_config_0_sram_id_table_59),
    .io_table_config_0_sram_id_table_60(pipe9_io_table_config_0_sram_id_table_60),
    .io_table_config_0_sram_id_table_61(pipe9_io_table_config_0_sram_id_table_61),
    .io_table_config_0_sram_id_table_62(pipe9_io_table_config_0_sram_id_table_62),
    .io_table_config_0_sram_id_table_63(pipe9_io_table_config_0_sram_id_table_63),
    .io_table_config_0_table_width(pipe9_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe9_io_table_config_0_table_depth),
    .io_table_config_1_sram_id_table_0(pipe9_io_table_config_1_sram_id_table_0),
    .io_table_config_1_sram_id_table_1(pipe9_io_table_config_1_sram_id_table_1),
    .io_table_config_1_sram_id_table_2(pipe9_io_table_config_1_sram_id_table_2),
    .io_table_config_1_sram_id_table_3(pipe9_io_table_config_1_sram_id_table_3),
    .io_table_config_1_sram_id_table_4(pipe9_io_table_config_1_sram_id_table_4),
    .io_table_config_1_sram_id_table_5(pipe9_io_table_config_1_sram_id_table_5),
    .io_table_config_1_sram_id_table_6(pipe9_io_table_config_1_sram_id_table_6),
    .io_table_config_1_sram_id_table_7(pipe9_io_table_config_1_sram_id_table_7),
    .io_table_config_1_sram_id_table_8(pipe9_io_table_config_1_sram_id_table_8),
    .io_table_config_1_sram_id_table_9(pipe9_io_table_config_1_sram_id_table_9),
    .io_table_config_1_sram_id_table_10(pipe9_io_table_config_1_sram_id_table_10),
    .io_table_config_1_sram_id_table_11(pipe9_io_table_config_1_sram_id_table_11),
    .io_table_config_1_sram_id_table_12(pipe9_io_table_config_1_sram_id_table_12),
    .io_table_config_1_sram_id_table_13(pipe9_io_table_config_1_sram_id_table_13),
    .io_table_config_1_sram_id_table_14(pipe9_io_table_config_1_sram_id_table_14),
    .io_table_config_1_sram_id_table_15(pipe9_io_table_config_1_sram_id_table_15),
    .io_table_config_1_sram_id_table_16(pipe9_io_table_config_1_sram_id_table_16),
    .io_table_config_1_sram_id_table_17(pipe9_io_table_config_1_sram_id_table_17),
    .io_table_config_1_sram_id_table_18(pipe9_io_table_config_1_sram_id_table_18),
    .io_table_config_1_sram_id_table_19(pipe9_io_table_config_1_sram_id_table_19),
    .io_table_config_1_sram_id_table_20(pipe9_io_table_config_1_sram_id_table_20),
    .io_table_config_1_sram_id_table_21(pipe9_io_table_config_1_sram_id_table_21),
    .io_table_config_1_sram_id_table_22(pipe9_io_table_config_1_sram_id_table_22),
    .io_table_config_1_sram_id_table_23(pipe9_io_table_config_1_sram_id_table_23),
    .io_table_config_1_sram_id_table_24(pipe9_io_table_config_1_sram_id_table_24),
    .io_table_config_1_sram_id_table_25(pipe9_io_table_config_1_sram_id_table_25),
    .io_table_config_1_sram_id_table_26(pipe9_io_table_config_1_sram_id_table_26),
    .io_table_config_1_sram_id_table_27(pipe9_io_table_config_1_sram_id_table_27),
    .io_table_config_1_sram_id_table_28(pipe9_io_table_config_1_sram_id_table_28),
    .io_table_config_1_sram_id_table_29(pipe9_io_table_config_1_sram_id_table_29),
    .io_table_config_1_sram_id_table_30(pipe9_io_table_config_1_sram_id_table_30),
    .io_table_config_1_sram_id_table_31(pipe9_io_table_config_1_sram_id_table_31),
    .io_table_config_1_sram_id_table_32(pipe9_io_table_config_1_sram_id_table_32),
    .io_table_config_1_sram_id_table_33(pipe9_io_table_config_1_sram_id_table_33),
    .io_table_config_1_sram_id_table_34(pipe9_io_table_config_1_sram_id_table_34),
    .io_table_config_1_sram_id_table_35(pipe9_io_table_config_1_sram_id_table_35),
    .io_table_config_1_sram_id_table_36(pipe9_io_table_config_1_sram_id_table_36),
    .io_table_config_1_sram_id_table_37(pipe9_io_table_config_1_sram_id_table_37),
    .io_table_config_1_sram_id_table_38(pipe9_io_table_config_1_sram_id_table_38),
    .io_table_config_1_sram_id_table_39(pipe9_io_table_config_1_sram_id_table_39),
    .io_table_config_1_sram_id_table_40(pipe9_io_table_config_1_sram_id_table_40),
    .io_table_config_1_sram_id_table_41(pipe9_io_table_config_1_sram_id_table_41),
    .io_table_config_1_sram_id_table_42(pipe9_io_table_config_1_sram_id_table_42),
    .io_table_config_1_sram_id_table_43(pipe9_io_table_config_1_sram_id_table_43),
    .io_table_config_1_sram_id_table_44(pipe9_io_table_config_1_sram_id_table_44),
    .io_table_config_1_sram_id_table_45(pipe9_io_table_config_1_sram_id_table_45),
    .io_table_config_1_sram_id_table_46(pipe9_io_table_config_1_sram_id_table_46),
    .io_table_config_1_sram_id_table_47(pipe9_io_table_config_1_sram_id_table_47),
    .io_table_config_1_sram_id_table_48(pipe9_io_table_config_1_sram_id_table_48),
    .io_table_config_1_sram_id_table_49(pipe9_io_table_config_1_sram_id_table_49),
    .io_table_config_1_sram_id_table_50(pipe9_io_table_config_1_sram_id_table_50),
    .io_table_config_1_sram_id_table_51(pipe9_io_table_config_1_sram_id_table_51),
    .io_table_config_1_sram_id_table_52(pipe9_io_table_config_1_sram_id_table_52),
    .io_table_config_1_sram_id_table_53(pipe9_io_table_config_1_sram_id_table_53),
    .io_table_config_1_sram_id_table_54(pipe9_io_table_config_1_sram_id_table_54),
    .io_table_config_1_sram_id_table_55(pipe9_io_table_config_1_sram_id_table_55),
    .io_table_config_1_sram_id_table_56(pipe9_io_table_config_1_sram_id_table_56),
    .io_table_config_1_sram_id_table_57(pipe9_io_table_config_1_sram_id_table_57),
    .io_table_config_1_sram_id_table_58(pipe9_io_table_config_1_sram_id_table_58),
    .io_table_config_1_sram_id_table_59(pipe9_io_table_config_1_sram_id_table_59),
    .io_table_config_1_sram_id_table_60(pipe9_io_table_config_1_sram_id_table_60),
    .io_table_config_1_sram_id_table_61(pipe9_io_table_config_1_sram_id_table_61),
    .io_table_config_1_sram_id_table_62(pipe9_io_table_config_1_sram_id_table_62),
    .io_table_config_1_sram_id_table_63(pipe9_io_table_config_1_sram_id_table_63),
    .io_table_config_1_table_width(pipe9_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe9_io_table_config_1_table_depth),
    .io_key_in(pipe9_io_key_in),
    .io_key_out(pipe9_io_key_out),
    .io_addr_in(pipe9_io_addr_in),
    .io_addr_out(pipe9_io_addr_out),
    .io_cs_in(pipe9_io_cs_in),
    .io_cs_out(pipe9_io_cs_out),
    .io_cs_vec_out_0(pipe9_io_cs_vec_out_0),
    .io_cs_vec_out_1(pipe9_io_cs_vec_out_1),
    .io_cs_vec_out_2(pipe9_io_cs_vec_out_2),
    .io_cs_vec_out_3(pipe9_io_cs_vec_out_3),
    .io_cs_vec_out_4(pipe9_io_cs_vec_out_4),
    .io_cs_vec_out_5(pipe9_io_cs_vec_out_5),
    .io_cs_vec_out_6(pipe9_io_cs_vec_out_6),
    .io_cs_vec_out_7(pipe9_io_cs_vec_out_7),
    .io_cs_vec_out_8(pipe9_io_cs_vec_out_8),
    .io_cs_vec_out_9(pipe9_io_cs_vec_out_9),
    .io_cs_vec_out_10(pipe9_io_cs_vec_out_10),
    .io_cs_vec_out_11(pipe9_io_cs_vec_out_11),
    .io_cs_vec_out_12(pipe9_io_cs_vec_out_12),
    .io_cs_vec_out_13(pipe9_io_cs_vec_out_13),
    .io_cs_vec_out_14(pipe9_io_cs_vec_out_14),
    .io_cs_vec_out_15(pipe9_io_cs_vec_out_15),
    .io_cs_vec_out_16(pipe9_io_cs_vec_out_16),
    .io_cs_vec_out_17(pipe9_io_cs_vec_out_17),
    .io_cs_vec_out_18(pipe9_io_cs_vec_out_18),
    .io_cs_vec_out_19(pipe9_io_cs_vec_out_19),
    .io_cs_vec_out_20(pipe9_io_cs_vec_out_20),
    .io_cs_vec_out_21(pipe9_io_cs_vec_out_21),
    .io_cs_vec_out_22(pipe9_io_cs_vec_out_22),
    .io_cs_vec_out_23(pipe9_io_cs_vec_out_23),
    .io_cs_vec_out_24(pipe9_io_cs_vec_out_24),
    .io_cs_vec_out_25(pipe9_io_cs_vec_out_25),
    .io_cs_vec_out_26(pipe9_io_cs_vec_out_26),
    .io_cs_vec_out_27(pipe9_io_cs_vec_out_27),
    .io_cs_vec_out_28(pipe9_io_cs_vec_out_28),
    .io_cs_vec_out_29(pipe9_io_cs_vec_out_29),
    .io_cs_vec_out_30(pipe9_io_cs_vec_out_30),
    .io_cs_vec_out_31(pipe9_io_cs_vec_out_31),
    .io_cs_vec_out_32(pipe9_io_cs_vec_out_32),
    .io_cs_vec_out_33(pipe9_io_cs_vec_out_33),
    .io_cs_vec_out_34(pipe9_io_cs_vec_out_34),
    .io_cs_vec_out_35(pipe9_io_cs_vec_out_35),
    .io_cs_vec_out_36(pipe9_io_cs_vec_out_36),
    .io_cs_vec_out_37(pipe9_io_cs_vec_out_37),
    .io_cs_vec_out_38(pipe9_io_cs_vec_out_38),
    .io_cs_vec_out_39(pipe9_io_cs_vec_out_39),
    .io_cs_vec_out_40(pipe9_io_cs_vec_out_40),
    .io_cs_vec_out_41(pipe9_io_cs_vec_out_41),
    .io_cs_vec_out_42(pipe9_io_cs_vec_out_42),
    .io_cs_vec_out_43(pipe9_io_cs_vec_out_43),
    .io_cs_vec_out_44(pipe9_io_cs_vec_out_44),
    .io_cs_vec_out_45(pipe9_io_cs_vec_out_45),
    .io_cs_vec_out_46(pipe9_io_cs_vec_out_46),
    .io_cs_vec_out_47(pipe9_io_cs_vec_out_47),
    .io_cs_vec_out_48(pipe9_io_cs_vec_out_48),
    .io_cs_vec_out_49(pipe9_io_cs_vec_out_49),
    .io_cs_vec_out_50(pipe9_io_cs_vec_out_50),
    .io_cs_vec_out_51(pipe9_io_cs_vec_out_51),
    .io_cs_vec_out_52(pipe9_io_cs_vec_out_52),
    .io_cs_vec_out_53(pipe9_io_cs_vec_out_53),
    .io_cs_vec_out_54(pipe9_io_cs_vec_out_54),
    .io_cs_vec_out_55(pipe9_io_cs_vec_out_55),
    .io_cs_vec_out_56(pipe9_io_cs_vec_out_56),
    .io_cs_vec_out_57(pipe9_io_cs_vec_out_57),
    .io_cs_vec_out_58(pipe9_io_cs_vec_out_58),
    .io_cs_vec_out_59(pipe9_io_cs_vec_out_59),
    .io_cs_vec_out_60(pipe9_io_cs_vec_out_60),
    .io_cs_vec_out_61(pipe9_io_cs_vec_out_61),
    .io_cs_vec_out_62(pipe9_io_cs_vec_out_62),
    .io_cs_vec_out_63(pipe9_io_cs_vec_out_63)
  );
  MatchReadData pipe10 ( // @[matcher.scala 347:24]
    .clock(pipe10_clock),
    .io_pipe_phv_in_data_0(pipe10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe10_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe10_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe10_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe10_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe10_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe10_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe10_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe10_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe10_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe10_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe10_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe10_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe10_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe10_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe10_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe10_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe10_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe10_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe10_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe10_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe10_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe10_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe10_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe10_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe10_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe10_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe10_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe10_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe10_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe10_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe10_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe10_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe10_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe10_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe10_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe10_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe10_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe10_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe10_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe10_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe10_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe10_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe10_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe10_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe10_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe10_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe10_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe10_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe10_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe10_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe10_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe10_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe10_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe10_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe10_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe10_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe10_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe10_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe10_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe10_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe10_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe10_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe10_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe10_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe10_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe10_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe10_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe10_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe10_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe10_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe10_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe10_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe10_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe10_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe10_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe10_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe10_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe10_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe10_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe10_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe10_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe10_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe10_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe10_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe10_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe10_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe10_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe10_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe10_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe10_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe10_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe10_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe10_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe10_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe10_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe10_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe10_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe10_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe10_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe10_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe10_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe10_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe10_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe10_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe10_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe10_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe10_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe10_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe10_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe10_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe10_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe10_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe10_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe10_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe10_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe10_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe10_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe10_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe10_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe10_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe10_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe10_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe10_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe10_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe10_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe10_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe10_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe10_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe10_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe10_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe10_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe10_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe10_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe10_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe10_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe10_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe10_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe10_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe10_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe10_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe10_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe10_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe10_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe10_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe10_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe10_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe10_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe10_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe10_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe10_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe10_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe10_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe10_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe10_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe10_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe10_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe10_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe10_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe10_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe10_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe10_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe10_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe10_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe10_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe10_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe10_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe10_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe10_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe10_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe10_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe10_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe10_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe10_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe10_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe10_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe10_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe10_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe10_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe10_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe10_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe10_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe10_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe10_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe10_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe10_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe10_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe10_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe10_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe10_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe10_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe10_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe10_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe10_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe10_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe10_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe10_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe10_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe10_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe10_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe10_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe10_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe10_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe10_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe10_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe10_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe10_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe10_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe10_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe10_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe10_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe10_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe10_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe10_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe10_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe10_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe10_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe10_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe10_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe10_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe10_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe10_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe10_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe10_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe10_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe10_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe10_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe10_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe10_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe10_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe10_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe10_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe10_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe10_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe10_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe10_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe10_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe10_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe10_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe10_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe10_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe10_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe10_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe10_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe10_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe10_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe10_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe10_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe10_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe10_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe10_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe10_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe10_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe10_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe10_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe10_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe10_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe10_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe10_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe10_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe10_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe10_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe10_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe10_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe10_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe10_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe10_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe10_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe10_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe10_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe10_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe10_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe10_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe10_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe10_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe10_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe10_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe10_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe10_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe10_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe10_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe10_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe10_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe10_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe10_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe10_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe10_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe10_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe10_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe10_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe10_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe10_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe10_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe10_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe10_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe10_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe10_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe10_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe10_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe10_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe10_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe10_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe10_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe10_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe10_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe10_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe10_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe10_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe10_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe10_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe10_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe10_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe10_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe10_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe10_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe10_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe10_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe10_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe10_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe10_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe10_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe10_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe10_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe10_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe10_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe10_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe10_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe10_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe10_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe10_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe10_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe10_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe10_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe10_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe10_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe10_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe10_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe10_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe10_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe10_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe10_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe10_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe10_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe10_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe10_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe10_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe10_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe10_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe10_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe10_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe10_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe10_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe10_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe10_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe10_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe10_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe10_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe10_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe10_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe10_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe10_io_key_in),
    .io_key_out(pipe10_io_key_out),
    .io_cs_in(pipe10_io_cs_in),
    .io_cs_out(pipe10_io_cs_out),
    .io_addr_in(pipe10_io_addr_in),
    .io_cs_vec_in_0(pipe10_io_cs_vec_in_0),
    .io_cs_vec_in_1(pipe10_io_cs_vec_in_1),
    .io_cs_vec_in_2(pipe10_io_cs_vec_in_2),
    .io_cs_vec_in_3(pipe10_io_cs_vec_in_3),
    .io_cs_vec_in_4(pipe10_io_cs_vec_in_4),
    .io_cs_vec_in_5(pipe10_io_cs_vec_in_5),
    .io_cs_vec_in_6(pipe10_io_cs_vec_in_6),
    .io_cs_vec_in_7(pipe10_io_cs_vec_in_7),
    .io_cs_vec_in_8(pipe10_io_cs_vec_in_8),
    .io_cs_vec_in_9(pipe10_io_cs_vec_in_9),
    .io_cs_vec_in_10(pipe10_io_cs_vec_in_10),
    .io_cs_vec_in_11(pipe10_io_cs_vec_in_11),
    .io_cs_vec_in_12(pipe10_io_cs_vec_in_12),
    .io_cs_vec_in_13(pipe10_io_cs_vec_in_13),
    .io_cs_vec_in_14(pipe10_io_cs_vec_in_14),
    .io_cs_vec_in_15(pipe10_io_cs_vec_in_15),
    .io_cs_vec_in_16(pipe10_io_cs_vec_in_16),
    .io_cs_vec_in_17(pipe10_io_cs_vec_in_17),
    .io_cs_vec_in_18(pipe10_io_cs_vec_in_18),
    .io_cs_vec_in_19(pipe10_io_cs_vec_in_19),
    .io_cs_vec_in_20(pipe10_io_cs_vec_in_20),
    .io_cs_vec_in_21(pipe10_io_cs_vec_in_21),
    .io_cs_vec_in_22(pipe10_io_cs_vec_in_22),
    .io_cs_vec_in_23(pipe10_io_cs_vec_in_23),
    .io_cs_vec_in_24(pipe10_io_cs_vec_in_24),
    .io_cs_vec_in_25(pipe10_io_cs_vec_in_25),
    .io_cs_vec_in_26(pipe10_io_cs_vec_in_26),
    .io_cs_vec_in_27(pipe10_io_cs_vec_in_27),
    .io_cs_vec_in_28(pipe10_io_cs_vec_in_28),
    .io_cs_vec_in_29(pipe10_io_cs_vec_in_29),
    .io_cs_vec_in_30(pipe10_io_cs_vec_in_30),
    .io_cs_vec_in_31(pipe10_io_cs_vec_in_31),
    .io_cs_vec_in_32(pipe10_io_cs_vec_in_32),
    .io_cs_vec_in_33(pipe10_io_cs_vec_in_33),
    .io_cs_vec_in_34(pipe10_io_cs_vec_in_34),
    .io_cs_vec_in_35(pipe10_io_cs_vec_in_35),
    .io_cs_vec_in_36(pipe10_io_cs_vec_in_36),
    .io_cs_vec_in_37(pipe10_io_cs_vec_in_37),
    .io_cs_vec_in_38(pipe10_io_cs_vec_in_38),
    .io_cs_vec_in_39(pipe10_io_cs_vec_in_39),
    .io_cs_vec_in_40(pipe10_io_cs_vec_in_40),
    .io_cs_vec_in_41(pipe10_io_cs_vec_in_41),
    .io_cs_vec_in_42(pipe10_io_cs_vec_in_42),
    .io_cs_vec_in_43(pipe10_io_cs_vec_in_43),
    .io_cs_vec_in_44(pipe10_io_cs_vec_in_44),
    .io_cs_vec_in_45(pipe10_io_cs_vec_in_45),
    .io_cs_vec_in_46(pipe10_io_cs_vec_in_46),
    .io_cs_vec_in_47(pipe10_io_cs_vec_in_47),
    .io_cs_vec_in_48(pipe10_io_cs_vec_in_48),
    .io_cs_vec_in_49(pipe10_io_cs_vec_in_49),
    .io_cs_vec_in_50(pipe10_io_cs_vec_in_50),
    .io_cs_vec_in_51(pipe10_io_cs_vec_in_51),
    .io_cs_vec_in_52(pipe10_io_cs_vec_in_52),
    .io_cs_vec_in_53(pipe10_io_cs_vec_in_53),
    .io_cs_vec_in_54(pipe10_io_cs_vec_in_54),
    .io_cs_vec_in_55(pipe10_io_cs_vec_in_55),
    .io_cs_vec_in_56(pipe10_io_cs_vec_in_56),
    .io_cs_vec_in_57(pipe10_io_cs_vec_in_57),
    .io_cs_vec_in_58(pipe10_io_cs_vec_in_58),
    .io_cs_vec_in_59(pipe10_io_cs_vec_in_59),
    .io_cs_vec_in_60(pipe10_io_cs_vec_in_60),
    .io_cs_vec_in_61(pipe10_io_cs_vec_in_61),
    .io_cs_vec_in_62(pipe10_io_cs_vec_in_62),
    .io_cs_vec_in_63(pipe10_io_cs_vec_in_63),
    .io_data_out_0(pipe10_io_data_out_0),
    .io_data_out_1(pipe10_io_data_out_1),
    .io_data_out_2(pipe10_io_data_out_2),
    .io_data_out_3(pipe10_io_data_out_3),
    .io_data_out_4(pipe10_io_data_out_4),
    .io_data_out_5(pipe10_io_data_out_5),
    .io_data_out_6(pipe10_io_data_out_6),
    .io_data_out_7(pipe10_io_data_out_7),
    .io_data_out_8(pipe10_io_data_out_8),
    .io_data_out_9(pipe10_io_data_out_9),
    .io_data_out_10(pipe10_io_data_out_10),
    .io_data_out_11(pipe10_io_data_out_11),
    .io_data_out_12(pipe10_io_data_out_12),
    .io_data_out_13(pipe10_io_data_out_13),
    .io_data_out_14(pipe10_io_data_out_14),
    .io_data_out_15(pipe10_io_data_out_15),
    .io_data_out_16(pipe10_io_data_out_16),
    .io_data_out_17(pipe10_io_data_out_17),
    .io_data_out_18(pipe10_io_data_out_18),
    .io_data_out_19(pipe10_io_data_out_19),
    .io_data_out_20(pipe10_io_data_out_20),
    .io_data_out_21(pipe10_io_data_out_21),
    .io_data_out_22(pipe10_io_data_out_22),
    .io_data_out_23(pipe10_io_data_out_23),
    .io_data_out_24(pipe10_io_data_out_24),
    .io_data_out_25(pipe10_io_data_out_25),
    .io_data_out_26(pipe10_io_data_out_26),
    .io_data_out_27(pipe10_io_data_out_27),
    .io_data_out_28(pipe10_io_data_out_28),
    .io_data_out_29(pipe10_io_data_out_29),
    .io_data_out_30(pipe10_io_data_out_30),
    .io_data_out_31(pipe10_io_data_out_31),
    .io_data_out_32(pipe10_io_data_out_32),
    .io_data_out_33(pipe10_io_data_out_33),
    .io_data_out_34(pipe10_io_data_out_34),
    .io_data_out_35(pipe10_io_data_out_35),
    .io_data_out_36(pipe10_io_data_out_36),
    .io_data_out_37(pipe10_io_data_out_37),
    .io_data_out_38(pipe10_io_data_out_38),
    .io_data_out_39(pipe10_io_data_out_39),
    .io_data_out_40(pipe10_io_data_out_40),
    .io_data_out_41(pipe10_io_data_out_41),
    .io_data_out_42(pipe10_io_data_out_42),
    .io_data_out_43(pipe10_io_data_out_43),
    .io_data_out_44(pipe10_io_data_out_44),
    .io_data_out_45(pipe10_io_data_out_45),
    .io_data_out_46(pipe10_io_data_out_46),
    .io_data_out_47(pipe10_io_data_out_47),
    .io_data_out_48(pipe10_io_data_out_48),
    .io_data_out_49(pipe10_io_data_out_49),
    .io_data_out_50(pipe10_io_data_out_50),
    .io_data_out_51(pipe10_io_data_out_51),
    .io_data_out_52(pipe10_io_data_out_52),
    .io_data_out_53(pipe10_io_data_out_53),
    .io_data_out_54(pipe10_io_data_out_54),
    .io_data_out_55(pipe10_io_data_out_55),
    .io_data_out_56(pipe10_io_data_out_56),
    .io_data_out_57(pipe10_io_data_out_57),
    .io_data_out_58(pipe10_io_data_out_58),
    .io_data_out_59(pipe10_io_data_out_59),
    .io_data_out_60(pipe10_io_data_out_60),
    .io_data_out_61(pipe10_io_data_out_61),
    .io_data_out_62(pipe10_io_data_out_62),
    .io_data_out_63(pipe10_io_data_out_63),
    .io_mem_cluster_0_en(pipe10_io_mem_cluster_0_en),
    .io_mem_cluster_0_addr(pipe10_io_mem_cluster_0_addr),
    .io_mem_cluster_0_data(pipe10_io_mem_cluster_0_data),
    .io_mem_cluster_1_en(pipe10_io_mem_cluster_1_en),
    .io_mem_cluster_1_addr(pipe10_io_mem_cluster_1_addr),
    .io_mem_cluster_1_data(pipe10_io_mem_cluster_1_data),
    .io_mem_cluster_2_en(pipe10_io_mem_cluster_2_en),
    .io_mem_cluster_2_addr(pipe10_io_mem_cluster_2_addr),
    .io_mem_cluster_2_data(pipe10_io_mem_cluster_2_data),
    .io_mem_cluster_3_en(pipe10_io_mem_cluster_3_en),
    .io_mem_cluster_3_addr(pipe10_io_mem_cluster_3_addr),
    .io_mem_cluster_3_data(pipe10_io_mem_cluster_3_data),
    .io_mem_cluster_4_en(pipe10_io_mem_cluster_4_en),
    .io_mem_cluster_4_addr(pipe10_io_mem_cluster_4_addr),
    .io_mem_cluster_4_data(pipe10_io_mem_cluster_4_data),
    .io_mem_cluster_5_en(pipe10_io_mem_cluster_5_en),
    .io_mem_cluster_5_addr(pipe10_io_mem_cluster_5_addr),
    .io_mem_cluster_5_data(pipe10_io_mem_cluster_5_data),
    .io_mem_cluster_6_en(pipe10_io_mem_cluster_6_en),
    .io_mem_cluster_6_addr(pipe10_io_mem_cluster_6_addr),
    .io_mem_cluster_6_data(pipe10_io_mem_cluster_6_data),
    .io_mem_cluster_7_en(pipe10_io_mem_cluster_7_en),
    .io_mem_cluster_7_addr(pipe10_io_mem_cluster_7_addr),
    .io_mem_cluster_7_data(pipe10_io_mem_cluster_7_data),
    .io_mem_cluster_8_en(pipe10_io_mem_cluster_8_en),
    .io_mem_cluster_8_addr(pipe10_io_mem_cluster_8_addr),
    .io_mem_cluster_8_data(pipe10_io_mem_cluster_8_data),
    .io_mem_cluster_9_en(pipe10_io_mem_cluster_9_en),
    .io_mem_cluster_9_addr(pipe10_io_mem_cluster_9_addr),
    .io_mem_cluster_9_data(pipe10_io_mem_cluster_9_data),
    .io_mem_cluster_10_en(pipe10_io_mem_cluster_10_en),
    .io_mem_cluster_10_addr(pipe10_io_mem_cluster_10_addr),
    .io_mem_cluster_10_data(pipe10_io_mem_cluster_10_data),
    .io_mem_cluster_11_en(pipe10_io_mem_cluster_11_en),
    .io_mem_cluster_11_addr(pipe10_io_mem_cluster_11_addr),
    .io_mem_cluster_11_data(pipe10_io_mem_cluster_11_data),
    .io_mem_cluster_12_en(pipe10_io_mem_cluster_12_en),
    .io_mem_cluster_12_addr(pipe10_io_mem_cluster_12_addr),
    .io_mem_cluster_12_data(pipe10_io_mem_cluster_12_data),
    .io_mem_cluster_13_en(pipe10_io_mem_cluster_13_en),
    .io_mem_cluster_13_addr(pipe10_io_mem_cluster_13_addr),
    .io_mem_cluster_13_data(pipe10_io_mem_cluster_13_data),
    .io_mem_cluster_14_en(pipe10_io_mem_cluster_14_en),
    .io_mem_cluster_14_addr(pipe10_io_mem_cluster_14_addr),
    .io_mem_cluster_14_data(pipe10_io_mem_cluster_14_data),
    .io_mem_cluster_15_en(pipe10_io_mem_cluster_15_en),
    .io_mem_cluster_15_addr(pipe10_io_mem_cluster_15_addr),
    .io_mem_cluster_15_data(pipe10_io_mem_cluster_15_data),
    .io_mem_cluster_16_en(pipe10_io_mem_cluster_16_en),
    .io_mem_cluster_16_addr(pipe10_io_mem_cluster_16_addr),
    .io_mem_cluster_16_data(pipe10_io_mem_cluster_16_data),
    .io_mem_cluster_17_en(pipe10_io_mem_cluster_17_en),
    .io_mem_cluster_17_addr(pipe10_io_mem_cluster_17_addr),
    .io_mem_cluster_17_data(pipe10_io_mem_cluster_17_data),
    .io_mem_cluster_18_en(pipe10_io_mem_cluster_18_en),
    .io_mem_cluster_18_addr(pipe10_io_mem_cluster_18_addr),
    .io_mem_cluster_18_data(pipe10_io_mem_cluster_18_data),
    .io_mem_cluster_19_en(pipe10_io_mem_cluster_19_en),
    .io_mem_cluster_19_addr(pipe10_io_mem_cluster_19_addr),
    .io_mem_cluster_19_data(pipe10_io_mem_cluster_19_data),
    .io_mem_cluster_20_en(pipe10_io_mem_cluster_20_en),
    .io_mem_cluster_20_addr(pipe10_io_mem_cluster_20_addr),
    .io_mem_cluster_20_data(pipe10_io_mem_cluster_20_data),
    .io_mem_cluster_21_en(pipe10_io_mem_cluster_21_en),
    .io_mem_cluster_21_addr(pipe10_io_mem_cluster_21_addr),
    .io_mem_cluster_21_data(pipe10_io_mem_cluster_21_data),
    .io_mem_cluster_22_en(pipe10_io_mem_cluster_22_en),
    .io_mem_cluster_22_addr(pipe10_io_mem_cluster_22_addr),
    .io_mem_cluster_22_data(pipe10_io_mem_cluster_22_data),
    .io_mem_cluster_23_en(pipe10_io_mem_cluster_23_en),
    .io_mem_cluster_23_addr(pipe10_io_mem_cluster_23_addr),
    .io_mem_cluster_23_data(pipe10_io_mem_cluster_23_data),
    .io_mem_cluster_24_en(pipe10_io_mem_cluster_24_en),
    .io_mem_cluster_24_addr(pipe10_io_mem_cluster_24_addr),
    .io_mem_cluster_24_data(pipe10_io_mem_cluster_24_data),
    .io_mem_cluster_25_en(pipe10_io_mem_cluster_25_en),
    .io_mem_cluster_25_addr(pipe10_io_mem_cluster_25_addr),
    .io_mem_cluster_25_data(pipe10_io_mem_cluster_25_data),
    .io_mem_cluster_26_en(pipe10_io_mem_cluster_26_en),
    .io_mem_cluster_26_addr(pipe10_io_mem_cluster_26_addr),
    .io_mem_cluster_26_data(pipe10_io_mem_cluster_26_data),
    .io_mem_cluster_27_en(pipe10_io_mem_cluster_27_en),
    .io_mem_cluster_27_addr(pipe10_io_mem_cluster_27_addr),
    .io_mem_cluster_27_data(pipe10_io_mem_cluster_27_data),
    .io_mem_cluster_28_en(pipe10_io_mem_cluster_28_en),
    .io_mem_cluster_28_addr(pipe10_io_mem_cluster_28_addr),
    .io_mem_cluster_28_data(pipe10_io_mem_cluster_28_data),
    .io_mem_cluster_29_en(pipe10_io_mem_cluster_29_en),
    .io_mem_cluster_29_addr(pipe10_io_mem_cluster_29_addr),
    .io_mem_cluster_29_data(pipe10_io_mem_cluster_29_data),
    .io_mem_cluster_30_en(pipe10_io_mem_cluster_30_en),
    .io_mem_cluster_30_addr(pipe10_io_mem_cluster_30_addr),
    .io_mem_cluster_30_data(pipe10_io_mem_cluster_30_data),
    .io_mem_cluster_31_en(pipe10_io_mem_cluster_31_en),
    .io_mem_cluster_31_addr(pipe10_io_mem_cluster_31_addr),
    .io_mem_cluster_31_data(pipe10_io_mem_cluster_31_data),
    .io_mem_cluster_32_en(pipe10_io_mem_cluster_32_en),
    .io_mem_cluster_32_addr(pipe10_io_mem_cluster_32_addr),
    .io_mem_cluster_32_data(pipe10_io_mem_cluster_32_data),
    .io_mem_cluster_33_en(pipe10_io_mem_cluster_33_en),
    .io_mem_cluster_33_addr(pipe10_io_mem_cluster_33_addr),
    .io_mem_cluster_33_data(pipe10_io_mem_cluster_33_data),
    .io_mem_cluster_34_en(pipe10_io_mem_cluster_34_en),
    .io_mem_cluster_34_addr(pipe10_io_mem_cluster_34_addr),
    .io_mem_cluster_34_data(pipe10_io_mem_cluster_34_data),
    .io_mem_cluster_35_en(pipe10_io_mem_cluster_35_en),
    .io_mem_cluster_35_addr(pipe10_io_mem_cluster_35_addr),
    .io_mem_cluster_35_data(pipe10_io_mem_cluster_35_data),
    .io_mem_cluster_36_en(pipe10_io_mem_cluster_36_en),
    .io_mem_cluster_36_addr(pipe10_io_mem_cluster_36_addr),
    .io_mem_cluster_36_data(pipe10_io_mem_cluster_36_data),
    .io_mem_cluster_37_en(pipe10_io_mem_cluster_37_en),
    .io_mem_cluster_37_addr(pipe10_io_mem_cluster_37_addr),
    .io_mem_cluster_37_data(pipe10_io_mem_cluster_37_data),
    .io_mem_cluster_38_en(pipe10_io_mem_cluster_38_en),
    .io_mem_cluster_38_addr(pipe10_io_mem_cluster_38_addr),
    .io_mem_cluster_38_data(pipe10_io_mem_cluster_38_data),
    .io_mem_cluster_39_en(pipe10_io_mem_cluster_39_en),
    .io_mem_cluster_39_addr(pipe10_io_mem_cluster_39_addr),
    .io_mem_cluster_39_data(pipe10_io_mem_cluster_39_data),
    .io_mem_cluster_40_en(pipe10_io_mem_cluster_40_en),
    .io_mem_cluster_40_addr(pipe10_io_mem_cluster_40_addr),
    .io_mem_cluster_40_data(pipe10_io_mem_cluster_40_data),
    .io_mem_cluster_41_en(pipe10_io_mem_cluster_41_en),
    .io_mem_cluster_41_addr(pipe10_io_mem_cluster_41_addr),
    .io_mem_cluster_41_data(pipe10_io_mem_cluster_41_data),
    .io_mem_cluster_42_en(pipe10_io_mem_cluster_42_en),
    .io_mem_cluster_42_addr(pipe10_io_mem_cluster_42_addr),
    .io_mem_cluster_42_data(pipe10_io_mem_cluster_42_data),
    .io_mem_cluster_43_en(pipe10_io_mem_cluster_43_en),
    .io_mem_cluster_43_addr(pipe10_io_mem_cluster_43_addr),
    .io_mem_cluster_43_data(pipe10_io_mem_cluster_43_data),
    .io_mem_cluster_44_en(pipe10_io_mem_cluster_44_en),
    .io_mem_cluster_44_addr(pipe10_io_mem_cluster_44_addr),
    .io_mem_cluster_44_data(pipe10_io_mem_cluster_44_data),
    .io_mem_cluster_45_en(pipe10_io_mem_cluster_45_en),
    .io_mem_cluster_45_addr(pipe10_io_mem_cluster_45_addr),
    .io_mem_cluster_45_data(pipe10_io_mem_cluster_45_data),
    .io_mem_cluster_46_en(pipe10_io_mem_cluster_46_en),
    .io_mem_cluster_46_addr(pipe10_io_mem_cluster_46_addr),
    .io_mem_cluster_46_data(pipe10_io_mem_cluster_46_data),
    .io_mem_cluster_47_en(pipe10_io_mem_cluster_47_en),
    .io_mem_cluster_47_addr(pipe10_io_mem_cluster_47_addr),
    .io_mem_cluster_47_data(pipe10_io_mem_cluster_47_data),
    .io_mem_cluster_48_en(pipe10_io_mem_cluster_48_en),
    .io_mem_cluster_48_addr(pipe10_io_mem_cluster_48_addr),
    .io_mem_cluster_48_data(pipe10_io_mem_cluster_48_data),
    .io_mem_cluster_49_en(pipe10_io_mem_cluster_49_en),
    .io_mem_cluster_49_addr(pipe10_io_mem_cluster_49_addr),
    .io_mem_cluster_49_data(pipe10_io_mem_cluster_49_data),
    .io_mem_cluster_50_en(pipe10_io_mem_cluster_50_en),
    .io_mem_cluster_50_addr(pipe10_io_mem_cluster_50_addr),
    .io_mem_cluster_50_data(pipe10_io_mem_cluster_50_data),
    .io_mem_cluster_51_en(pipe10_io_mem_cluster_51_en),
    .io_mem_cluster_51_addr(pipe10_io_mem_cluster_51_addr),
    .io_mem_cluster_51_data(pipe10_io_mem_cluster_51_data),
    .io_mem_cluster_52_en(pipe10_io_mem_cluster_52_en),
    .io_mem_cluster_52_addr(pipe10_io_mem_cluster_52_addr),
    .io_mem_cluster_52_data(pipe10_io_mem_cluster_52_data),
    .io_mem_cluster_53_en(pipe10_io_mem_cluster_53_en),
    .io_mem_cluster_53_addr(pipe10_io_mem_cluster_53_addr),
    .io_mem_cluster_53_data(pipe10_io_mem_cluster_53_data),
    .io_mem_cluster_54_en(pipe10_io_mem_cluster_54_en),
    .io_mem_cluster_54_addr(pipe10_io_mem_cluster_54_addr),
    .io_mem_cluster_54_data(pipe10_io_mem_cluster_54_data),
    .io_mem_cluster_55_en(pipe10_io_mem_cluster_55_en),
    .io_mem_cluster_55_addr(pipe10_io_mem_cluster_55_addr),
    .io_mem_cluster_55_data(pipe10_io_mem_cluster_55_data),
    .io_mem_cluster_56_en(pipe10_io_mem_cluster_56_en),
    .io_mem_cluster_56_addr(pipe10_io_mem_cluster_56_addr),
    .io_mem_cluster_56_data(pipe10_io_mem_cluster_56_data),
    .io_mem_cluster_57_en(pipe10_io_mem_cluster_57_en),
    .io_mem_cluster_57_addr(pipe10_io_mem_cluster_57_addr),
    .io_mem_cluster_57_data(pipe10_io_mem_cluster_57_data),
    .io_mem_cluster_58_en(pipe10_io_mem_cluster_58_en),
    .io_mem_cluster_58_addr(pipe10_io_mem_cluster_58_addr),
    .io_mem_cluster_58_data(pipe10_io_mem_cluster_58_data),
    .io_mem_cluster_59_en(pipe10_io_mem_cluster_59_en),
    .io_mem_cluster_59_addr(pipe10_io_mem_cluster_59_addr),
    .io_mem_cluster_59_data(pipe10_io_mem_cluster_59_data),
    .io_mem_cluster_60_en(pipe10_io_mem_cluster_60_en),
    .io_mem_cluster_60_addr(pipe10_io_mem_cluster_60_addr),
    .io_mem_cluster_60_data(pipe10_io_mem_cluster_60_data),
    .io_mem_cluster_61_en(pipe10_io_mem_cluster_61_en),
    .io_mem_cluster_61_addr(pipe10_io_mem_cluster_61_addr),
    .io_mem_cluster_61_data(pipe10_io_mem_cluster_61_data),
    .io_mem_cluster_62_en(pipe10_io_mem_cluster_62_en),
    .io_mem_cluster_62_addr(pipe10_io_mem_cluster_62_addr),
    .io_mem_cluster_62_data(pipe10_io_mem_cluster_62_data),
    .io_mem_cluster_63_en(pipe10_io_mem_cluster_63_en),
    .io_mem_cluster_63_addr(pipe10_io_mem_cluster_63_addr),
    .io_mem_cluster_63_data(pipe10_io_mem_cluster_63_data)
  );
  MatchDataReshape pipe11 ( // @[matcher.scala 348:24]
    .clock(pipe11_clock),
    .io_pipe_phv_in_data_0(pipe11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe11_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe11_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe11_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe11_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe11_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe11_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe11_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe11_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe11_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe11_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe11_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe11_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe11_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe11_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe11_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe11_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe11_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe11_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe11_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe11_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe11_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe11_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe11_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe11_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe11_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe11_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe11_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe11_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe11_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe11_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe11_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe11_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe11_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe11_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe11_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe11_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe11_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe11_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe11_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe11_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe11_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe11_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe11_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe11_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe11_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe11_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe11_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe11_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe11_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe11_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe11_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe11_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe11_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe11_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe11_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe11_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe11_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe11_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe11_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe11_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe11_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe11_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe11_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe11_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe11_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe11_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe11_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe11_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe11_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe11_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe11_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe11_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe11_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe11_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe11_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe11_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe11_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe11_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe11_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe11_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe11_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe11_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe11_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe11_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe11_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe11_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe11_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe11_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe11_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe11_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe11_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe11_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe11_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe11_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe11_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe11_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe11_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe11_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe11_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe11_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe11_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe11_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe11_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe11_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe11_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe11_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe11_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe11_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe11_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe11_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe11_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe11_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe11_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe11_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe11_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe11_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe11_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe11_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe11_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe11_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe11_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe11_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe11_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe11_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe11_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe11_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe11_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe11_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe11_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe11_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe11_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe11_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe11_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe11_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe11_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe11_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe11_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe11_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe11_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe11_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe11_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe11_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe11_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe11_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe11_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe11_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe11_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe11_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe11_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe11_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe11_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe11_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe11_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe11_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe11_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe11_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe11_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe11_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe11_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe11_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe11_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe11_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe11_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe11_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe11_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe11_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe11_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe11_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe11_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe11_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe11_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe11_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe11_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe11_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe11_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe11_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe11_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe11_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe11_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe11_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe11_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe11_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe11_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe11_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe11_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe11_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe11_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe11_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe11_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe11_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe11_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe11_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe11_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe11_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe11_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe11_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe11_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe11_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe11_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe11_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe11_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe11_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe11_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe11_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe11_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe11_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe11_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe11_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe11_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe11_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe11_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe11_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe11_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe11_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe11_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe11_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe11_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe11_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe11_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe11_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe11_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe11_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe11_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe11_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe11_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe11_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe11_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe11_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe11_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe11_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe11_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe11_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe11_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe11_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe11_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe11_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe11_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe11_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe11_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe11_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe11_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe11_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe11_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe11_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe11_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe11_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe11_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe11_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe11_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe11_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe11_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe11_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe11_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe11_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe11_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe11_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe11_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe11_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe11_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe11_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe11_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe11_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe11_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe11_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe11_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe11_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe11_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe11_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe11_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe11_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe11_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe11_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe11_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe11_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe11_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe11_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe11_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe11_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe11_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe11_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe11_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe11_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe11_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe11_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe11_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe11_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe11_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe11_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe11_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe11_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe11_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe11_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe11_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe11_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe11_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe11_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe11_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe11_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe11_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe11_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe11_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe11_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe11_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe11_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe11_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe11_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe11_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe11_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe11_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe11_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe11_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe11_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe11_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe11_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe11_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe11_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe11_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe11_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe11_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe11_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe11_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe11_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe11_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe11_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe11_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe11_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe11_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe11_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe11_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe11_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe11_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe11_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe11_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe11_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe11_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe11_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe11_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe11_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe11_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe11_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe11_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe11_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe11_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe11_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe11_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe11_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe11_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe11_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe11_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe11_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe11_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe11_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe11_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe11_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe11_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe11_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe11_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe11_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe11_io_pipe_phv_out_is_valid_processor),
    .io_table_config_0_table_width(pipe11_io_table_config_0_table_width),
    .io_table_config_0_table_depth(pipe11_io_table_config_0_table_depth),
    .io_table_config_1_table_width(pipe11_io_table_config_1_table_width),
    .io_table_config_1_table_depth(pipe11_io_table_config_1_table_depth),
    .io_key_in(pipe11_io_key_in),
    .io_key_out(pipe11_io_key_out),
    .io_cs_in(pipe11_io_cs_in),
    .io_data_in_0(pipe11_io_data_in_0),
    .io_data_in_1(pipe11_io_data_in_1),
    .io_data_in_2(pipe11_io_data_in_2),
    .io_data_in_3(pipe11_io_data_in_3),
    .io_data_in_4(pipe11_io_data_in_4),
    .io_data_in_5(pipe11_io_data_in_5),
    .io_data_in_6(pipe11_io_data_in_6),
    .io_data_in_7(pipe11_io_data_in_7),
    .io_data_in_8(pipe11_io_data_in_8),
    .io_data_in_9(pipe11_io_data_in_9),
    .io_data_in_10(pipe11_io_data_in_10),
    .io_data_in_11(pipe11_io_data_in_11),
    .io_data_in_12(pipe11_io_data_in_12),
    .io_data_in_13(pipe11_io_data_in_13),
    .io_data_in_14(pipe11_io_data_in_14),
    .io_data_in_15(pipe11_io_data_in_15),
    .io_data_in_16(pipe11_io_data_in_16),
    .io_data_in_17(pipe11_io_data_in_17),
    .io_data_in_18(pipe11_io_data_in_18),
    .io_data_in_19(pipe11_io_data_in_19),
    .io_data_in_20(pipe11_io_data_in_20),
    .io_data_in_21(pipe11_io_data_in_21),
    .io_data_in_22(pipe11_io_data_in_22),
    .io_data_in_23(pipe11_io_data_in_23),
    .io_data_in_24(pipe11_io_data_in_24),
    .io_data_in_25(pipe11_io_data_in_25),
    .io_data_in_26(pipe11_io_data_in_26),
    .io_data_in_27(pipe11_io_data_in_27),
    .io_data_in_28(pipe11_io_data_in_28),
    .io_data_in_29(pipe11_io_data_in_29),
    .io_data_in_30(pipe11_io_data_in_30),
    .io_data_in_31(pipe11_io_data_in_31),
    .io_data_in_32(pipe11_io_data_in_32),
    .io_data_in_33(pipe11_io_data_in_33),
    .io_data_in_34(pipe11_io_data_in_34),
    .io_data_in_35(pipe11_io_data_in_35),
    .io_data_in_36(pipe11_io_data_in_36),
    .io_data_in_37(pipe11_io_data_in_37),
    .io_data_in_38(pipe11_io_data_in_38),
    .io_data_in_39(pipe11_io_data_in_39),
    .io_data_in_40(pipe11_io_data_in_40),
    .io_data_in_41(pipe11_io_data_in_41),
    .io_data_in_42(pipe11_io_data_in_42),
    .io_data_in_43(pipe11_io_data_in_43),
    .io_data_in_44(pipe11_io_data_in_44),
    .io_data_in_45(pipe11_io_data_in_45),
    .io_data_in_46(pipe11_io_data_in_46),
    .io_data_in_47(pipe11_io_data_in_47),
    .io_data_in_48(pipe11_io_data_in_48),
    .io_data_in_49(pipe11_io_data_in_49),
    .io_data_in_50(pipe11_io_data_in_50),
    .io_data_in_51(pipe11_io_data_in_51),
    .io_data_in_52(pipe11_io_data_in_52),
    .io_data_in_53(pipe11_io_data_in_53),
    .io_data_in_54(pipe11_io_data_in_54),
    .io_data_in_55(pipe11_io_data_in_55),
    .io_data_in_56(pipe11_io_data_in_56),
    .io_data_in_57(pipe11_io_data_in_57),
    .io_data_in_58(pipe11_io_data_in_58),
    .io_data_in_59(pipe11_io_data_in_59),
    .io_data_in_60(pipe11_io_data_in_60),
    .io_data_in_61(pipe11_io_data_in_61),
    .io_data_in_62(pipe11_io_data_in_62),
    .io_data_in_63(pipe11_io_data_in_63),
    .io_data_out(pipe11_io_data_out)
  );
  MatchResult pipe12 ( // @[matcher.scala 349:24]
    .clock(pipe12_clock),
    .io_pipe_phv_in_data_0(pipe12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe12_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe12_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe12_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe12_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe12_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe12_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe12_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe12_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe12_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe12_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe12_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe12_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe12_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe12_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe12_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe12_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe12_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe12_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe12_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe12_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe12_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe12_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe12_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe12_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe12_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe12_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe12_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe12_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe12_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe12_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe12_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe12_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe12_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe12_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe12_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe12_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe12_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe12_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe12_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe12_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe12_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe12_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe12_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe12_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe12_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe12_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe12_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe12_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe12_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe12_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe12_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe12_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe12_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe12_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe12_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe12_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe12_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe12_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe12_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe12_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe12_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe12_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe12_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe12_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe12_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe12_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe12_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe12_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe12_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe12_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe12_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe12_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe12_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe12_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe12_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe12_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe12_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe12_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe12_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe12_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe12_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe12_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe12_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe12_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe12_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe12_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe12_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe12_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe12_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe12_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe12_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe12_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe12_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe12_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe12_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe12_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe12_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe12_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe12_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe12_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe12_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe12_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe12_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe12_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe12_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe12_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe12_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe12_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe12_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe12_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe12_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe12_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe12_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe12_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe12_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe12_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe12_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe12_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe12_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe12_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe12_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe12_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe12_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe12_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe12_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe12_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe12_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe12_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe12_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe12_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe12_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe12_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe12_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe12_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe12_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe12_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe12_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe12_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe12_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe12_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe12_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe12_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe12_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe12_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe12_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe12_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe12_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe12_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe12_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe12_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe12_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe12_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe12_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe12_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe12_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe12_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe12_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe12_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe12_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe12_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe12_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe12_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe12_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe12_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe12_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe12_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe12_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe12_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe12_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe12_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe12_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe12_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe12_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe12_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe12_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe12_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe12_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe12_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe12_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe12_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe12_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe12_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe12_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe12_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe12_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe12_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe12_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe12_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe12_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe12_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe12_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe12_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe12_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe12_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe12_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe12_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe12_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe12_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe12_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe12_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe12_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe12_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe12_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe12_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe12_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe12_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe12_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe12_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe12_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe12_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe12_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe12_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe12_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe12_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe12_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe12_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe12_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe12_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe12_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe12_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe12_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe12_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe12_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe12_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe12_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe12_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe12_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe12_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe12_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe12_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe12_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe12_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe12_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe12_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe12_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe12_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe12_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe12_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe12_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe12_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe12_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe12_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe12_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe12_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe12_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe12_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe12_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe12_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe12_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe12_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe12_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe12_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe12_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe12_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe12_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe12_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe12_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe12_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe12_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe12_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe12_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe12_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe12_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe12_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe12_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe12_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe12_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe12_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe12_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe12_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe12_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe12_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe12_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe12_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe12_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe12_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe12_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe12_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe12_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe12_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe12_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe12_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe12_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe12_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe12_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe12_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe12_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe12_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe12_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe12_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe12_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe12_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe12_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe12_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe12_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe12_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe12_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe12_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe12_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe12_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe12_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe12_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe12_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe12_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe12_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe12_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe12_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe12_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe12_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe12_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe12_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe12_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe12_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe12_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe12_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe12_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe12_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe12_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe12_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe12_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe12_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe12_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe12_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe12_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe12_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe12_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe12_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe12_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe12_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe12_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe12_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe12_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe12_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe12_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe12_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe12_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe12_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe12_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe12_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe12_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe12_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe12_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe12_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe12_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe12_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe12_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe12_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe12_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe12_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe12_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe12_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe12_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe12_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe12_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe12_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe12_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe12_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe12_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe12_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe12_io_pipe_phv_out_is_valid_processor),
    .io_key_config_0_key_length(pipe12_io_key_config_0_key_length),
    .io_key_config_1_key_length(pipe12_io_key_config_1_key_length),
    .io_key_in(pipe12_io_key_in),
    .io_data_in(pipe12_io_data_in),
    .io_hit(pipe12_io_hit),
    .io_match_value(pipe12_io_match_value)
  );
  assign io_pipe_phv_out_data_0 = pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_1 = pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_2 = pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_3 = pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_4 = pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_5 = pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_6 = pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_7 = pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_8 = pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_9 = pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_10 = pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_11 = pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_12 = pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_13 = pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_14 = pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_15 = pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_16 = pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_17 = pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_18 = pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_19 = pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_20 = pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_21 = pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_22 = pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_23 = pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_24 = pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_25 = pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_26 = pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_27 = pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_28 = pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_29 = pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_30 = pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_31 = pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_32 = pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_33 = pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_34 = pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_35 = pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_36 = pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_37 = pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_38 = pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_39 = pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_40 = pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_41 = pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_42 = pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_43 = pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_44 = pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_45 = pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_46 = pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_47 = pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_48 = pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_49 = pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_50 = pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_51 = pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_52 = pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_53 = pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_54 = pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_55 = pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_56 = pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_57 = pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_58 = pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_59 = pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_60 = pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_61 = pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_62 = pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_63 = pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_64 = pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_65 = pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_66 = pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_67 = pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_68 = pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_69 = pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_70 = pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_71 = pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_72 = pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_73 = pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_74 = pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_75 = pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_76 = pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_77 = pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_78 = pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_79 = pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_80 = pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_81 = pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_82 = pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_83 = pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_84 = pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_85 = pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_86 = pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_87 = pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_88 = pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_89 = pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_90 = pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_91 = pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_92 = pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_93 = pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_94 = pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_95 = pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_96 = pipe12_io_pipe_phv_out_data_96; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_97 = pipe12_io_pipe_phv_out_data_97; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_98 = pipe12_io_pipe_phv_out_data_98; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_99 = pipe12_io_pipe_phv_out_data_99; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_100 = pipe12_io_pipe_phv_out_data_100; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_101 = pipe12_io_pipe_phv_out_data_101; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_102 = pipe12_io_pipe_phv_out_data_102; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_103 = pipe12_io_pipe_phv_out_data_103; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_104 = pipe12_io_pipe_phv_out_data_104; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_105 = pipe12_io_pipe_phv_out_data_105; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_106 = pipe12_io_pipe_phv_out_data_106; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_107 = pipe12_io_pipe_phv_out_data_107; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_108 = pipe12_io_pipe_phv_out_data_108; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_109 = pipe12_io_pipe_phv_out_data_109; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_110 = pipe12_io_pipe_phv_out_data_110; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_111 = pipe12_io_pipe_phv_out_data_111; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_112 = pipe12_io_pipe_phv_out_data_112; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_113 = pipe12_io_pipe_phv_out_data_113; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_114 = pipe12_io_pipe_phv_out_data_114; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_115 = pipe12_io_pipe_phv_out_data_115; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_116 = pipe12_io_pipe_phv_out_data_116; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_117 = pipe12_io_pipe_phv_out_data_117; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_118 = pipe12_io_pipe_phv_out_data_118; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_119 = pipe12_io_pipe_phv_out_data_119; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_120 = pipe12_io_pipe_phv_out_data_120; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_121 = pipe12_io_pipe_phv_out_data_121; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_122 = pipe12_io_pipe_phv_out_data_122; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_123 = pipe12_io_pipe_phv_out_data_123; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_124 = pipe12_io_pipe_phv_out_data_124; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_125 = pipe12_io_pipe_phv_out_data_125; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_126 = pipe12_io_pipe_phv_out_data_126; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_127 = pipe12_io_pipe_phv_out_data_127; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_128 = pipe12_io_pipe_phv_out_data_128; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_129 = pipe12_io_pipe_phv_out_data_129; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_130 = pipe12_io_pipe_phv_out_data_130; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_131 = pipe12_io_pipe_phv_out_data_131; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_132 = pipe12_io_pipe_phv_out_data_132; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_133 = pipe12_io_pipe_phv_out_data_133; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_134 = pipe12_io_pipe_phv_out_data_134; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_135 = pipe12_io_pipe_phv_out_data_135; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_136 = pipe12_io_pipe_phv_out_data_136; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_137 = pipe12_io_pipe_phv_out_data_137; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_138 = pipe12_io_pipe_phv_out_data_138; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_139 = pipe12_io_pipe_phv_out_data_139; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_140 = pipe12_io_pipe_phv_out_data_140; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_141 = pipe12_io_pipe_phv_out_data_141; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_142 = pipe12_io_pipe_phv_out_data_142; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_143 = pipe12_io_pipe_phv_out_data_143; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_144 = pipe12_io_pipe_phv_out_data_144; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_145 = pipe12_io_pipe_phv_out_data_145; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_146 = pipe12_io_pipe_phv_out_data_146; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_147 = pipe12_io_pipe_phv_out_data_147; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_148 = pipe12_io_pipe_phv_out_data_148; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_149 = pipe12_io_pipe_phv_out_data_149; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_150 = pipe12_io_pipe_phv_out_data_150; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_151 = pipe12_io_pipe_phv_out_data_151; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_152 = pipe12_io_pipe_phv_out_data_152; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_153 = pipe12_io_pipe_phv_out_data_153; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_154 = pipe12_io_pipe_phv_out_data_154; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_155 = pipe12_io_pipe_phv_out_data_155; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_156 = pipe12_io_pipe_phv_out_data_156; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_157 = pipe12_io_pipe_phv_out_data_157; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_158 = pipe12_io_pipe_phv_out_data_158; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_159 = pipe12_io_pipe_phv_out_data_159; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_160 = pipe12_io_pipe_phv_out_data_160; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_161 = pipe12_io_pipe_phv_out_data_161; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_162 = pipe12_io_pipe_phv_out_data_162; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_163 = pipe12_io_pipe_phv_out_data_163; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_164 = pipe12_io_pipe_phv_out_data_164; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_165 = pipe12_io_pipe_phv_out_data_165; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_166 = pipe12_io_pipe_phv_out_data_166; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_167 = pipe12_io_pipe_phv_out_data_167; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_168 = pipe12_io_pipe_phv_out_data_168; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_169 = pipe12_io_pipe_phv_out_data_169; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_170 = pipe12_io_pipe_phv_out_data_170; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_171 = pipe12_io_pipe_phv_out_data_171; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_172 = pipe12_io_pipe_phv_out_data_172; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_173 = pipe12_io_pipe_phv_out_data_173; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_174 = pipe12_io_pipe_phv_out_data_174; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_175 = pipe12_io_pipe_phv_out_data_175; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_176 = pipe12_io_pipe_phv_out_data_176; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_177 = pipe12_io_pipe_phv_out_data_177; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_178 = pipe12_io_pipe_phv_out_data_178; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_179 = pipe12_io_pipe_phv_out_data_179; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_180 = pipe12_io_pipe_phv_out_data_180; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_181 = pipe12_io_pipe_phv_out_data_181; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_182 = pipe12_io_pipe_phv_out_data_182; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_183 = pipe12_io_pipe_phv_out_data_183; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_184 = pipe12_io_pipe_phv_out_data_184; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_185 = pipe12_io_pipe_phv_out_data_185; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_186 = pipe12_io_pipe_phv_out_data_186; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_187 = pipe12_io_pipe_phv_out_data_187; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_188 = pipe12_io_pipe_phv_out_data_188; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_189 = pipe12_io_pipe_phv_out_data_189; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_190 = pipe12_io_pipe_phv_out_data_190; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_191 = pipe12_io_pipe_phv_out_data_191; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_192 = pipe12_io_pipe_phv_out_data_192; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_193 = pipe12_io_pipe_phv_out_data_193; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_194 = pipe12_io_pipe_phv_out_data_194; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_195 = pipe12_io_pipe_phv_out_data_195; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_196 = pipe12_io_pipe_phv_out_data_196; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_197 = pipe12_io_pipe_phv_out_data_197; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_198 = pipe12_io_pipe_phv_out_data_198; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_199 = pipe12_io_pipe_phv_out_data_199; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_200 = pipe12_io_pipe_phv_out_data_200; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_201 = pipe12_io_pipe_phv_out_data_201; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_202 = pipe12_io_pipe_phv_out_data_202; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_203 = pipe12_io_pipe_phv_out_data_203; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_204 = pipe12_io_pipe_phv_out_data_204; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_205 = pipe12_io_pipe_phv_out_data_205; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_206 = pipe12_io_pipe_phv_out_data_206; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_207 = pipe12_io_pipe_phv_out_data_207; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_208 = pipe12_io_pipe_phv_out_data_208; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_209 = pipe12_io_pipe_phv_out_data_209; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_210 = pipe12_io_pipe_phv_out_data_210; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_211 = pipe12_io_pipe_phv_out_data_211; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_212 = pipe12_io_pipe_phv_out_data_212; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_213 = pipe12_io_pipe_phv_out_data_213; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_214 = pipe12_io_pipe_phv_out_data_214; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_215 = pipe12_io_pipe_phv_out_data_215; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_216 = pipe12_io_pipe_phv_out_data_216; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_217 = pipe12_io_pipe_phv_out_data_217; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_218 = pipe12_io_pipe_phv_out_data_218; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_219 = pipe12_io_pipe_phv_out_data_219; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_220 = pipe12_io_pipe_phv_out_data_220; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_221 = pipe12_io_pipe_phv_out_data_221; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_222 = pipe12_io_pipe_phv_out_data_222; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_223 = pipe12_io_pipe_phv_out_data_223; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_224 = pipe12_io_pipe_phv_out_data_224; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_225 = pipe12_io_pipe_phv_out_data_225; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_226 = pipe12_io_pipe_phv_out_data_226; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_227 = pipe12_io_pipe_phv_out_data_227; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_228 = pipe12_io_pipe_phv_out_data_228; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_229 = pipe12_io_pipe_phv_out_data_229; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_230 = pipe12_io_pipe_phv_out_data_230; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_231 = pipe12_io_pipe_phv_out_data_231; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_232 = pipe12_io_pipe_phv_out_data_232; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_233 = pipe12_io_pipe_phv_out_data_233; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_234 = pipe12_io_pipe_phv_out_data_234; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_235 = pipe12_io_pipe_phv_out_data_235; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_236 = pipe12_io_pipe_phv_out_data_236; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_237 = pipe12_io_pipe_phv_out_data_237; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_238 = pipe12_io_pipe_phv_out_data_238; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_239 = pipe12_io_pipe_phv_out_data_239; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_240 = pipe12_io_pipe_phv_out_data_240; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_241 = pipe12_io_pipe_phv_out_data_241; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_242 = pipe12_io_pipe_phv_out_data_242; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_243 = pipe12_io_pipe_phv_out_data_243; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_244 = pipe12_io_pipe_phv_out_data_244; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_245 = pipe12_io_pipe_phv_out_data_245; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_246 = pipe12_io_pipe_phv_out_data_246; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_247 = pipe12_io_pipe_phv_out_data_247; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_248 = pipe12_io_pipe_phv_out_data_248; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_249 = pipe12_io_pipe_phv_out_data_249; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_250 = pipe12_io_pipe_phv_out_data_250; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_251 = pipe12_io_pipe_phv_out_data_251; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_252 = pipe12_io_pipe_phv_out_data_252; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_253 = pipe12_io_pipe_phv_out_data_253; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_254 = pipe12_io_pipe_phv_out_data_254; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_255 = pipe12_io_pipe_phv_out_data_255; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_0 = pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_1 = pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_2 = pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_3 = pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_4 = pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_5 = pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_6 = pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_7 = pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_8 = pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_9 = pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_10 = pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_11 = pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_12 = pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_13 = pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_14 = pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_15 = pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_current_state = pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_current_offset = pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_transition_field = pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_next_processor_id = pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_next_config_id = pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_is_valid_processor = pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 388:27]
  assign io_hit = pipe12_io_hit; // @[matcher.scala 389:27]
  assign io_match_value = pipe12_io_match_value; // @[matcher.scala 390:27]
  assign io_mem_cluster_0_en = pipe10_io_mem_cluster_0_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_0_addr = pipe10_io_mem_cluster_0_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_1_en = pipe10_io_mem_cluster_1_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_1_addr = pipe10_io_mem_cluster_1_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_2_en = pipe10_io_mem_cluster_2_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_2_addr = pipe10_io_mem_cluster_2_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_3_en = pipe10_io_mem_cluster_3_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_3_addr = pipe10_io_mem_cluster_3_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_4_en = pipe10_io_mem_cluster_4_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_4_addr = pipe10_io_mem_cluster_4_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_5_en = pipe10_io_mem_cluster_5_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_5_addr = pipe10_io_mem_cluster_5_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_6_en = pipe10_io_mem_cluster_6_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_6_addr = pipe10_io_mem_cluster_6_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_7_en = pipe10_io_mem_cluster_7_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_7_addr = pipe10_io_mem_cluster_7_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_8_en = pipe10_io_mem_cluster_8_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_8_addr = pipe10_io_mem_cluster_8_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_9_en = pipe10_io_mem_cluster_9_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_9_addr = pipe10_io_mem_cluster_9_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_10_en = pipe10_io_mem_cluster_10_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_10_addr = pipe10_io_mem_cluster_10_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_11_en = pipe10_io_mem_cluster_11_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_11_addr = pipe10_io_mem_cluster_11_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_12_en = pipe10_io_mem_cluster_12_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_12_addr = pipe10_io_mem_cluster_12_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_13_en = pipe10_io_mem_cluster_13_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_13_addr = pipe10_io_mem_cluster_13_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_14_en = pipe10_io_mem_cluster_14_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_14_addr = pipe10_io_mem_cluster_14_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_15_en = pipe10_io_mem_cluster_15_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_15_addr = pipe10_io_mem_cluster_15_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_16_en = pipe10_io_mem_cluster_16_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_16_addr = pipe10_io_mem_cluster_16_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_17_en = pipe10_io_mem_cluster_17_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_17_addr = pipe10_io_mem_cluster_17_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_18_en = pipe10_io_mem_cluster_18_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_18_addr = pipe10_io_mem_cluster_18_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_19_en = pipe10_io_mem_cluster_19_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_19_addr = pipe10_io_mem_cluster_19_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_20_en = pipe10_io_mem_cluster_20_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_20_addr = pipe10_io_mem_cluster_20_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_21_en = pipe10_io_mem_cluster_21_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_21_addr = pipe10_io_mem_cluster_21_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_22_en = pipe10_io_mem_cluster_22_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_22_addr = pipe10_io_mem_cluster_22_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_23_en = pipe10_io_mem_cluster_23_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_23_addr = pipe10_io_mem_cluster_23_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_24_en = pipe10_io_mem_cluster_24_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_24_addr = pipe10_io_mem_cluster_24_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_25_en = pipe10_io_mem_cluster_25_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_25_addr = pipe10_io_mem_cluster_25_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_26_en = pipe10_io_mem_cluster_26_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_26_addr = pipe10_io_mem_cluster_26_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_27_en = pipe10_io_mem_cluster_27_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_27_addr = pipe10_io_mem_cluster_27_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_28_en = pipe10_io_mem_cluster_28_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_28_addr = pipe10_io_mem_cluster_28_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_29_en = pipe10_io_mem_cluster_29_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_29_addr = pipe10_io_mem_cluster_29_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_30_en = pipe10_io_mem_cluster_30_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_30_addr = pipe10_io_mem_cluster_30_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_31_en = pipe10_io_mem_cluster_31_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_31_addr = pipe10_io_mem_cluster_31_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_32_en = pipe10_io_mem_cluster_32_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_32_addr = pipe10_io_mem_cluster_32_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_33_en = pipe10_io_mem_cluster_33_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_33_addr = pipe10_io_mem_cluster_33_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_34_en = pipe10_io_mem_cluster_34_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_34_addr = pipe10_io_mem_cluster_34_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_35_en = pipe10_io_mem_cluster_35_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_35_addr = pipe10_io_mem_cluster_35_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_36_en = pipe10_io_mem_cluster_36_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_36_addr = pipe10_io_mem_cluster_36_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_37_en = pipe10_io_mem_cluster_37_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_37_addr = pipe10_io_mem_cluster_37_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_38_en = pipe10_io_mem_cluster_38_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_38_addr = pipe10_io_mem_cluster_38_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_39_en = pipe10_io_mem_cluster_39_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_39_addr = pipe10_io_mem_cluster_39_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_40_en = pipe10_io_mem_cluster_40_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_40_addr = pipe10_io_mem_cluster_40_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_41_en = pipe10_io_mem_cluster_41_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_41_addr = pipe10_io_mem_cluster_41_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_42_en = pipe10_io_mem_cluster_42_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_42_addr = pipe10_io_mem_cluster_42_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_43_en = pipe10_io_mem_cluster_43_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_43_addr = pipe10_io_mem_cluster_43_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_44_en = pipe10_io_mem_cluster_44_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_44_addr = pipe10_io_mem_cluster_44_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_45_en = pipe10_io_mem_cluster_45_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_45_addr = pipe10_io_mem_cluster_45_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_46_en = pipe10_io_mem_cluster_46_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_46_addr = pipe10_io_mem_cluster_46_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_47_en = pipe10_io_mem_cluster_47_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_47_addr = pipe10_io_mem_cluster_47_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_48_en = pipe10_io_mem_cluster_48_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_48_addr = pipe10_io_mem_cluster_48_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_49_en = pipe10_io_mem_cluster_49_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_49_addr = pipe10_io_mem_cluster_49_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_50_en = pipe10_io_mem_cluster_50_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_50_addr = pipe10_io_mem_cluster_50_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_51_en = pipe10_io_mem_cluster_51_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_51_addr = pipe10_io_mem_cluster_51_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_52_en = pipe10_io_mem_cluster_52_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_52_addr = pipe10_io_mem_cluster_52_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_53_en = pipe10_io_mem_cluster_53_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_53_addr = pipe10_io_mem_cluster_53_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_54_en = pipe10_io_mem_cluster_54_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_54_addr = pipe10_io_mem_cluster_54_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_55_en = pipe10_io_mem_cluster_55_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_55_addr = pipe10_io_mem_cluster_55_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_56_en = pipe10_io_mem_cluster_56_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_56_addr = pipe10_io_mem_cluster_56_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_57_en = pipe10_io_mem_cluster_57_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_57_addr = pipe10_io_mem_cluster_57_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_58_en = pipe10_io_mem_cluster_58_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_58_addr = pipe10_io_mem_cluster_58_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_59_en = pipe10_io_mem_cluster_59_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_59_addr = pipe10_io_mem_cluster_59_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_60_en = pipe10_io_mem_cluster_60_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_60_addr = pipe10_io_mem_cluster_60_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_61_en = pipe10_io_mem_cluster_61_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_61_addr = pipe10_io_mem_cluster_61_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_62_en = pipe10_io_mem_cluster_62_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_62_addr = pipe10_io_mem_cluster_62_addr; // @[matcher.scala 375:27]
  assign io_mem_cluster_63_en = pipe10_io_mem_cluster_63_en; // @[matcher.scala 375:27]
  assign io_mem_cluster_63_addr = pipe10_io_mem_cluster_63_addr; // @[matcher.scala 375:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[matcher.scala 351:26]
  assign pipe1_io_key_config_0_header_id = key_config_0_header_id; // @[matcher.scala 352:26]
  assign pipe1_io_key_config_0_internal_offset = key_config_0_internal_offset; // @[matcher.scala 352:26]
  assign pipe1_io_key_config_1_header_id = key_config_1_header_id; // @[matcher.scala 352:26]
  assign pipe1_io_key_config_1_internal_offset = key_config_1_internal_offset; // @[matcher.scala 352:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 354:26]
  assign pipe2_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 356:26]
  assign pipe2_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 356:26]
  assign pipe2_io_key_offset = pipe1_io_key_offset; // @[matcher.scala 355:26]
  assign pipe3to8_clock = clock;
  assign pipe3to8_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 358:29]
  assign pipe3to8_io_mod_hash_depth_mod = io_mod_en; // @[matcher.scala 359:36]
  assign pipe3to8_io_mod_config_id = io_mod_config_id; // @[matcher.scala 360:36]
  assign pipe3to8_io_mod_hash_depth = io_mod_table_mod_table_depth[5:0]; // @[matcher.scala 361:36]
  assign pipe3to8_io_key_in = pipe2_io_match_key; // @[matcher.scala 362:26]
  assign pipe9_clock = clock;
  assign pipe9_io_pipe_phv_in_data_0 = pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_1 = pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_2 = pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_3 = pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_4 = pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_5 = pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_6 = pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_7 = pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_8 = pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_9 = pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_10 = pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_11 = pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_12 = pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_13 = pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_14 = pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_15 = pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_16 = pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_17 = pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_18 = pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_19 = pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_20 = pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_21 = pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_22 = pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_23 = pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_24 = pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_25 = pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_26 = pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_27 = pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_28 = pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_29 = pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_30 = pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_31 = pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_32 = pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_33 = pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_34 = pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_35 = pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_36 = pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_37 = pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_38 = pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_39 = pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_40 = pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_41 = pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_42 = pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_43 = pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_44 = pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_45 = pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_46 = pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_47 = pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_48 = pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_49 = pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_50 = pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_51 = pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_52 = pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_53 = pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_54 = pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_55 = pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_56 = pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_57 = pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_58 = pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_59 = pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_60 = pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_61 = pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_62 = pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_63 = pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_64 = pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_65 = pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_66 = pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_67 = pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_68 = pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_69 = pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_70 = pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_71 = pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_72 = pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_73 = pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_74 = pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_75 = pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_76 = pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_77 = pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_78 = pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_79 = pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_80 = pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_81 = pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_82 = pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_83 = pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_84 = pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_85 = pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_86 = pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_87 = pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_88 = pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_89 = pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_90 = pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_91 = pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_92 = pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_93 = pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_94 = pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_95 = pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_96 = pipe3to8_io_pipe_phv_out_data_96; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_97 = pipe3to8_io_pipe_phv_out_data_97; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_98 = pipe3to8_io_pipe_phv_out_data_98; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_99 = pipe3to8_io_pipe_phv_out_data_99; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_100 = pipe3to8_io_pipe_phv_out_data_100; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_101 = pipe3to8_io_pipe_phv_out_data_101; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_102 = pipe3to8_io_pipe_phv_out_data_102; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_103 = pipe3to8_io_pipe_phv_out_data_103; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_104 = pipe3to8_io_pipe_phv_out_data_104; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_105 = pipe3to8_io_pipe_phv_out_data_105; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_106 = pipe3to8_io_pipe_phv_out_data_106; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_107 = pipe3to8_io_pipe_phv_out_data_107; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_108 = pipe3to8_io_pipe_phv_out_data_108; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_109 = pipe3to8_io_pipe_phv_out_data_109; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_110 = pipe3to8_io_pipe_phv_out_data_110; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_111 = pipe3to8_io_pipe_phv_out_data_111; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_112 = pipe3to8_io_pipe_phv_out_data_112; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_113 = pipe3to8_io_pipe_phv_out_data_113; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_114 = pipe3to8_io_pipe_phv_out_data_114; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_115 = pipe3to8_io_pipe_phv_out_data_115; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_116 = pipe3to8_io_pipe_phv_out_data_116; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_117 = pipe3to8_io_pipe_phv_out_data_117; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_118 = pipe3to8_io_pipe_phv_out_data_118; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_119 = pipe3to8_io_pipe_phv_out_data_119; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_120 = pipe3to8_io_pipe_phv_out_data_120; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_121 = pipe3to8_io_pipe_phv_out_data_121; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_122 = pipe3to8_io_pipe_phv_out_data_122; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_123 = pipe3to8_io_pipe_phv_out_data_123; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_124 = pipe3to8_io_pipe_phv_out_data_124; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_125 = pipe3to8_io_pipe_phv_out_data_125; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_126 = pipe3to8_io_pipe_phv_out_data_126; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_127 = pipe3to8_io_pipe_phv_out_data_127; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_128 = pipe3to8_io_pipe_phv_out_data_128; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_129 = pipe3to8_io_pipe_phv_out_data_129; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_130 = pipe3to8_io_pipe_phv_out_data_130; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_131 = pipe3to8_io_pipe_phv_out_data_131; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_132 = pipe3to8_io_pipe_phv_out_data_132; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_133 = pipe3to8_io_pipe_phv_out_data_133; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_134 = pipe3to8_io_pipe_phv_out_data_134; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_135 = pipe3to8_io_pipe_phv_out_data_135; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_136 = pipe3to8_io_pipe_phv_out_data_136; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_137 = pipe3to8_io_pipe_phv_out_data_137; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_138 = pipe3to8_io_pipe_phv_out_data_138; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_139 = pipe3to8_io_pipe_phv_out_data_139; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_140 = pipe3to8_io_pipe_phv_out_data_140; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_141 = pipe3to8_io_pipe_phv_out_data_141; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_142 = pipe3to8_io_pipe_phv_out_data_142; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_143 = pipe3to8_io_pipe_phv_out_data_143; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_144 = pipe3to8_io_pipe_phv_out_data_144; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_145 = pipe3to8_io_pipe_phv_out_data_145; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_146 = pipe3to8_io_pipe_phv_out_data_146; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_147 = pipe3to8_io_pipe_phv_out_data_147; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_148 = pipe3to8_io_pipe_phv_out_data_148; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_149 = pipe3to8_io_pipe_phv_out_data_149; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_150 = pipe3to8_io_pipe_phv_out_data_150; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_151 = pipe3to8_io_pipe_phv_out_data_151; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_152 = pipe3to8_io_pipe_phv_out_data_152; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_153 = pipe3to8_io_pipe_phv_out_data_153; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_154 = pipe3to8_io_pipe_phv_out_data_154; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_155 = pipe3to8_io_pipe_phv_out_data_155; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_156 = pipe3to8_io_pipe_phv_out_data_156; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_157 = pipe3to8_io_pipe_phv_out_data_157; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_158 = pipe3to8_io_pipe_phv_out_data_158; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_159 = pipe3to8_io_pipe_phv_out_data_159; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_160 = pipe3to8_io_pipe_phv_out_data_160; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_161 = pipe3to8_io_pipe_phv_out_data_161; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_162 = pipe3to8_io_pipe_phv_out_data_162; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_163 = pipe3to8_io_pipe_phv_out_data_163; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_164 = pipe3to8_io_pipe_phv_out_data_164; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_165 = pipe3to8_io_pipe_phv_out_data_165; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_166 = pipe3to8_io_pipe_phv_out_data_166; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_167 = pipe3to8_io_pipe_phv_out_data_167; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_168 = pipe3to8_io_pipe_phv_out_data_168; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_169 = pipe3to8_io_pipe_phv_out_data_169; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_170 = pipe3to8_io_pipe_phv_out_data_170; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_171 = pipe3to8_io_pipe_phv_out_data_171; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_172 = pipe3to8_io_pipe_phv_out_data_172; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_173 = pipe3to8_io_pipe_phv_out_data_173; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_174 = pipe3to8_io_pipe_phv_out_data_174; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_175 = pipe3to8_io_pipe_phv_out_data_175; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_176 = pipe3to8_io_pipe_phv_out_data_176; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_177 = pipe3to8_io_pipe_phv_out_data_177; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_178 = pipe3to8_io_pipe_phv_out_data_178; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_179 = pipe3to8_io_pipe_phv_out_data_179; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_180 = pipe3to8_io_pipe_phv_out_data_180; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_181 = pipe3to8_io_pipe_phv_out_data_181; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_182 = pipe3to8_io_pipe_phv_out_data_182; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_183 = pipe3to8_io_pipe_phv_out_data_183; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_184 = pipe3to8_io_pipe_phv_out_data_184; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_185 = pipe3to8_io_pipe_phv_out_data_185; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_186 = pipe3to8_io_pipe_phv_out_data_186; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_187 = pipe3to8_io_pipe_phv_out_data_187; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_188 = pipe3to8_io_pipe_phv_out_data_188; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_189 = pipe3to8_io_pipe_phv_out_data_189; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_190 = pipe3to8_io_pipe_phv_out_data_190; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_191 = pipe3to8_io_pipe_phv_out_data_191; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_192 = pipe3to8_io_pipe_phv_out_data_192; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_193 = pipe3to8_io_pipe_phv_out_data_193; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_194 = pipe3to8_io_pipe_phv_out_data_194; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_195 = pipe3to8_io_pipe_phv_out_data_195; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_196 = pipe3to8_io_pipe_phv_out_data_196; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_197 = pipe3to8_io_pipe_phv_out_data_197; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_198 = pipe3to8_io_pipe_phv_out_data_198; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_199 = pipe3to8_io_pipe_phv_out_data_199; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_200 = pipe3to8_io_pipe_phv_out_data_200; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_201 = pipe3to8_io_pipe_phv_out_data_201; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_202 = pipe3to8_io_pipe_phv_out_data_202; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_203 = pipe3to8_io_pipe_phv_out_data_203; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_204 = pipe3to8_io_pipe_phv_out_data_204; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_205 = pipe3to8_io_pipe_phv_out_data_205; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_206 = pipe3to8_io_pipe_phv_out_data_206; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_207 = pipe3to8_io_pipe_phv_out_data_207; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_208 = pipe3to8_io_pipe_phv_out_data_208; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_209 = pipe3to8_io_pipe_phv_out_data_209; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_210 = pipe3to8_io_pipe_phv_out_data_210; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_211 = pipe3to8_io_pipe_phv_out_data_211; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_212 = pipe3to8_io_pipe_phv_out_data_212; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_213 = pipe3to8_io_pipe_phv_out_data_213; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_214 = pipe3to8_io_pipe_phv_out_data_214; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_215 = pipe3to8_io_pipe_phv_out_data_215; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_216 = pipe3to8_io_pipe_phv_out_data_216; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_217 = pipe3to8_io_pipe_phv_out_data_217; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_218 = pipe3to8_io_pipe_phv_out_data_218; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_219 = pipe3to8_io_pipe_phv_out_data_219; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_220 = pipe3to8_io_pipe_phv_out_data_220; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_221 = pipe3to8_io_pipe_phv_out_data_221; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_222 = pipe3to8_io_pipe_phv_out_data_222; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_223 = pipe3to8_io_pipe_phv_out_data_223; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_224 = pipe3to8_io_pipe_phv_out_data_224; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_225 = pipe3to8_io_pipe_phv_out_data_225; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_226 = pipe3to8_io_pipe_phv_out_data_226; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_227 = pipe3to8_io_pipe_phv_out_data_227; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_228 = pipe3to8_io_pipe_phv_out_data_228; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_229 = pipe3to8_io_pipe_phv_out_data_229; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_230 = pipe3to8_io_pipe_phv_out_data_230; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_231 = pipe3to8_io_pipe_phv_out_data_231; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_232 = pipe3to8_io_pipe_phv_out_data_232; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_233 = pipe3to8_io_pipe_phv_out_data_233; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_234 = pipe3to8_io_pipe_phv_out_data_234; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_235 = pipe3to8_io_pipe_phv_out_data_235; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_236 = pipe3to8_io_pipe_phv_out_data_236; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_237 = pipe3to8_io_pipe_phv_out_data_237; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_238 = pipe3to8_io_pipe_phv_out_data_238; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_239 = pipe3to8_io_pipe_phv_out_data_239; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_240 = pipe3to8_io_pipe_phv_out_data_240; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_241 = pipe3to8_io_pipe_phv_out_data_241; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_242 = pipe3to8_io_pipe_phv_out_data_242; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_243 = pipe3to8_io_pipe_phv_out_data_243; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_244 = pipe3to8_io_pipe_phv_out_data_244; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_245 = pipe3to8_io_pipe_phv_out_data_245; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_246 = pipe3to8_io_pipe_phv_out_data_246; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_247 = pipe3to8_io_pipe_phv_out_data_247; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_248 = pipe3to8_io_pipe_phv_out_data_248; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_249 = pipe3to8_io_pipe_phv_out_data_249; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_250 = pipe3to8_io_pipe_phv_out_data_250; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_251 = pipe3to8_io_pipe_phv_out_data_251; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_252 = pipe3to8_io_pipe_phv_out_data_252; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_253 = pipe3to8_io_pipe_phv_out_data_253; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_254 = pipe3to8_io_pipe_phv_out_data_254; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_255 = pipe3to8_io_pipe_phv_out_data_255; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_0 = pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_1 = pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_2 = pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_3 = pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_4 = pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_5 = pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_6 = pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_7 = pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_8 = pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_9 = pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_10 = pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_11 = pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_12 = pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_13 = pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_14 = pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_15 = pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_current_state = pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_current_offset = pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_transition_field = pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_next_processor_id = pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_next_config_id = pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_is_valid_processor = pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 364:27]
  assign pipe9_io_table_config_0_sram_id_table_0 = table_config_0_sram_id_table_0; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_1 = table_config_0_sram_id_table_1; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_2 = table_config_0_sram_id_table_2; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_3 = table_config_0_sram_id_table_3; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_4 = table_config_0_sram_id_table_4; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_5 = table_config_0_sram_id_table_5; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_6 = table_config_0_sram_id_table_6; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_7 = table_config_0_sram_id_table_7; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_8 = table_config_0_sram_id_table_8; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_9 = table_config_0_sram_id_table_9; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_10 = table_config_0_sram_id_table_10; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_11 = table_config_0_sram_id_table_11; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_12 = table_config_0_sram_id_table_12; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_13 = table_config_0_sram_id_table_13; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_14 = table_config_0_sram_id_table_14; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_15 = table_config_0_sram_id_table_15; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_16 = table_config_0_sram_id_table_16; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_17 = table_config_0_sram_id_table_17; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_18 = table_config_0_sram_id_table_18; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_19 = table_config_0_sram_id_table_19; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_20 = table_config_0_sram_id_table_20; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_21 = table_config_0_sram_id_table_21; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_22 = table_config_0_sram_id_table_22; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_23 = table_config_0_sram_id_table_23; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_24 = table_config_0_sram_id_table_24; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_25 = table_config_0_sram_id_table_25; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_26 = table_config_0_sram_id_table_26; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_27 = table_config_0_sram_id_table_27; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_28 = table_config_0_sram_id_table_28; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_29 = table_config_0_sram_id_table_29; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_30 = table_config_0_sram_id_table_30; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_31 = table_config_0_sram_id_table_31; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_32 = table_config_0_sram_id_table_32; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_33 = table_config_0_sram_id_table_33; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_34 = table_config_0_sram_id_table_34; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_35 = table_config_0_sram_id_table_35; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_36 = table_config_0_sram_id_table_36; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_37 = table_config_0_sram_id_table_37; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_38 = table_config_0_sram_id_table_38; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_39 = table_config_0_sram_id_table_39; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_40 = table_config_0_sram_id_table_40; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_41 = table_config_0_sram_id_table_41; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_42 = table_config_0_sram_id_table_42; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_43 = table_config_0_sram_id_table_43; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_44 = table_config_0_sram_id_table_44; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_45 = table_config_0_sram_id_table_45; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_46 = table_config_0_sram_id_table_46; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_47 = table_config_0_sram_id_table_47; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_48 = table_config_0_sram_id_table_48; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_49 = table_config_0_sram_id_table_49; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_50 = table_config_0_sram_id_table_50; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_51 = table_config_0_sram_id_table_51; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_52 = table_config_0_sram_id_table_52; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_53 = table_config_0_sram_id_table_53; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_54 = table_config_0_sram_id_table_54; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_55 = table_config_0_sram_id_table_55; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_56 = table_config_0_sram_id_table_56; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_57 = table_config_0_sram_id_table_57; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_58 = table_config_0_sram_id_table_58; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_59 = table_config_0_sram_id_table_59; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_60 = table_config_0_sram_id_table_60; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_61 = table_config_0_sram_id_table_61; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_62 = table_config_0_sram_id_table_62; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_sram_id_table_63 = table_config_0_sram_id_table_63; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_0 = table_config_1_sram_id_table_0; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_1 = table_config_1_sram_id_table_1; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_2 = table_config_1_sram_id_table_2; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_3 = table_config_1_sram_id_table_3; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_4 = table_config_1_sram_id_table_4; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_5 = table_config_1_sram_id_table_5; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_6 = table_config_1_sram_id_table_6; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_7 = table_config_1_sram_id_table_7; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_8 = table_config_1_sram_id_table_8; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_9 = table_config_1_sram_id_table_9; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_10 = table_config_1_sram_id_table_10; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_11 = table_config_1_sram_id_table_11; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_12 = table_config_1_sram_id_table_12; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_13 = table_config_1_sram_id_table_13; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_14 = table_config_1_sram_id_table_14; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_15 = table_config_1_sram_id_table_15; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_16 = table_config_1_sram_id_table_16; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_17 = table_config_1_sram_id_table_17; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_18 = table_config_1_sram_id_table_18; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_19 = table_config_1_sram_id_table_19; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_20 = table_config_1_sram_id_table_20; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_21 = table_config_1_sram_id_table_21; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_22 = table_config_1_sram_id_table_22; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_23 = table_config_1_sram_id_table_23; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_24 = table_config_1_sram_id_table_24; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_25 = table_config_1_sram_id_table_25; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_26 = table_config_1_sram_id_table_26; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_27 = table_config_1_sram_id_table_27; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_28 = table_config_1_sram_id_table_28; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_29 = table_config_1_sram_id_table_29; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_30 = table_config_1_sram_id_table_30; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_31 = table_config_1_sram_id_table_31; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_32 = table_config_1_sram_id_table_32; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_33 = table_config_1_sram_id_table_33; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_34 = table_config_1_sram_id_table_34; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_35 = table_config_1_sram_id_table_35; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_36 = table_config_1_sram_id_table_36; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_37 = table_config_1_sram_id_table_37; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_38 = table_config_1_sram_id_table_38; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_39 = table_config_1_sram_id_table_39; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_40 = table_config_1_sram_id_table_40; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_41 = table_config_1_sram_id_table_41; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_42 = table_config_1_sram_id_table_42; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_43 = table_config_1_sram_id_table_43; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_44 = table_config_1_sram_id_table_44; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_45 = table_config_1_sram_id_table_45; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_46 = table_config_1_sram_id_table_46; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_47 = table_config_1_sram_id_table_47; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_48 = table_config_1_sram_id_table_48; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_49 = table_config_1_sram_id_table_49; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_50 = table_config_1_sram_id_table_50; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_51 = table_config_1_sram_id_table_51; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_52 = table_config_1_sram_id_table_52; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_53 = table_config_1_sram_id_table_53; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_54 = table_config_1_sram_id_table_54; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_55 = table_config_1_sram_id_table_55; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_56 = table_config_1_sram_id_table_56; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_57 = table_config_1_sram_id_table_57; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_58 = table_config_1_sram_id_table_58; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_59 = table_config_1_sram_id_table_59; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_60 = table_config_1_sram_id_table_60; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_61 = table_config_1_sram_id_table_61; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_62 = table_config_1_sram_id_table_62; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_sram_id_table_63 = table_config_1_sram_id_table_63; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 368:27]
  assign pipe9_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 368:27]
  assign pipe9_io_key_in = pipe3to8_io_key_out; // @[matcher.scala 365:27]
  assign pipe9_io_addr_in = pipe3to8_io_hash_val; // @[matcher.scala 366:27]
  assign pipe9_io_cs_in = pipe3to8_io_hash_val_cs; // @[matcher.scala 367:27]
  assign pipe10_clock = clock;
  assign pipe10_io_pipe_phv_in_data_0 = pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_1 = pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_2 = pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_3 = pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_4 = pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_5 = pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_6 = pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_7 = pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_8 = pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_9 = pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_10 = pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_11 = pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_12 = pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_13 = pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_14 = pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_15 = pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_16 = pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_17 = pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_18 = pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_19 = pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_20 = pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_21 = pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_22 = pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_23 = pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_24 = pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_25 = pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_26 = pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_27 = pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_28 = pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_29 = pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_30 = pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_31 = pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_32 = pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_33 = pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_34 = pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_35 = pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_36 = pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_37 = pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_38 = pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_39 = pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_40 = pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_41 = pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_42 = pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_43 = pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_44 = pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_45 = pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_46 = pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_47 = pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_48 = pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_49 = pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_50 = pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_51 = pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_52 = pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_53 = pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_54 = pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_55 = pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_56 = pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_57 = pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_58 = pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_59 = pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_60 = pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_61 = pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_62 = pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_63 = pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_64 = pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_65 = pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_66 = pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_67 = pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_68 = pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_69 = pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_70 = pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_71 = pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_72 = pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_73 = pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_74 = pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_75 = pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_76 = pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_77 = pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_78 = pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_79 = pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_80 = pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_81 = pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_82 = pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_83 = pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_84 = pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_85 = pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_86 = pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_87 = pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_88 = pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_89 = pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_90 = pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_91 = pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_92 = pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_93 = pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_94 = pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_95 = pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_96 = pipe9_io_pipe_phv_out_data_96; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_97 = pipe9_io_pipe_phv_out_data_97; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_98 = pipe9_io_pipe_phv_out_data_98; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_99 = pipe9_io_pipe_phv_out_data_99; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_100 = pipe9_io_pipe_phv_out_data_100; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_101 = pipe9_io_pipe_phv_out_data_101; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_102 = pipe9_io_pipe_phv_out_data_102; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_103 = pipe9_io_pipe_phv_out_data_103; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_104 = pipe9_io_pipe_phv_out_data_104; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_105 = pipe9_io_pipe_phv_out_data_105; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_106 = pipe9_io_pipe_phv_out_data_106; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_107 = pipe9_io_pipe_phv_out_data_107; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_108 = pipe9_io_pipe_phv_out_data_108; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_109 = pipe9_io_pipe_phv_out_data_109; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_110 = pipe9_io_pipe_phv_out_data_110; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_111 = pipe9_io_pipe_phv_out_data_111; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_112 = pipe9_io_pipe_phv_out_data_112; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_113 = pipe9_io_pipe_phv_out_data_113; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_114 = pipe9_io_pipe_phv_out_data_114; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_115 = pipe9_io_pipe_phv_out_data_115; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_116 = pipe9_io_pipe_phv_out_data_116; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_117 = pipe9_io_pipe_phv_out_data_117; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_118 = pipe9_io_pipe_phv_out_data_118; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_119 = pipe9_io_pipe_phv_out_data_119; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_120 = pipe9_io_pipe_phv_out_data_120; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_121 = pipe9_io_pipe_phv_out_data_121; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_122 = pipe9_io_pipe_phv_out_data_122; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_123 = pipe9_io_pipe_phv_out_data_123; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_124 = pipe9_io_pipe_phv_out_data_124; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_125 = pipe9_io_pipe_phv_out_data_125; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_126 = pipe9_io_pipe_phv_out_data_126; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_127 = pipe9_io_pipe_phv_out_data_127; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_128 = pipe9_io_pipe_phv_out_data_128; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_129 = pipe9_io_pipe_phv_out_data_129; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_130 = pipe9_io_pipe_phv_out_data_130; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_131 = pipe9_io_pipe_phv_out_data_131; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_132 = pipe9_io_pipe_phv_out_data_132; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_133 = pipe9_io_pipe_phv_out_data_133; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_134 = pipe9_io_pipe_phv_out_data_134; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_135 = pipe9_io_pipe_phv_out_data_135; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_136 = pipe9_io_pipe_phv_out_data_136; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_137 = pipe9_io_pipe_phv_out_data_137; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_138 = pipe9_io_pipe_phv_out_data_138; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_139 = pipe9_io_pipe_phv_out_data_139; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_140 = pipe9_io_pipe_phv_out_data_140; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_141 = pipe9_io_pipe_phv_out_data_141; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_142 = pipe9_io_pipe_phv_out_data_142; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_143 = pipe9_io_pipe_phv_out_data_143; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_144 = pipe9_io_pipe_phv_out_data_144; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_145 = pipe9_io_pipe_phv_out_data_145; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_146 = pipe9_io_pipe_phv_out_data_146; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_147 = pipe9_io_pipe_phv_out_data_147; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_148 = pipe9_io_pipe_phv_out_data_148; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_149 = pipe9_io_pipe_phv_out_data_149; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_150 = pipe9_io_pipe_phv_out_data_150; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_151 = pipe9_io_pipe_phv_out_data_151; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_152 = pipe9_io_pipe_phv_out_data_152; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_153 = pipe9_io_pipe_phv_out_data_153; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_154 = pipe9_io_pipe_phv_out_data_154; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_155 = pipe9_io_pipe_phv_out_data_155; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_156 = pipe9_io_pipe_phv_out_data_156; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_157 = pipe9_io_pipe_phv_out_data_157; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_158 = pipe9_io_pipe_phv_out_data_158; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_159 = pipe9_io_pipe_phv_out_data_159; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_160 = pipe9_io_pipe_phv_out_data_160; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_161 = pipe9_io_pipe_phv_out_data_161; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_162 = pipe9_io_pipe_phv_out_data_162; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_163 = pipe9_io_pipe_phv_out_data_163; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_164 = pipe9_io_pipe_phv_out_data_164; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_165 = pipe9_io_pipe_phv_out_data_165; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_166 = pipe9_io_pipe_phv_out_data_166; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_167 = pipe9_io_pipe_phv_out_data_167; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_168 = pipe9_io_pipe_phv_out_data_168; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_169 = pipe9_io_pipe_phv_out_data_169; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_170 = pipe9_io_pipe_phv_out_data_170; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_171 = pipe9_io_pipe_phv_out_data_171; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_172 = pipe9_io_pipe_phv_out_data_172; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_173 = pipe9_io_pipe_phv_out_data_173; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_174 = pipe9_io_pipe_phv_out_data_174; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_175 = pipe9_io_pipe_phv_out_data_175; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_176 = pipe9_io_pipe_phv_out_data_176; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_177 = pipe9_io_pipe_phv_out_data_177; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_178 = pipe9_io_pipe_phv_out_data_178; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_179 = pipe9_io_pipe_phv_out_data_179; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_180 = pipe9_io_pipe_phv_out_data_180; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_181 = pipe9_io_pipe_phv_out_data_181; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_182 = pipe9_io_pipe_phv_out_data_182; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_183 = pipe9_io_pipe_phv_out_data_183; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_184 = pipe9_io_pipe_phv_out_data_184; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_185 = pipe9_io_pipe_phv_out_data_185; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_186 = pipe9_io_pipe_phv_out_data_186; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_187 = pipe9_io_pipe_phv_out_data_187; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_188 = pipe9_io_pipe_phv_out_data_188; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_189 = pipe9_io_pipe_phv_out_data_189; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_190 = pipe9_io_pipe_phv_out_data_190; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_191 = pipe9_io_pipe_phv_out_data_191; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_192 = pipe9_io_pipe_phv_out_data_192; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_193 = pipe9_io_pipe_phv_out_data_193; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_194 = pipe9_io_pipe_phv_out_data_194; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_195 = pipe9_io_pipe_phv_out_data_195; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_196 = pipe9_io_pipe_phv_out_data_196; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_197 = pipe9_io_pipe_phv_out_data_197; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_198 = pipe9_io_pipe_phv_out_data_198; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_199 = pipe9_io_pipe_phv_out_data_199; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_200 = pipe9_io_pipe_phv_out_data_200; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_201 = pipe9_io_pipe_phv_out_data_201; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_202 = pipe9_io_pipe_phv_out_data_202; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_203 = pipe9_io_pipe_phv_out_data_203; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_204 = pipe9_io_pipe_phv_out_data_204; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_205 = pipe9_io_pipe_phv_out_data_205; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_206 = pipe9_io_pipe_phv_out_data_206; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_207 = pipe9_io_pipe_phv_out_data_207; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_208 = pipe9_io_pipe_phv_out_data_208; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_209 = pipe9_io_pipe_phv_out_data_209; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_210 = pipe9_io_pipe_phv_out_data_210; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_211 = pipe9_io_pipe_phv_out_data_211; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_212 = pipe9_io_pipe_phv_out_data_212; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_213 = pipe9_io_pipe_phv_out_data_213; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_214 = pipe9_io_pipe_phv_out_data_214; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_215 = pipe9_io_pipe_phv_out_data_215; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_216 = pipe9_io_pipe_phv_out_data_216; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_217 = pipe9_io_pipe_phv_out_data_217; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_218 = pipe9_io_pipe_phv_out_data_218; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_219 = pipe9_io_pipe_phv_out_data_219; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_220 = pipe9_io_pipe_phv_out_data_220; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_221 = pipe9_io_pipe_phv_out_data_221; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_222 = pipe9_io_pipe_phv_out_data_222; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_223 = pipe9_io_pipe_phv_out_data_223; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_224 = pipe9_io_pipe_phv_out_data_224; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_225 = pipe9_io_pipe_phv_out_data_225; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_226 = pipe9_io_pipe_phv_out_data_226; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_227 = pipe9_io_pipe_phv_out_data_227; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_228 = pipe9_io_pipe_phv_out_data_228; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_229 = pipe9_io_pipe_phv_out_data_229; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_230 = pipe9_io_pipe_phv_out_data_230; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_231 = pipe9_io_pipe_phv_out_data_231; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_232 = pipe9_io_pipe_phv_out_data_232; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_233 = pipe9_io_pipe_phv_out_data_233; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_234 = pipe9_io_pipe_phv_out_data_234; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_235 = pipe9_io_pipe_phv_out_data_235; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_236 = pipe9_io_pipe_phv_out_data_236; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_237 = pipe9_io_pipe_phv_out_data_237; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_238 = pipe9_io_pipe_phv_out_data_238; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_239 = pipe9_io_pipe_phv_out_data_239; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_240 = pipe9_io_pipe_phv_out_data_240; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_241 = pipe9_io_pipe_phv_out_data_241; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_242 = pipe9_io_pipe_phv_out_data_242; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_243 = pipe9_io_pipe_phv_out_data_243; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_244 = pipe9_io_pipe_phv_out_data_244; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_245 = pipe9_io_pipe_phv_out_data_245; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_246 = pipe9_io_pipe_phv_out_data_246; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_247 = pipe9_io_pipe_phv_out_data_247; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_248 = pipe9_io_pipe_phv_out_data_248; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_249 = pipe9_io_pipe_phv_out_data_249; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_250 = pipe9_io_pipe_phv_out_data_250; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_251 = pipe9_io_pipe_phv_out_data_251; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_252 = pipe9_io_pipe_phv_out_data_252; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_253 = pipe9_io_pipe_phv_out_data_253; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_254 = pipe9_io_pipe_phv_out_data_254; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_255 = pipe9_io_pipe_phv_out_data_255; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_0 = pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_1 = pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_2 = pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_3 = pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_4 = pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_5 = pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_6 = pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_7 = pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_8 = pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_9 = pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_10 = pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_11 = pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_12 = pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_13 = pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_14 = pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_15 = pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_current_state = pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_current_offset = pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_transition_field = pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_next_processor_id = pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_next_config_id = pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_is_valid_processor = pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 370:27]
  assign pipe10_io_key_in = pipe9_io_key_out; // @[matcher.scala 371:27]
  assign pipe10_io_cs_in = pipe9_io_cs_out; // @[matcher.scala 372:27]
  assign pipe10_io_addr_in = pipe9_io_addr_out; // @[matcher.scala 373:27]
  assign pipe10_io_cs_vec_in_0 = pipe9_io_cs_vec_out_0; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_1 = pipe9_io_cs_vec_out_1; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_2 = pipe9_io_cs_vec_out_2; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_3 = pipe9_io_cs_vec_out_3; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_4 = pipe9_io_cs_vec_out_4; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_5 = pipe9_io_cs_vec_out_5; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_6 = pipe9_io_cs_vec_out_6; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_7 = pipe9_io_cs_vec_out_7; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_8 = pipe9_io_cs_vec_out_8; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_9 = pipe9_io_cs_vec_out_9; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_10 = pipe9_io_cs_vec_out_10; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_11 = pipe9_io_cs_vec_out_11; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_12 = pipe9_io_cs_vec_out_12; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_13 = pipe9_io_cs_vec_out_13; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_14 = pipe9_io_cs_vec_out_14; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_15 = pipe9_io_cs_vec_out_15; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_16 = pipe9_io_cs_vec_out_16; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_17 = pipe9_io_cs_vec_out_17; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_18 = pipe9_io_cs_vec_out_18; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_19 = pipe9_io_cs_vec_out_19; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_20 = pipe9_io_cs_vec_out_20; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_21 = pipe9_io_cs_vec_out_21; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_22 = pipe9_io_cs_vec_out_22; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_23 = pipe9_io_cs_vec_out_23; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_24 = pipe9_io_cs_vec_out_24; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_25 = pipe9_io_cs_vec_out_25; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_26 = pipe9_io_cs_vec_out_26; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_27 = pipe9_io_cs_vec_out_27; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_28 = pipe9_io_cs_vec_out_28; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_29 = pipe9_io_cs_vec_out_29; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_30 = pipe9_io_cs_vec_out_30; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_31 = pipe9_io_cs_vec_out_31; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_32 = pipe9_io_cs_vec_out_32; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_33 = pipe9_io_cs_vec_out_33; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_34 = pipe9_io_cs_vec_out_34; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_35 = pipe9_io_cs_vec_out_35; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_36 = pipe9_io_cs_vec_out_36; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_37 = pipe9_io_cs_vec_out_37; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_38 = pipe9_io_cs_vec_out_38; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_39 = pipe9_io_cs_vec_out_39; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_40 = pipe9_io_cs_vec_out_40; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_41 = pipe9_io_cs_vec_out_41; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_42 = pipe9_io_cs_vec_out_42; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_43 = pipe9_io_cs_vec_out_43; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_44 = pipe9_io_cs_vec_out_44; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_45 = pipe9_io_cs_vec_out_45; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_46 = pipe9_io_cs_vec_out_46; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_47 = pipe9_io_cs_vec_out_47; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_48 = pipe9_io_cs_vec_out_48; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_49 = pipe9_io_cs_vec_out_49; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_50 = pipe9_io_cs_vec_out_50; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_51 = pipe9_io_cs_vec_out_51; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_52 = pipe9_io_cs_vec_out_52; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_53 = pipe9_io_cs_vec_out_53; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_54 = pipe9_io_cs_vec_out_54; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_55 = pipe9_io_cs_vec_out_55; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_56 = pipe9_io_cs_vec_out_56; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_57 = pipe9_io_cs_vec_out_57; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_58 = pipe9_io_cs_vec_out_58; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_59 = pipe9_io_cs_vec_out_59; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_60 = pipe9_io_cs_vec_out_60; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_61 = pipe9_io_cs_vec_out_61; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_62 = pipe9_io_cs_vec_out_62; // @[matcher.scala 374:27]
  assign pipe10_io_cs_vec_in_63 = pipe9_io_cs_vec_out_63; // @[matcher.scala 374:27]
  assign pipe10_io_mem_cluster_0_data = io_mem_cluster_0_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_1_data = io_mem_cluster_1_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_2_data = io_mem_cluster_2_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_3_data = io_mem_cluster_3_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_4_data = io_mem_cluster_4_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_5_data = io_mem_cluster_5_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_6_data = io_mem_cluster_6_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_7_data = io_mem_cluster_7_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_8_data = io_mem_cluster_8_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_9_data = io_mem_cluster_9_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_10_data = io_mem_cluster_10_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_11_data = io_mem_cluster_11_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_12_data = io_mem_cluster_12_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_13_data = io_mem_cluster_13_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_14_data = io_mem_cluster_14_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_15_data = io_mem_cluster_15_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_16_data = io_mem_cluster_16_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_17_data = io_mem_cluster_17_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_18_data = io_mem_cluster_18_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_19_data = io_mem_cluster_19_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_20_data = io_mem_cluster_20_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_21_data = io_mem_cluster_21_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_22_data = io_mem_cluster_22_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_23_data = io_mem_cluster_23_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_24_data = io_mem_cluster_24_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_25_data = io_mem_cluster_25_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_26_data = io_mem_cluster_26_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_27_data = io_mem_cluster_27_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_28_data = io_mem_cluster_28_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_29_data = io_mem_cluster_29_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_30_data = io_mem_cluster_30_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_31_data = io_mem_cluster_31_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_32_data = io_mem_cluster_32_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_33_data = io_mem_cluster_33_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_34_data = io_mem_cluster_34_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_35_data = io_mem_cluster_35_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_36_data = io_mem_cluster_36_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_37_data = io_mem_cluster_37_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_38_data = io_mem_cluster_38_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_39_data = io_mem_cluster_39_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_40_data = io_mem_cluster_40_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_41_data = io_mem_cluster_41_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_42_data = io_mem_cluster_42_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_43_data = io_mem_cluster_43_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_44_data = io_mem_cluster_44_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_45_data = io_mem_cluster_45_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_46_data = io_mem_cluster_46_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_47_data = io_mem_cluster_47_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_48_data = io_mem_cluster_48_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_49_data = io_mem_cluster_49_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_50_data = io_mem_cluster_50_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_51_data = io_mem_cluster_51_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_52_data = io_mem_cluster_52_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_53_data = io_mem_cluster_53_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_54_data = io_mem_cluster_54_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_55_data = io_mem_cluster_55_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_56_data = io_mem_cluster_56_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_57_data = io_mem_cluster_57_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_58_data = io_mem_cluster_58_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_59_data = io_mem_cluster_59_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_60_data = io_mem_cluster_60_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_61_data = io_mem_cluster_61_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_62_data = io_mem_cluster_62_data; // @[matcher.scala 375:27]
  assign pipe10_io_mem_cluster_63_data = io_mem_cluster_63_data; // @[matcher.scala 375:27]
  assign pipe11_clock = clock;
  assign pipe11_io_pipe_phv_in_data_0 = pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_1 = pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_2 = pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_3 = pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_4 = pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_5 = pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_6 = pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_7 = pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_8 = pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_9 = pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_10 = pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_11 = pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_12 = pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_13 = pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_14 = pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_15 = pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_16 = pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_17 = pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_18 = pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_19 = pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_20 = pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_21 = pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_22 = pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_23 = pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_24 = pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_25 = pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_26 = pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_27 = pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_28 = pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_29 = pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_30 = pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_31 = pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_32 = pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_33 = pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_34 = pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_35 = pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_36 = pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_37 = pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_38 = pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_39 = pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_40 = pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_41 = pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_42 = pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_43 = pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_44 = pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_45 = pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_46 = pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_47 = pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_48 = pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_49 = pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_50 = pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_51 = pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_52 = pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_53 = pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_54 = pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_55 = pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_56 = pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_57 = pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_58 = pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_59 = pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_60 = pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_61 = pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_62 = pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_63 = pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_64 = pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_65 = pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_66 = pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_67 = pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_68 = pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_69 = pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_70 = pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_71 = pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_72 = pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_73 = pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_74 = pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_75 = pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_76 = pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_77 = pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_78 = pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_79 = pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_80 = pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_81 = pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_82 = pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_83 = pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_84 = pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_85 = pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_86 = pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_87 = pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_88 = pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_89 = pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_90 = pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_91 = pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_92 = pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_93 = pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_94 = pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_95 = pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_96 = pipe10_io_pipe_phv_out_data_96; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_97 = pipe10_io_pipe_phv_out_data_97; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_98 = pipe10_io_pipe_phv_out_data_98; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_99 = pipe10_io_pipe_phv_out_data_99; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_100 = pipe10_io_pipe_phv_out_data_100; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_101 = pipe10_io_pipe_phv_out_data_101; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_102 = pipe10_io_pipe_phv_out_data_102; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_103 = pipe10_io_pipe_phv_out_data_103; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_104 = pipe10_io_pipe_phv_out_data_104; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_105 = pipe10_io_pipe_phv_out_data_105; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_106 = pipe10_io_pipe_phv_out_data_106; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_107 = pipe10_io_pipe_phv_out_data_107; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_108 = pipe10_io_pipe_phv_out_data_108; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_109 = pipe10_io_pipe_phv_out_data_109; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_110 = pipe10_io_pipe_phv_out_data_110; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_111 = pipe10_io_pipe_phv_out_data_111; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_112 = pipe10_io_pipe_phv_out_data_112; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_113 = pipe10_io_pipe_phv_out_data_113; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_114 = pipe10_io_pipe_phv_out_data_114; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_115 = pipe10_io_pipe_phv_out_data_115; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_116 = pipe10_io_pipe_phv_out_data_116; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_117 = pipe10_io_pipe_phv_out_data_117; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_118 = pipe10_io_pipe_phv_out_data_118; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_119 = pipe10_io_pipe_phv_out_data_119; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_120 = pipe10_io_pipe_phv_out_data_120; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_121 = pipe10_io_pipe_phv_out_data_121; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_122 = pipe10_io_pipe_phv_out_data_122; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_123 = pipe10_io_pipe_phv_out_data_123; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_124 = pipe10_io_pipe_phv_out_data_124; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_125 = pipe10_io_pipe_phv_out_data_125; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_126 = pipe10_io_pipe_phv_out_data_126; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_127 = pipe10_io_pipe_phv_out_data_127; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_128 = pipe10_io_pipe_phv_out_data_128; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_129 = pipe10_io_pipe_phv_out_data_129; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_130 = pipe10_io_pipe_phv_out_data_130; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_131 = pipe10_io_pipe_phv_out_data_131; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_132 = pipe10_io_pipe_phv_out_data_132; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_133 = pipe10_io_pipe_phv_out_data_133; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_134 = pipe10_io_pipe_phv_out_data_134; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_135 = pipe10_io_pipe_phv_out_data_135; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_136 = pipe10_io_pipe_phv_out_data_136; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_137 = pipe10_io_pipe_phv_out_data_137; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_138 = pipe10_io_pipe_phv_out_data_138; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_139 = pipe10_io_pipe_phv_out_data_139; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_140 = pipe10_io_pipe_phv_out_data_140; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_141 = pipe10_io_pipe_phv_out_data_141; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_142 = pipe10_io_pipe_phv_out_data_142; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_143 = pipe10_io_pipe_phv_out_data_143; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_144 = pipe10_io_pipe_phv_out_data_144; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_145 = pipe10_io_pipe_phv_out_data_145; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_146 = pipe10_io_pipe_phv_out_data_146; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_147 = pipe10_io_pipe_phv_out_data_147; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_148 = pipe10_io_pipe_phv_out_data_148; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_149 = pipe10_io_pipe_phv_out_data_149; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_150 = pipe10_io_pipe_phv_out_data_150; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_151 = pipe10_io_pipe_phv_out_data_151; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_152 = pipe10_io_pipe_phv_out_data_152; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_153 = pipe10_io_pipe_phv_out_data_153; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_154 = pipe10_io_pipe_phv_out_data_154; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_155 = pipe10_io_pipe_phv_out_data_155; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_156 = pipe10_io_pipe_phv_out_data_156; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_157 = pipe10_io_pipe_phv_out_data_157; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_158 = pipe10_io_pipe_phv_out_data_158; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_159 = pipe10_io_pipe_phv_out_data_159; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_160 = pipe10_io_pipe_phv_out_data_160; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_161 = pipe10_io_pipe_phv_out_data_161; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_162 = pipe10_io_pipe_phv_out_data_162; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_163 = pipe10_io_pipe_phv_out_data_163; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_164 = pipe10_io_pipe_phv_out_data_164; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_165 = pipe10_io_pipe_phv_out_data_165; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_166 = pipe10_io_pipe_phv_out_data_166; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_167 = pipe10_io_pipe_phv_out_data_167; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_168 = pipe10_io_pipe_phv_out_data_168; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_169 = pipe10_io_pipe_phv_out_data_169; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_170 = pipe10_io_pipe_phv_out_data_170; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_171 = pipe10_io_pipe_phv_out_data_171; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_172 = pipe10_io_pipe_phv_out_data_172; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_173 = pipe10_io_pipe_phv_out_data_173; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_174 = pipe10_io_pipe_phv_out_data_174; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_175 = pipe10_io_pipe_phv_out_data_175; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_176 = pipe10_io_pipe_phv_out_data_176; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_177 = pipe10_io_pipe_phv_out_data_177; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_178 = pipe10_io_pipe_phv_out_data_178; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_179 = pipe10_io_pipe_phv_out_data_179; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_180 = pipe10_io_pipe_phv_out_data_180; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_181 = pipe10_io_pipe_phv_out_data_181; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_182 = pipe10_io_pipe_phv_out_data_182; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_183 = pipe10_io_pipe_phv_out_data_183; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_184 = pipe10_io_pipe_phv_out_data_184; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_185 = pipe10_io_pipe_phv_out_data_185; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_186 = pipe10_io_pipe_phv_out_data_186; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_187 = pipe10_io_pipe_phv_out_data_187; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_188 = pipe10_io_pipe_phv_out_data_188; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_189 = pipe10_io_pipe_phv_out_data_189; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_190 = pipe10_io_pipe_phv_out_data_190; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_191 = pipe10_io_pipe_phv_out_data_191; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_192 = pipe10_io_pipe_phv_out_data_192; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_193 = pipe10_io_pipe_phv_out_data_193; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_194 = pipe10_io_pipe_phv_out_data_194; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_195 = pipe10_io_pipe_phv_out_data_195; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_196 = pipe10_io_pipe_phv_out_data_196; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_197 = pipe10_io_pipe_phv_out_data_197; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_198 = pipe10_io_pipe_phv_out_data_198; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_199 = pipe10_io_pipe_phv_out_data_199; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_200 = pipe10_io_pipe_phv_out_data_200; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_201 = pipe10_io_pipe_phv_out_data_201; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_202 = pipe10_io_pipe_phv_out_data_202; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_203 = pipe10_io_pipe_phv_out_data_203; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_204 = pipe10_io_pipe_phv_out_data_204; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_205 = pipe10_io_pipe_phv_out_data_205; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_206 = pipe10_io_pipe_phv_out_data_206; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_207 = pipe10_io_pipe_phv_out_data_207; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_208 = pipe10_io_pipe_phv_out_data_208; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_209 = pipe10_io_pipe_phv_out_data_209; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_210 = pipe10_io_pipe_phv_out_data_210; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_211 = pipe10_io_pipe_phv_out_data_211; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_212 = pipe10_io_pipe_phv_out_data_212; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_213 = pipe10_io_pipe_phv_out_data_213; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_214 = pipe10_io_pipe_phv_out_data_214; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_215 = pipe10_io_pipe_phv_out_data_215; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_216 = pipe10_io_pipe_phv_out_data_216; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_217 = pipe10_io_pipe_phv_out_data_217; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_218 = pipe10_io_pipe_phv_out_data_218; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_219 = pipe10_io_pipe_phv_out_data_219; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_220 = pipe10_io_pipe_phv_out_data_220; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_221 = pipe10_io_pipe_phv_out_data_221; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_222 = pipe10_io_pipe_phv_out_data_222; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_223 = pipe10_io_pipe_phv_out_data_223; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_224 = pipe10_io_pipe_phv_out_data_224; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_225 = pipe10_io_pipe_phv_out_data_225; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_226 = pipe10_io_pipe_phv_out_data_226; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_227 = pipe10_io_pipe_phv_out_data_227; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_228 = pipe10_io_pipe_phv_out_data_228; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_229 = pipe10_io_pipe_phv_out_data_229; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_230 = pipe10_io_pipe_phv_out_data_230; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_231 = pipe10_io_pipe_phv_out_data_231; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_232 = pipe10_io_pipe_phv_out_data_232; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_233 = pipe10_io_pipe_phv_out_data_233; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_234 = pipe10_io_pipe_phv_out_data_234; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_235 = pipe10_io_pipe_phv_out_data_235; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_236 = pipe10_io_pipe_phv_out_data_236; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_237 = pipe10_io_pipe_phv_out_data_237; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_238 = pipe10_io_pipe_phv_out_data_238; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_239 = pipe10_io_pipe_phv_out_data_239; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_240 = pipe10_io_pipe_phv_out_data_240; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_241 = pipe10_io_pipe_phv_out_data_241; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_242 = pipe10_io_pipe_phv_out_data_242; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_243 = pipe10_io_pipe_phv_out_data_243; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_244 = pipe10_io_pipe_phv_out_data_244; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_245 = pipe10_io_pipe_phv_out_data_245; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_246 = pipe10_io_pipe_phv_out_data_246; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_247 = pipe10_io_pipe_phv_out_data_247; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_248 = pipe10_io_pipe_phv_out_data_248; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_249 = pipe10_io_pipe_phv_out_data_249; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_250 = pipe10_io_pipe_phv_out_data_250; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_251 = pipe10_io_pipe_phv_out_data_251; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_252 = pipe10_io_pipe_phv_out_data_252; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_253 = pipe10_io_pipe_phv_out_data_253; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_254 = pipe10_io_pipe_phv_out_data_254; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_255 = pipe10_io_pipe_phv_out_data_255; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_0 = pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_1 = pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_2 = pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_3 = pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_4 = pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_5 = pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_6 = pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_7 = pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_8 = pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_9 = pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_10 = pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_11 = pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_12 = pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_13 = pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_14 = pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_15 = pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_current_state = pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_current_offset = pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_transition_field = pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_next_processor_id = pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_next_config_id = pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_is_valid_processor = pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 377:27]
  assign pipe11_io_table_config_0_table_width = table_config_0_table_width; // @[matcher.scala 381:28]
  assign pipe11_io_table_config_0_table_depth = table_config_0_table_depth; // @[matcher.scala 381:28]
  assign pipe11_io_table_config_1_table_width = table_config_1_table_width; // @[matcher.scala 381:28]
  assign pipe11_io_table_config_1_table_depth = table_config_1_table_depth; // @[matcher.scala 381:28]
  assign pipe11_io_key_in = pipe10_io_key_out; // @[matcher.scala 378:27]
  assign pipe11_io_cs_in = pipe10_io_cs_out; // @[matcher.scala 379:27]
  assign pipe11_io_data_in_0 = pipe10_io_data_out_0; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_1 = pipe10_io_data_out_1; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_2 = pipe10_io_data_out_2; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_3 = pipe10_io_data_out_3; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_4 = pipe10_io_data_out_4; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_5 = pipe10_io_data_out_5; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_6 = pipe10_io_data_out_6; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_7 = pipe10_io_data_out_7; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_8 = pipe10_io_data_out_8; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_9 = pipe10_io_data_out_9; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_10 = pipe10_io_data_out_10; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_11 = pipe10_io_data_out_11; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_12 = pipe10_io_data_out_12; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_13 = pipe10_io_data_out_13; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_14 = pipe10_io_data_out_14; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_15 = pipe10_io_data_out_15; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_16 = pipe10_io_data_out_16; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_17 = pipe10_io_data_out_17; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_18 = pipe10_io_data_out_18; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_19 = pipe10_io_data_out_19; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_20 = pipe10_io_data_out_20; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_21 = pipe10_io_data_out_21; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_22 = pipe10_io_data_out_22; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_23 = pipe10_io_data_out_23; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_24 = pipe10_io_data_out_24; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_25 = pipe10_io_data_out_25; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_26 = pipe10_io_data_out_26; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_27 = pipe10_io_data_out_27; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_28 = pipe10_io_data_out_28; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_29 = pipe10_io_data_out_29; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_30 = pipe10_io_data_out_30; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_31 = pipe10_io_data_out_31; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_32 = pipe10_io_data_out_32; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_33 = pipe10_io_data_out_33; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_34 = pipe10_io_data_out_34; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_35 = pipe10_io_data_out_35; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_36 = pipe10_io_data_out_36; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_37 = pipe10_io_data_out_37; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_38 = pipe10_io_data_out_38; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_39 = pipe10_io_data_out_39; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_40 = pipe10_io_data_out_40; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_41 = pipe10_io_data_out_41; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_42 = pipe10_io_data_out_42; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_43 = pipe10_io_data_out_43; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_44 = pipe10_io_data_out_44; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_45 = pipe10_io_data_out_45; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_46 = pipe10_io_data_out_46; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_47 = pipe10_io_data_out_47; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_48 = pipe10_io_data_out_48; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_49 = pipe10_io_data_out_49; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_50 = pipe10_io_data_out_50; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_51 = pipe10_io_data_out_51; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_52 = pipe10_io_data_out_52; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_53 = pipe10_io_data_out_53; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_54 = pipe10_io_data_out_54; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_55 = pipe10_io_data_out_55; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_56 = pipe10_io_data_out_56; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_57 = pipe10_io_data_out_57; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_58 = pipe10_io_data_out_58; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_59 = pipe10_io_data_out_59; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_60 = pipe10_io_data_out_60; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_61 = pipe10_io_data_out_61; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_62 = pipe10_io_data_out_62; // @[matcher.scala 380:27]
  assign pipe11_io_data_in_63 = pipe10_io_data_out_63; // @[matcher.scala 380:27]
  assign pipe12_clock = clock;
  assign pipe12_io_pipe_phv_in_data_0 = pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_1 = pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_2 = pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_3 = pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_4 = pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_5 = pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_6 = pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_7 = pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_8 = pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_9 = pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_10 = pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_11 = pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_12 = pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_13 = pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_14 = pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_15 = pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_16 = pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_17 = pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_18 = pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_19 = pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_20 = pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_21 = pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_22 = pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_23 = pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_24 = pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_25 = pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_26 = pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_27 = pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_28 = pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_29 = pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_30 = pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_31 = pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_32 = pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_33 = pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_34 = pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_35 = pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_36 = pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_37 = pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_38 = pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_39 = pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_40 = pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_41 = pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_42 = pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_43 = pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_44 = pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_45 = pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_46 = pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_47 = pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_48 = pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_49 = pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_50 = pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_51 = pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_52 = pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_53 = pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_54 = pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_55 = pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_56 = pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_57 = pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_58 = pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_59 = pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_60 = pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_61 = pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_62 = pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_63 = pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_64 = pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_65 = pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_66 = pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_67 = pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_68 = pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_69 = pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_70 = pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_71 = pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_72 = pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_73 = pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_74 = pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_75 = pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_76 = pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_77 = pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_78 = pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_79 = pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_80 = pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_81 = pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_82 = pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_83 = pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_84 = pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_85 = pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_86 = pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_87 = pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_88 = pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_89 = pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_90 = pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_91 = pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_92 = pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_93 = pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_94 = pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_95 = pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_96 = pipe11_io_pipe_phv_out_data_96; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_97 = pipe11_io_pipe_phv_out_data_97; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_98 = pipe11_io_pipe_phv_out_data_98; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_99 = pipe11_io_pipe_phv_out_data_99; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_100 = pipe11_io_pipe_phv_out_data_100; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_101 = pipe11_io_pipe_phv_out_data_101; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_102 = pipe11_io_pipe_phv_out_data_102; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_103 = pipe11_io_pipe_phv_out_data_103; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_104 = pipe11_io_pipe_phv_out_data_104; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_105 = pipe11_io_pipe_phv_out_data_105; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_106 = pipe11_io_pipe_phv_out_data_106; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_107 = pipe11_io_pipe_phv_out_data_107; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_108 = pipe11_io_pipe_phv_out_data_108; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_109 = pipe11_io_pipe_phv_out_data_109; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_110 = pipe11_io_pipe_phv_out_data_110; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_111 = pipe11_io_pipe_phv_out_data_111; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_112 = pipe11_io_pipe_phv_out_data_112; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_113 = pipe11_io_pipe_phv_out_data_113; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_114 = pipe11_io_pipe_phv_out_data_114; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_115 = pipe11_io_pipe_phv_out_data_115; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_116 = pipe11_io_pipe_phv_out_data_116; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_117 = pipe11_io_pipe_phv_out_data_117; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_118 = pipe11_io_pipe_phv_out_data_118; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_119 = pipe11_io_pipe_phv_out_data_119; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_120 = pipe11_io_pipe_phv_out_data_120; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_121 = pipe11_io_pipe_phv_out_data_121; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_122 = pipe11_io_pipe_phv_out_data_122; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_123 = pipe11_io_pipe_phv_out_data_123; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_124 = pipe11_io_pipe_phv_out_data_124; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_125 = pipe11_io_pipe_phv_out_data_125; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_126 = pipe11_io_pipe_phv_out_data_126; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_127 = pipe11_io_pipe_phv_out_data_127; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_128 = pipe11_io_pipe_phv_out_data_128; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_129 = pipe11_io_pipe_phv_out_data_129; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_130 = pipe11_io_pipe_phv_out_data_130; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_131 = pipe11_io_pipe_phv_out_data_131; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_132 = pipe11_io_pipe_phv_out_data_132; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_133 = pipe11_io_pipe_phv_out_data_133; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_134 = pipe11_io_pipe_phv_out_data_134; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_135 = pipe11_io_pipe_phv_out_data_135; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_136 = pipe11_io_pipe_phv_out_data_136; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_137 = pipe11_io_pipe_phv_out_data_137; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_138 = pipe11_io_pipe_phv_out_data_138; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_139 = pipe11_io_pipe_phv_out_data_139; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_140 = pipe11_io_pipe_phv_out_data_140; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_141 = pipe11_io_pipe_phv_out_data_141; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_142 = pipe11_io_pipe_phv_out_data_142; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_143 = pipe11_io_pipe_phv_out_data_143; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_144 = pipe11_io_pipe_phv_out_data_144; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_145 = pipe11_io_pipe_phv_out_data_145; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_146 = pipe11_io_pipe_phv_out_data_146; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_147 = pipe11_io_pipe_phv_out_data_147; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_148 = pipe11_io_pipe_phv_out_data_148; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_149 = pipe11_io_pipe_phv_out_data_149; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_150 = pipe11_io_pipe_phv_out_data_150; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_151 = pipe11_io_pipe_phv_out_data_151; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_152 = pipe11_io_pipe_phv_out_data_152; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_153 = pipe11_io_pipe_phv_out_data_153; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_154 = pipe11_io_pipe_phv_out_data_154; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_155 = pipe11_io_pipe_phv_out_data_155; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_156 = pipe11_io_pipe_phv_out_data_156; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_157 = pipe11_io_pipe_phv_out_data_157; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_158 = pipe11_io_pipe_phv_out_data_158; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_159 = pipe11_io_pipe_phv_out_data_159; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_160 = pipe11_io_pipe_phv_out_data_160; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_161 = pipe11_io_pipe_phv_out_data_161; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_162 = pipe11_io_pipe_phv_out_data_162; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_163 = pipe11_io_pipe_phv_out_data_163; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_164 = pipe11_io_pipe_phv_out_data_164; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_165 = pipe11_io_pipe_phv_out_data_165; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_166 = pipe11_io_pipe_phv_out_data_166; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_167 = pipe11_io_pipe_phv_out_data_167; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_168 = pipe11_io_pipe_phv_out_data_168; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_169 = pipe11_io_pipe_phv_out_data_169; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_170 = pipe11_io_pipe_phv_out_data_170; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_171 = pipe11_io_pipe_phv_out_data_171; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_172 = pipe11_io_pipe_phv_out_data_172; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_173 = pipe11_io_pipe_phv_out_data_173; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_174 = pipe11_io_pipe_phv_out_data_174; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_175 = pipe11_io_pipe_phv_out_data_175; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_176 = pipe11_io_pipe_phv_out_data_176; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_177 = pipe11_io_pipe_phv_out_data_177; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_178 = pipe11_io_pipe_phv_out_data_178; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_179 = pipe11_io_pipe_phv_out_data_179; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_180 = pipe11_io_pipe_phv_out_data_180; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_181 = pipe11_io_pipe_phv_out_data_181; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_182 = pipe11_io_pipe_phv_out_data_182; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_183 = pipe11_io_pipe_phv_out_data_183; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_184 = pipe11_io_pipe_phv_out_data_184; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_185 = pipe11_io_pipe_phv_out_data_185; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_186 = pipe11_io_pipe_phv_out_data_186; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_187 = pipe11_io_pipe_phv_out_data_187; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_188 = pipe11_io_pipe_phv_out_data_188; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_189 = pipe11_io_pipe_phv_out_data_189; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_190 = pipe11_io_pipe_phv_out_data_190; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_191 = pipe11_io_pipe_phv_out_data_191; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_192 = pipe11_io_pipe_phv_out_data_192; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_193 = pipe11_io_pipe_phv_out_data_193; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_194 = pipe11_io_pipe_phv_out_data_194; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_195 = pipe11_io_pipe_phv_out_data_195; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_196 = pipe11_io_pipe_phv_out_data_196; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_197 = pipe11_io_pipe_phv_out_data_197; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_198 = pipe11_io_pipe_phv_out_data_198; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_199 = pipe11_io_pipe_phv_out_data_199; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_200 = pipe11_io_pipe_phv_out_data_200; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_201 = pipe11_io_pipe_phv_out_data_201; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_202 = pipe11_io_pipe_phv_out_data_202; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_203 = pipe11_io_pipe_phv_out_data_203; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_204 = pipe11_io_pipe_phv_out_data_204; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_205 = pipe11_io_pipe_phv_out_data_205; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_206 = pipe11_io_pipe_phv_out_data_206; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_207 = pipe11_io_pipe_phv_out_data_207; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_208 = pipe11_io_pipe_phv_out_data_208; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_209 = pipe11_io_pipe_phv_out_data_209; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_210 = pipe11_io_pipe_phv_out_data_210; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_211 = pipe11_io_pipe_phv_out_data_211; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_212 = pipe11_io_pipe_phv_out_data_212; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_213 = pipe11_io_pipe_phv_out_data_213; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_214 = pipe11_io_pipe_phv_out_data_214; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_215 = pipe11_io_pipe_phv_out_data_215; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_216 = pipe11_io_pipe_phv_out_data_216; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_217 = pipe11_io_pipe_phv_out_data_217; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_218 = pipe11_io_pipe_phv_out_data_218; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_219 = pipe11_io_pipe_phv_out_data_219; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_220 = pipe11_io_pipe_phv_out_data_220; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_221 = pipe11_io_pipe_phv_out_data_221; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_222 = pipe11_io_pipe_phv_out_data_222; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_223 = pipe11_io_pipe_phv_out_data_223; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_224 = pipe11_io_pipe_phv_out_data_224; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_225 = pipe11_io_pipe_phv_out_data_225; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_226 = pipe11_io_pipe_phv_out_data_226; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_227 = pipe11_io_pipe_phv_out_data_227; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_228 = pipe11_io_pipe_phv_out_data_228; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_229 = pipe11_io_pipe_phv_out_data_229; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_230 = pipe11_io_pipe_phv_out_data_230; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_231 = pipe11_io_pipe_phv_out_data_231; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_232 = pipe11_io_pipe_phv_out_data_232; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_233 = pipe11_io_pipe_phv_out_data_233; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_234 = pipe11_io_pipe_phv_out_data_234; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_235 = pipe11_io_pipe_phv_out_data_235; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_236 = pipe11_io_pipe_phv_out_data_236; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_237 = pipe11_io_pipe_phv_out_data_237; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_238 = pipe11_io_pipe_phv_out_data_238; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_239 = pipe11_io_pipe_phv_out_data_239; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_240 = pipe11_io_pipe_phv_out_data_240; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_241 = pipe11_io_pipe_phv_out_data_241; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_242 = pipe11_io_pipe_phv_out_data_242; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_243 = pipe11_io_pipe_phv_out_data_243; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_244 = pipe11_io_pipe_phv_out_data_244; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_245 = pipe11_io_pipe_phv_out_data_245; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_246 = pipe11_io_pipe_phv_out_data_246; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_247 = pipe11_io_pipe_phv_out_data_247; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_248 = pipe11_io_pipe_phv_out_data_248; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_249 = pipe11_io_pipe_phv_out_data_249; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_250 = pipe11_io_pipe_phv_out_data_250; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_251 = pipe11_io_pipe_phv_out_data_251; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_252 = pipe11_io_pipe_phv_out_data_252; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_253 = pipe11_io_pipe_phv_out_data_253; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_254 = pipe11_io_pipe_phv_out_data_254; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_255 = pipe11_io_pipe_phv_out_data_255; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_0 = pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_1 = pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_2 = pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_3 = pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_4 = pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_5 = pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_6 = pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_7 = pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_8 = pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_9 = pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_10 = pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_11 = pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_12 = pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_13 = pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_14 = pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_15 = pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_current_state = pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_current_offset = pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_transition_field = pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_next_processor_id = pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_next_config_id = pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_is_valid_processor = pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 383:27]
  assign pipe12_io_key_config_0_key_length = key_config_0_key_length; // @[matcher.scala 386:27]
  assign pipe12_io_key_config_1_key_length = key_config_1_key_length; // @[matcher.scala 386:27]
  assign pipe12_io_key_in = pipe11_io_key_out; // @[matcher.scala 384:27]
  assign pipe12_io_data_in = pipe11_io_data_out; // @[matcher.scala 385:27]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_0_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_header_id <= io_mod_key_mod_header_id; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_internal_offset <= io_mod_key_mod_internal_offset; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 21:40]
        key_config_1_key_length <= io_mod_key_mod_key_length; // @[matcher.scala 21:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_0 <= io_mod_table_mod_sram_id_table_0; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_1 <= io_mod_table_mod_sram_id_table_1; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_2 <= io_mod_table_mod_sram_id_table_2; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_3 <= io_mod_table_mod_sram_id_table_3; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_4 <= io_mod_table_mod_sram_id_table_4; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_5 <= io_mod_table_mod_sram_id_table_5; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_6 <= io_mod_table_mod_sram_id_table_6; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_7 <= io_mod_table_mod_sram_id_table_7; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_8 <= io_mod_table_mod_sram_id_table_8; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_9 <= io_mod_table_mod_sram_id_table_9; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_10 <= io_mod_table_mod_sram_id_table_10; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_11 <= io_mod_table_mod_sram_id_table_11; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_12 <= io_mod_table_mod_sram_id_table_12; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_13 <= io_mod_table_mod_sram_id_table_13; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_14 <= io_mod_table_mod_sram_id_table_14; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_15 <= io_mod_table_mod_sram_id_table_15; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_16 <= io_mod_table_mod_sram_id_table_16; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_17 <= io_mod_table_mod_sram_id_table_17; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_18 <= io_mod_table_mod_sram_id_table_18; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_19 <= io_mod_table_mod_sram_id_table_19; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_20 <= io_mod_table_mod_sram_id_table_20; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_21 <= io_mod_table_mod_sram_id_table_21; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_22 <= io_mod_table_mod_sram_id_table_22; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_23 <= io_mod_table_mod_sram_id_table_23; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_24 <= io_mod_table_mod_sram_id_table_24; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_25 <= io_mod_table_mod_sram_id_table_25; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_26 <= io_mod_table_mod_sram_id_table_26; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_27 <= io_mod_table_mod_sram_id_table_27; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_28 <= io_mod_table_mod_sram_id_table_28; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_29 <= io_mod_table_mod_sram_id_table_29; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_30 <= io_mod_table_mod_sram_id_table_30; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_31 <= io_mod_table_mod_sram_id_table_31; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_32 <= io_mod_table_mod_sram_id_table_32; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_33 <= io_mod_table_mod_sram_id_table_33; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_34 <= io_mod_table_mod_sram_id_table_34; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_35 <= io_mod_table_mod_sram_id_table_35; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_36 <= io_mod_table_mod_sram_id_table_36; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_37 <= io_mod_table_mod_sram_id_table_37; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_38 <= io_mod_table_mod_sram_id_table_38; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_39 <= io_mod_table_mod_sram_id_table_39; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_40 <= io_mod_table_mod_sram_id_table_40; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_41 <= io_mod_table_mod_sram_id_table_41; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_42 <= io_mod_table_mod_sram_id_table_42; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_43 <= io_mod_table_mod_sram_id_table_43; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_44 <= io_mod_table_mod_sram_id_table_44; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_45 <= io_mod_table_mod_sram_id_table_45; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_46 <= io_mod_table_mod_sram_id_table_46; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_47 <= io_mod_table_mod_sram_id_table_47; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_48 <= io_mod_table_mod_sram_id_table_48; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_49 <= io_mod_table_mod_sram_id_table_49; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_50 <= io_mod_table_mod_sram_id_table_50; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_51 <= io_mod_table_mod_sram_id_table_51; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_52 <= io_mod_table_mod_sram_id_table_52; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_53 <= io_mod_table_mod_sram_id_table_53; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_54 <= io_mod_table_mod_sram_id_table_54; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_55 <= io_mod_table_mod_sram_id_table_55; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_56 <= io_mod_table_mod_sram_id_table_56; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_57 <= io_mod_table_mod_sram_id_table_57; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_58 <= io_mod_table_mod_sram_id_table_58; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_59 <= io_mod_table_mod_sram_id_table_59; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_60 <= io_mod_table_mod_sram_id_table_60; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_61 <= io_mod_table_mod_sram_id_table_61; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_62 <= io_mod_table_mod_sram_id_table_62; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_sram_id_table_63 <= io_mod_table_mod_sram_id_table_63; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (~io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_0_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_0 <= io_mod_table_mod_sram_id_table_0; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_1 <= io_mod_table_mod_sram_id_table_1; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_2 <= io_mod_table_mod_sram_id_table_2; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_3 <= io_mod_table_mod_sram_id_table_3; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_4 <= io_mod_table_mod_sram_id_table_4; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_5 <= io_mod_table_mod_sram_id_table_5; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_6 <= io_mod_table_mod_sram_id_table_6; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_7 <= io_mod_table_mod_sram_id_table_7; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_8 <= io_mod_table_mod_sram_id_table_8; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_9 <= io_mod_table_mod_sram_id_table_9; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_10 <= io_mod_table_mod_sram_id_table_10; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_11 <= io_mod_table_mod_sram_id_table_11; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_12 <= io_mod_table_mod_sram_id_table_12; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_13 <= io_mod_table_mod_sram_id_table_13; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_14 <= io_mod_table_mod_sram_id_table_14; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_15 <= io_mod_table_mod_sram_id_table_15; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_16 <= io_mod_table_mod_sram_id_table_16; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_17 <= io_mod_table_mod_sram_id_table_17; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_18 <= io_mod_table_mod_sram_id_table_18; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_19 <= io_mod_table_mod_sram_id_table_19; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_20 <= io_mod_table_mod_sram_id_table_20; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_21 <= io_mod_table_mod_sram_id_table_21; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_22 <= io_mod_table_mod_sram_id_table_22; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_23 <= io_mod_table_mod_sram_id_table_23; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_24 <= io_mod_table_mod_sram_id_table_24; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_25 <= io_mod_table_mod_sram_id_table_25; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_26 <= io_mod_table_mod_sram_id_table_26; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_27 <= io_mod_table_mod_sram_id_table_27; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_28 <= io_mod_table_mod_sram_id_table_28; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_29 <= io_mod_table_mod_sram_id_table_29; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_30 <= io_mod_table_mod_sram_id_table_30; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_31 <= io_mod_table_mod_sram_id_table_31; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_32 <= io_mod_table_mod_sram_id_table_32; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_33 <= io_mod_table_mod_sram_id_table_33; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_34 <= io_mod_table_mod_sram_id_table_34; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_35 <= io_mod_table_mod_sram_id_table_35; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_36 <= io_mod_table_mod_sram_id_table_36; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_37 <= io_mod_table_mod_sram_id_table_37; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_38 <= io_mod_table_mod_sram_id_table_38; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_39 <= io_mod_table_mod_sram_id_table_39; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_40 <= io_mod_table_mod_sram_id_table_40; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_41 <= io_mod_table_mod_sram_id_table_41; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_42 <= io_mod_table_mod_sram_id_table_42; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_43 <= io_mod_table_mod_sram_id_table_43; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_44 <= io_mod_table_mod_sram_id_table_44; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_45 <= io_mod_table_mod_sram_id_table_45; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_46 <= io_mod_table_mod_sram_id_table_46; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_47 <= io_mod_table_mod_sram_id_table_47; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_48 <= io_mod_table_mod_sram_id_table_48; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_49 <= io_mod_table_mod_sram_id_table_49; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_50 <= io_mod_table_mod_sram_id_table_50; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_51 <= io_mod_table_mod_sram_id_table_51; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_52 <= io_mod_table_mod_sram_id_table_52; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_53 <= io_mod_table_mod_sram_id_table_53; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_54 <= io_mod_table_mod_sram_id_table_54; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_55 <= io_mod_table_mod_sram_id_table_55; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_56 <= io_mod_table_mod_sram_id_table_56; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_57 <= io_mod_table_mod_sram_id_table_57; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_58 <= io_mod_table_mod_sram_id_table_58; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_59 <= io_mod_table_mod_sram_id_table_59; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_60 <= io_mod_table_mod_sram_id_table_60; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_61 <= io_mod_table_mod_sram_id_table_61; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_62 <= io_mod_table_mod_sram_id_table_62; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_sram_id_table_63 <= io_mod_table_mod_sram_id_table_63; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_width <= io_mod_table_mod_table_width; // @[matcher.scala 22:40]
      end
    end
    if (io_mod_en) begin // @[matcher.scala 20:22]
      if (io_mod_config_id) begin // @[matcher.scala 22:40]
        table_config_1_table_depth <= io_mod_table_mod_table_depth; // @[matcher.scala 22:40]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  key_config_0_header_id = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  key_config_0_internal_offset = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  key_config_0_key_length = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  key_config_1_header_id = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  key_config_1_internal_offset = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  key_config_1_key_length = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  table_config_0_sram_id_table_0 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  table_config_0_sram_id_table_1 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  table_config_0_sram_id_table_2 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  table_config_0_sram_id_table_3 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  table_config_0_sram_id_table_4 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  table_config_0_sram_id_table_5 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  table_config_0_sram_id_table_6 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  table_config_0_sram_id_table_7 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  table_config_0_sram_id_table_8 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  table_config_0_sram_id_table_9 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  table_config_0_sram_id_table_10 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  table_config_0_sram_id_table_11 = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  table_config_0_sram_id_table_12 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  table_config_0_sram_id_table_13 = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  table_config_0_sram_id_table_14 = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  table_config_0_sram_id_table_15 = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  table_config_0_sram_id_table_16 = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  table_config_0_sram_id_table_17 = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  table_config_0_sram_id_table_18 = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  table_config_0_sram_id_table_19 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  table_config_0_sram_id_table_20 = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  table_config_0_sram_id_table_21 = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  table_config_0_sram_id_table_22 = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  table_config_0_sram_id_table_23 = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  table_config_0_sram_id_table_24 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  table_config_0_sram_id_table_25 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  table_config_0_sram_id_table_26 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  table_config_0_sram_id_table_27 = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  table_config_0_sram_id_table_28 = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  table_config_0_sram_id_table_29 = _RAND_35[5:0];
  _RAND_36 = {1{`RANDOM}};
  table_config_0_sram_id_table_30 = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  table_config_0_sram_id_table_31 = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  table_config_0_sram_id_table_32 = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  table_config_0_sram_id_table_33 = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  table_config_0_sram_id_table_34 = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  table_config_0_sram_id_table_35 = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  table_config_0_sram_id_table_36 = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  table_config_0_sram_id_table_37 = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  table_config_0_sram_id_table_38 = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  table_config_0_sram_id_table_39 = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  table_config_0_sram_id_table_40 = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  table_config_0_sram_id_table_41 = _RAND_47[5:0];
  _RAND_48 = {1{`RANDOM}};
  table_config_0_sram_id_table_42 = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  table_config_0_sram_id_table_43 = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  table_config_0_sram_id_table_44 = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  table_config_0_sram_id_table_45 = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
  table_config_0_sram_id_table_46 = _RAND_52[5:0];
  _RAND_53 = {1{`RANDOM}};
  table_config_0_sram_id_table_47 = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  table_config_0_sram_id_table_48 = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  table_config_0_sram_id_table_49 = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  table_config_0_sram_id_table_50 = _RAND_56[5:0];
  _RAND_57 = {1{`RANDOM}};
  table_config_0_sram_id_table_51 = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  table_config_0_sram_id_table_52 = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  table_config_0_sram_id_table_53 = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  table_config_0_sram_id_table_54 = _RAND_60[5:0];
  _RAND_61 = {1{`RANDOM}};
  table_config_0_sram_id_table_55 = _RAND_61[5:0];
  _RAND_62 = {1{`RANDOM}};
  table_config_0_sram_id_table_56 = _RAND_62[5:0];
  _RAND_63 = {1{`RANDOM}};
  table_config_0_sram_id_table_57 = _RAND_63[5:0];
  _RAND_64 = {1{`RANDOM}};
  table_config_0_sram_id_table_58 = _RAND_64[5:0];
  _RAND_65 = {1{`RANDOM}};
  table_config_0_sram_id_table_59 = _RAND_65[5:0];
  _RAND_66 = {1{`RANDOM}};
  table_config_0_sram_id_table_60 = _RAND_66[5:0];
  _RAND_67 = {1{`RANDOM}};
  table_config_0_sram_id_table_61 = _RAND_67[5:0];
  _RAND_68 = {1{`RANDOM}};
  table_config_0_sram_id_table_62 = _RAND_68[5:0];
  _RAND_69 = {1{`RANDOM}};
  table_config_0_sram_id_table_63 = _RAND_69[5:0];
  _RAND_70 = {1{`RANDOM}};
  table_config_0_table_width = _RAND_70[6:0];
  _RAND_71 = {1{`RANDOM}};
  table_config_0_table_depth = _RAND_71[6:0];
  _RAND_72 = {1{`RANDOM}};
  table_config_1_sram_id_table_0 = _RAND_72[5:0];
  _RAND_73 = {1{`RANDOM}};
  table_config_1_sram_id_table_1 = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  table_config_1_sram_id_table_2 = _RAND_74[5:0];
  _RAND_75 = {1{`RANDOM}};
  table_config_1_sram_id_table_3 = _RAND_75[5:0];
  _RAND_76 = {1{`RANDOM}};
  table_config_1_sram_id_table_4 = _RAND_76[5:0];
  _RAND_77 = {1{`RANDOM}};
  table_config_1_sram_id_table_5 = _RAND_77[5:0];
  _RAND_78 = {1{`RANDOM}};
  table_config_1_sram_id_table_6 = _RAND_78[5:0];
  _RAND_79 = {1{`RANDOM}};
  table_config_1_sram_id_table_7 = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  table_config_1_sram_id_table_8 = _RAND_80[5:0];
  _RAND_81 = {1{`RANDOM}};
  table_config_1_sram_id_table_9 = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  table_config_1_sram_id_table_10 = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  table_config_1_sram_id_table_11 = _RAND_83[5:0];
  _RAND_84 = {1{`RANDOM}};
  table_config_1_sram_id_table_12 = _RAND_84[5:0];
  _RAND_85 = {1{`RANDOM}};
  table_config_1_sram_id_table_13 = _RAND_85[5:0];
  _RAND_86 = {1{`RANDOM}};
  table_config_1_sram_id_table_14 = _RAND_86[5:0];
  _RAND_87 = {1{`RANDOM}};
  table_config_1_sram_id_table_15 = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  table_config_1_sram_id_table_16 = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  table_config_1_sram_id_table_17 = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  table_config_1_sram_id_table_18 = _RAND_90[5:0];
  _RAND_91 = {1{`RANDOM}};
  table_config_1_sram_id_table_19 = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  table_config_1_sram_id_table_20 = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  table_config_1_sram_id_table_21 = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  table_config_1_sram_id_table_22 = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  table_config_1_sram_id_table_23 = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  table_config_1_sram_id_table_24 = _RAND_96[5:0];
  _RAND_97 = {1{`RANDOM}};
  table_config_1_sram_id_table_25 = _RAND_97[5:0];
  _RAND_98 = {1{`RANDOM}};
  table_config_1_sram_id_table_26 = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  table_config_1_sram_id_table_27 = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  table_config_1_sram_id_table_28 = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  table_config_1_sram_id_table_29 = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  table_config_1_sram_id_table_30 = _RAND_102[5:0];
  _RAND_103 = {1{`RANDOM}};
  table_config_1_sram_id_table_31 = _RAND_103[5:0];
  _RAND_104 = {1{`RANDOM}};
  table_config_1_sram_id_table_32 = _RAND_104[5:0];
  _RAND_105 = {1{`RANDOM}};
  table_config_1_sram_id_table_33 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  table_config_1_sram_id_table_34 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  table_config_1_sram_id_table_35 = _RAND_107[5:0];
  _RAND_108 = {1{`RANDOM}};
  table_config_1_sram_id_table_36 = _RAND_108[5:0];
  _RAND_109 = {1{`RANDOM}};
  table_config_1_sram_id_table_37 = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  table_config_1_sram_id_table_38 = _RAND_110[5:0];
  _RAND_111 = {1{`RANDOM}};
  table_config_1_sram_id_table_39 = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  table_config_1_sram_id_table_40 = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  table_config_1_sram_id_table_41 = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  table_config_1_sram_id_table_42 = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  table_config_1_sram_id_table_43 = _RAND_115[5:0];
  _RAND_116 = {1{`RANDOM}};
  table_config_1_sram_id_table_44 = _RAND_116[5:0];
  _RAND_117 = {1{`RANDOM}};
  table_config_1_sram_id_table_45 = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  table_config_1_sram_id_table_46 = _RAND_118[5:0];
  _RAND_119 = {1{`RANDOM}};
  table_config_1_sram_id_table_47 = _RAND_119[5:0];
  _RAND_120 = {1{`RANDOM}};
  table_config_1_sram_id_table_48 = _RAND_120[5:0];
  _RAND_121 = {1{`RANDOM}};
  table_config_1_sram_id_table_49 = _RAND_121[5:0];
  _RAND_122 = {1{`RANDOM}};
  table_config_1_sram_id_table_50 = _RAND_122[5:0];
  _RAND_123 = {1{`RANDOM}};
  table_config_1_sram_id_table_51 = _RAND_123[5:0];
  _RAND_124 = {1{`RANDOM}};
  table_config_1_sram_id_table_52 = _RAND_124[5:0];
  _RAND_125 = {1{`RANDOM}};
  table_config_1_sram_id_table_53 = _RAND_125[5:0];
  _RAND_126 = {1{`RANDOM}};
  table_config_1_sram_id_table_54 = _RAND_126[5:0];
  _RAND_127 = {1{`RANDOM}};
  table_config_1_sram_id_table_55 = _RAND_127[5:0];
  _RAND_128 = {1{`RANDOM}};
  table_config_1_sram_id_table_56 = _RAND_128[5:0];
  _RAND_129 = {1{`RANDOM}};
  table_config_1_sram_id_table_57 = _RAND_129[5:0];
  _RAND_130 = {1{`RANDOM}};
  table_config_1_sram_id_table_58 = _RAND_130[5:0];
  _RAND_131 = {1{`RANDOM}};
  table_config_1_sram_id_table_59 = _RAND_131[5:0];
  _RAND_132 = {1{`RANDOM}};
  table_config_1_sram_id_table_60 = _RAND_132[5:0];
  _RAND_133 = {1{`RANDOM}};
  table_config_1_sram_id_table_61 = _RAND_133[5:0];
  _RAND_134 = {1{`RANDOM}};
  table_config_1_sram_id_table_62 = _RAND_134[5:0];
  _RAND_135 = {1{`RANDOM}};
  table_config_1_sram_id_table_63 = _RAND_135[5:0];
  _RAND_136 = {1{`RANDOM}};
  table_config_1_table_width = _RAND_136[6:0];
  _RAND_137 = {1{`RANDOM}};
  table_config_1_table_depth = _RAND_137[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
