module PISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  input         io_mod_par_mod_en,
  input         io_mod_par_mod_last_mau_id_mod,
  input  [3:0]  io_mod_par_mod_last_mau_id,
  input  [2:0]  io_mod_par_mod_cs,
  input         io_mod_par_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_par_mod_module_mod_state_id,
  input         io_mod_par_mod_module_mod_sram_w_cs,
  input         io_mod_par_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_par_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_par_mod_module_mod_sram_w_data,
  input         io_mod_proc_mod_0_mat_mod_en,
  input         io_mod_proc_mod_0_mat_mod_config_id,
  input         io_mod_proc_mod_0_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_0_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_0_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_0_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_0_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_0_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_0_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_0_mat_mod_w_data,
  input         io_mod_proc_mod_0_exe_mod_en_0,
  input         io_mod_proc_mod_0_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_0_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_0_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_0_exe_mod_data_1,
  input         io_mod_proc_mod_1_mat_mod_en,
  input         io_mod_proc_mod_1_mat_mod_config_id,
  input         io_mod_proc_mod_1_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_1_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_1_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_1_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_1_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_1_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_1_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_1_mat_mod_w_data,
  input         io_mod_proc_mod_1_exe_mod_en_0,
  input         io_mod_proc_mod_1_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_1_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_1_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_1_exe_mod_data_1,
  input         io_mod_proc_mod_2_mat_mod_en,
  input         io_mod_proc_mod_2_mat_mod_config_id,
  input         io_mod_proc_mod_2_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_2_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_2_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_2_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_2_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_2_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_2_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_2_mat_mod_w_data,
  input         io_mod_proc_mod_2_exe_mod_en_0,
  input         io_mod_proc_mod_2_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_2_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_2_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_2_exe_mod_data_1,
  input         io_mod_proc_mod_3_mat_mod_en,
  input         io_mod_proc_mod_3_mat_mod_config_id,
  input         io_mod_proc_mod_3_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_3_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_3_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_3_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_3_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_3_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_3_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_3_mat_mod_w_data,
  input         io_mod_proc_mod_3_exe_mod_en_0,
  input         io_mod_proc_mod_3_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_3_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_3_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_3_exe_mod_data_1,
  input         io_mod_proc_mod_4_mat_mod_en,
  input         io_mod_proc_mod_4_mat_mod_config_id,
  input         io_mod_proc_mod_4_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_4_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_4_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_4_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_4_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_4_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_4_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_4_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_4_mat_mod_w_data,
  input         io_mod_proc_mod_4_exe_mod_en_0,
  input         io_mod_proc_mod_4_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_4_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_4_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_4_exe_mod_data_1,
  input         io_mod_proc_mod_5_mat_mod_en,
  input         io_mod_proc_mod_5_mat_mod_config_id,
  input         io_mod_proc_mod_5_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_5_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_5_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_5_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_5_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_5_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_5_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_5_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_5_mat_mod_w_data,
  input         io_mod_proc_mod_5_exe_mod_en_0,
  input         io_mod_proc_mod_5_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_5_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_5_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_5_exe_mod_data_1,
  input         io_mod_proc_mod_6_mat_mod_en,
  input         io_mod_proc_mod_6_mat_mod_config_id,
  input         io_mod_proc_mod_6_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_6_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_6_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_6_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_6_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_6_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_6_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_6_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_6_mat_mod_w_data,
  input         io_mod_proc_mod_6_exe_mod_en_0,
  input         io_mod_proc_mod_6_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_6_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_6_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_6_exe_mod_data_1,
  input         io_mod_proc_mod_7_mat_mod_en,
  input         io_mod_proc_mod_7_mat_mod_config_id,
  input         io_mod_proc_mod_7_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_7_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_7_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_7_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_7_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_7_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_7_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_7_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_7_mat_mod_w_data,
  input         io_mod_proc_mod_7_exe_mod_en_0,
  input         io_mod_proc_mod_7_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_7_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_7_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_7_exe_mod_data_1,
  input         io_mod_proc_mod_8_mat_mod_en,
  input         io_mod_proc_mod_8_mat_mod_config_id,
  input         io_mod_proc_mod_8_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_8_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_8_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_8_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_8_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_8_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_8_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_8_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_8_mat_mod_w_data,
  input         io_mod_proc_mod_8_exe_mod_en_0,
  input         io_mod_proc_mod_8_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_8_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_8_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_8_exe_mod_data_1,
  input         io_mod_proc_mod_9_mat_mod_en,
  input         io_mod_proc_mod_9_mat_mod_config_id,
  input         io_mod_proc_mod_9_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_9_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_9_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_9_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_9_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_9_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_9_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_9_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_9_mat_mod_w_data,
  input         io_mod_proc_mod_9_exe_mod_en_0,
  input         io_mod_proc_mod_9_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_9_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_9_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_9_exe_mod_data_1,
  input         io_mod_proc_mod_10_mat_mod_en,
  input         io_mod_proc_mod_10_mat_mod_config_id,
  input         io_mod_proc_mod_10_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_10_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_10_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_10_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_10_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_10_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_10_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_10_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_10_mat_mod_w_data,
  input         io_mod_proc_mod_10_exe_mod_en_0,
  input         io_mod_proc_mod_10_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_10_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_10_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_10_exe_mod_data_1,
  input         io_mod_proc_mod_11_mat_mod_en,
  input         io_mod_proc_mod_11_mat_mod_config_id,
  input         io_mod_proc_mod_11_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_11_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_11_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_11_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_11_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_11_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_11_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_11_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_11_mat_mod_w_data,
  input         io_mod_proc_mod_11_exe_mod_en_0,
  input         io_mod_proc_mod_11_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_11_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_11_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_11_exe_mod_data_1,
  input         io_mod_proc_mod_12_mat_mod_en,
  input         io_mod_proc_mod_12_mat_mod_config_id,
  input         io_mod_proc_mod_12_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_12_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_12_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_12_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_12_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_12_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_12_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_12_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_12_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_12_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_12_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_12_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_12_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_12_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_12_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_12_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_12_mat_mod_w_data,
  input         io_mod_proc_mod_12_exe_mod_en_0,
  input         io_mod_proc_mod_12_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_12_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_12_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_12_exe_mod_data_1,
  input         io_mod_proc_mod_13_mat_mod_en,
  input         io_mod_proc_mod_13_mat_mod_config_id,
  input         io_mod_proc_mod_13_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_13_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_13_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_13_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_13_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_13_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_13_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_13_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_13_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_13_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_13_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_13_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_13_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_13_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_13_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_13_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_13_mat_mod_w_data,
  input         io_mod_proc_mod_13_exe_mod_en_0,
  input         io_mod_proc_mod_13_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_13_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_13_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_13_exe_mod_data_1,
  input         io_mod_proc_mod_14_mat_mod_en,
  input         io_mod_proc_mod_14_mat_mod_config_id,
  input         io_mod_proc_mod_14_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_14_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_14_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_14_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_14_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_14_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_14_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_14_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_14_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_14_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_14_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_14_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_14_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_14_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_14_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_14_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_14_mat_mod_w_data,
  input         io_mod_proc_mod_14_exe_mod_en_0,
  input         io_mod_proc_mod_14_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_14_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_14_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_14_exe_mod_data_1,
  input         io_mod_proc_mod_15_mat_mod_en,
  input         io_mod_proc_mod_15_mat_mod_config_id,
  input         io_mod_proc_mod_15_mat_mod_key_mod_en,
  input  [2:0]  io_mod_proc_mod_15_mat_mod_key_mod_group_index,
  input  [1:0]  io_mod_proc_mod_15_mat_mod_key_mod_group_config,
  input         io_mod_proc_mod_15_mat_mod_key_mod_group_mask_0,
  input         io_mod_proc_mod_15_mat_mod_key_mod_group_mask_1,
  input         io_mod_proc_mod_15_mat_mod_key_mod_group_mask_2,
  input         io_mod_proc_mod_15_mat_mod_key_mod_group_mask_3,
  input  [6:0]  io_mod_proc_mod_15_mat_mod_key_mod_group_id_0,
  input  [6:0]  io_mod_proc_mod_15_mat_mod_key_mod_group_id_1,
  input  [6:0]  io_mod_proc_mod_15_mat_mod_key_mod_group_id_2,
  input  [6:0]  io_mod_proc_mod_15_mat_mod_key_mod_group_id_3,
  input  [4:0]  io_mod_proc_mod_15_mat_mod_table_mod_table_depth,
  input  [4:0]  io_mod_proc_mod_15_mat_mod_table_mod_table_width,
  input         io_mod_proc_mod_15_mat_mod_w_en,
  input  [3:0]  io_mod_proc_mod_15_mat_mod_w_sram_id,
  input  [7:0]  io_mod_proc_mod_15_mat_mod_w_addr,
  input  [63:0] io_mod_proc_mod_15_mat_mod_w_data,
  input         io_mod_proc_mod_15_exe_mod_en_0,
  input         io_mod_proc_mod_15_exe_mod_en_1,
  input  [7:0]  io_mod_proc_mod_15_exe_mod_addr,
  input  [63:0] io_mod_proc_mod_15_exe_mod_data_0,
  input  [63:0] io_mod_proc_mod_15_exe_mod_data_1
);
  wire  init_clock; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_0; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_1; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_2; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_3; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_4; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_5; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_6; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_7; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_8; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_9; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_10; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_11; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_12; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_13; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_14; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_15; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_16; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_17; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_18; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_19; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_20; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_21; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_22; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_23; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_24; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_25; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_26; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_27; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_28; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_29; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_30; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_31; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_32; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_33; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_34; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_35; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_36; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_37; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_38; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_39; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_40; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_41; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_42; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_43; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_44; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_45; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_46; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_47; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_48; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_49; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_50; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_51; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_52; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_53; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_54; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_55; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_56; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_57; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_58; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_59; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_60; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_61; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_62; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_63; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_64; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_65; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_66; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_67; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_68; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_69; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_70; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_71; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_72; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_73; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_74; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_75; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_76; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_77; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_78; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_79; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_80; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_81; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_82; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_83; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_84; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_85; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_86; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_87; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_88; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_89; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_90; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_91; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_92; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_93; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_94; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_95; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_96; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_97; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_98; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_99; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_100; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_101; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_102; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_103; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_104; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_105; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_106; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_107; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_108; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_109; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_110; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_111; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_112; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_113; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_114; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_115; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_116; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_117; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_118; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_119; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_120; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_121; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_122; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_123; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_124; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_125; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_126; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_in_data_127; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_0; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_1; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_2; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_3; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_4; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_5; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_6; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_7; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_8; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_9; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_10; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_11; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_12; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_13; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_14; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_15; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_16; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_17; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_18; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_19; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_20; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_21; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_22; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_23; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_24; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_25; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_26; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_27; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_28; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_29; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_30; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_31; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_32; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_33; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_34; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_35; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_36; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_37; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_38; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_39; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_40; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_41; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_42; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_43; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_44; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_45; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_46; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_47; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_48; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_49; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_50; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_51; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_52; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_53; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_54; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_55; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_56; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_57; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_58; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_59; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_60; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_61; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_62; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_63; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_64; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_65; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_66; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_67; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_68; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_69; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_70; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_71; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_72; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_73; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_74; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_75; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_76; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_77; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_78; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_79; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_80; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_81; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_82; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_83; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_84; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_85; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_86; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_87; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_88; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_89; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_90; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_91; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_92; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_93; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_94; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_95; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_96; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_97; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_98; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_99; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_100; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_101; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_102; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_103; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_104; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_105; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_106; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_107; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_108; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_109; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_110; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_111; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_112; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_113; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_114; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_115; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_116; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_117; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_118; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_119; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_120; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_121; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_122; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_123; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_124; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_125; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_126; // @[pisa.scala 19:22]
  wire [7:0] init_io_pipe_phv_out_data_127; // @[pisa.scala 19:22]
  wire  PAR_clock; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_0; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_1; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_2; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_3; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_4; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_5; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_6; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_7; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_8; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_9; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_10; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_11; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_12; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_13; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_14; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_15; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_16; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_17; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_18; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_19; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_20; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_21; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_22; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_23; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_24; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_25; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_26; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_27; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_28; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_29; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_30; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_31; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_32; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_33; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_34; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_35; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_36; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_37; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_38; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_39; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_40; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_41; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_42; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_43; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_44; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_45; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_46; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_47; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_48; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_49; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_50; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_51; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_52; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_53; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_54; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_55; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_56; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_57; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_58; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_59; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_60; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_61; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_62; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_63; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_64; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_65; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_66; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_67; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_68; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_69; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_70; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_71; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_72; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_73; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_74; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_75; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_76; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_77; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_78; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_79; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_80; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_81; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_82; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_83; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_84; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_85; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_86; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_87; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_88; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_89; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_90; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_91; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_92; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_93; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_94; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_95; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_96; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_97; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_98; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_99; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_100; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_101; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_102; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_103; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_104; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_105; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_106; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_107; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_108; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_109; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_110; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_111; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_112; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_113; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_114; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_115; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_116; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_117; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_118; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_119; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_120; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_121; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_122; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_123; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_124; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_125; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_126; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_in_data_127; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_0; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_1; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_2; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_3; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_4; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_5; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_6; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_7; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_8; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_9; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_10; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_11; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_12; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_13; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_14; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_15; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_16; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_17; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_18; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_19; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_20; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_21; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_22; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_23; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_24; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_25; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_26; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_27; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_28; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_29; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_30; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_31; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_32; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_33; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_34; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_35; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_36; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_37; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_38; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_39; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_40; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_41; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_42; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_43; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_44; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_45; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_46; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_47; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_48; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_49; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_50; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_51; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_52; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_53; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_54; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_55; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_56; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_57; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_58; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_59; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_60; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_61; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_62; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_63; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_64; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_65; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_66; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_67; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_68; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_69; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_70; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_71; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_72; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_73; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_74; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_75; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_76; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_77; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_78; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_79; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_80; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_81; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_82; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_83; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_84; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_85; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_86; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_87; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_88; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_89; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_90; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_91; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_92; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_93; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_94; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_95; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_96; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_97; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_98; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_99; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_100; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_101; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_102; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_103; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_104; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_105; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_106; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_107; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_108; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_109; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_110; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_111; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_112; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_113; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_114; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_115; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_116; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_117; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_118; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_119; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_120; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_121; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_122; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_123; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_124; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_125; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_126; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_127; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_128; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_129; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_130; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_131; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_132; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_133; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_134; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_135; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_136; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_137; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_138; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_139; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_140; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_141; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_142; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_143; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_144; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_145; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_146; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_147; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_148; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_149; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_150; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_151; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_152; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_153; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_154; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_155; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_156; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_157; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_158; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_pipe_phv_out_data_159; // @[pisa.scala 23:21]
  wire [3:0] PAR_io_pipe_phv_out_next_processor_id; // @[pisa.scala 23:21]
  wire  PAR_io_pipe_phv_out_next_config_id; // @[pisa.scala 23:21]
  wire  PAR_io_pipe_phv_out_valid; // @[pisa.scala 23:21]
  wire  PAR_io_mod_en; // @[pisa.scala 23:21]
  wire  PAR_io_mod_last_mau_id_mod; // @[pisa.scala 23:21]
  wire [3:0] PAR_io_mod_last_mau_id; // @[pisa.scala 23:21]
  wire [2:0] PAR_io_mod_cs; // @[pisa.scala 23:21]
  wire  PAR_io_mod_module_mod_state_id_mod; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_mod_module_mod_state_id; // @[pisa.scala 23:21]
  wire  PAR_io_mod_module_mod_sram_w_cs; // @[pisa.scala 23:21]
  wire  PAR_io_mod_module_mod_sram_w_en; // @[pisa.scala 23:21]
  wire [7:0] PAR_io_mod_module_mod_sram_w_addr; // @[pisa.scala 23:21]
  wire [63:0] PAR_io_mod_module_mod_sram_w_data; // @[pisa.scala 23:21]
  wire  proc_0_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_0_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_0_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_0_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_0_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_0_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_0_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_0_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_0_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_0_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_0_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_0_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_0_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_0_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_0_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_1_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_1_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_1_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_1_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_1_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_1_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_1_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_1_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_1_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_1_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_1_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_1_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_1_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_1_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_1_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_2_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_2_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_2_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_2_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_2_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_2_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_2_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_2_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_2_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_2_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_2_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_2_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_2_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_2_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_2_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_3_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_3_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_3_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_3_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_3_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_3_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_3_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_3_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_3_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_3_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_3_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_3_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_3_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_3_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_3_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_4_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_4_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_4_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_4_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_4_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_4_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_4_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_4_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_4_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_4_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_4_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_4_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_4_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_4_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_4_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_5_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_5_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_5_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_5_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_5_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_5_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_5_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_5_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_5_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_5_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_5_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_5_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_5_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_5_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_5_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_6_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_6_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_6_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_6_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_6_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_6_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_6_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_6_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_6_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_6_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_6_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_6_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_6_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_6_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_6_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_7_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_7_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_7_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_7_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_7_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_7_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_7_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_7_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_7_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_7_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_7_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_7_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_7_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_7_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_7_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_8_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_8_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_8_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_8_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_8_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_8_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_8_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_8_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_8_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_8_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_8_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_8_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_8_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_8_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_8_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_9_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_9_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_9_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_9_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_9_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_9_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_9_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_9_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_9_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_9_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_9_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_9_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_9_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_9_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_9_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_10_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_10_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_10_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_10_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_10_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_10_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_10_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_10_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_10_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_10_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_10_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_10_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_10_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_10_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_10_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_11_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_11_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_11_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_11_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_11_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_11_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_11_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_11_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_11_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_11_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_11_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_11_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_11_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_11_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_11_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_12_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_12_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_12_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_12_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_12_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_12_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_12_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_12_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_12_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_12_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_12_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_12_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_12_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_12_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_12_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_12_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_12_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_12_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_12_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_12_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_12_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_12_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_13_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_13_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_13_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_13_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_13_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_13_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_13_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_13_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_13_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_13_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_13_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_13_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_13_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_13_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_13_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_13_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_13_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_13_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_13_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_13_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_13_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_13_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_14_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_14_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_14_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_14_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_14_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_14_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_14_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_14_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_14_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_14_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_14_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_14_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_14_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_14_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_14_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_14_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_14_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_14_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_14_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_14_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_14_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_14_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  wire  proc_15_clock; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_in_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_15_io_pipe_phv_in_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_15_io_pipe_phv_in_next_config_id; // @[pisa.scala 28:25]
  wire  proc_15_io_pipe_phv_in_is_valid_processor; // @[pisa.scala 28:25]
  wire  proc_15_io_pipe_phv_in_valid; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_0; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_1; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_2; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_3; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_4; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_5; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_6; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_7; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_8; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_9; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_10; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_11; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_12; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_13; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_14; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_15; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_16; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_17; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_18; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_19; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_20; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_21; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_22; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_23; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_24; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_25; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_26; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_27; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_28; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_29; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_30; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_31; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_32; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_33; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_34; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_35; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_36; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_37; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_38; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_39; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_40; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_41; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_42; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_43; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_44; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_45; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_46; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_47; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_48; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_49; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_50; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_51; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_52; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_53; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_54; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_55; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_56; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_57; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_58; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_59; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_60; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_61; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_62; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_63; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_64; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_65; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_66; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_67; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_68; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_69; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_70; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_71; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_72; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_73; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_74; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_75; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_76; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_77; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_78; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_79; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_80; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_81; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_82; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_83; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_84; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_85; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_86; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_87; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_88; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_89; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_90; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_91; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_92; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_93; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_94; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_95; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_96; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_97; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_98; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_99; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_100; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_101; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_102; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_103; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_104; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_105; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_106; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_107; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_108; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_109; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_110; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_111; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_112; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_113; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_114; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_115; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_116; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_117; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_118; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_119; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_120; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_121; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_122; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_123; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_124; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_125; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_126; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_127; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_128; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_129; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_130; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_131; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_132; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_133; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_134; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_135; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_136; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_137; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_138; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_139; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_140; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_141; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_142; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_143; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_144; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_145; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_146; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_147; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_148; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_149; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_150; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_151; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_152; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_153; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_154; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_155; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_156; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_157; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_158; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_pipe_phv_out_data_159; // @[pisa.scala 28:25]
  wire [3:0] proc_15_io_pipe_phv_out_next_processor_id; // @[pisa.scala 28:25]
  wire  proc_15_io_pipe_phv_out_next_config_id; // @[pisa.scala 28:25]
  wire  proc_15_io_pipe_phv_out_valid; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_en; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_config_id; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_key_mod_en; // @[pisa.scala 28:25]
  wire [2:0] proc_15_io_mod_mat_mod_key_mod_group_index; // @[pisa.scala 28:25]
  wire [1:0] proc_15_io_mod_mat_mod_key_mod_group_config; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_key_mod_group_mask_0; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_key_mod_group_mask_1; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_key_mod_group_mask_2; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_key_mod_group_mask_3; // @[pisa.scala 28:25]
  wire [6:0] proc_15_io_mod_mat_mod_key_mod_group_id_0; // @[pisa.scala 28:25]
  wire [6:0] proc_15_io_mod_mat_mod_key_mod_group_id_1; // @[pisa.scala 28:25]
  wire [6:0] proc_15_io_mod_mat_mod_key_mod_group_id_2; // @[pisa.scala 28:25]
  wire [6:0] proc_15_io_mod_mat_mod_key_mod_group_id_3; // @[pisa.scala 28:25]
  wire [4:0] proc_15_io_mod_mat_mod_table_mod_table_depth; // @[pisa.scala 28:25]
  wire [4:0] proc_15_io_mod_mat_mod_table_mod_table_width; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_mat_mod_w_en; // @[pisa.scala 28:25]
  wire [3:0] proc_15_io_mod_mat_mod_w_sram_id; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_mod_mat_mod_w_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_15_io_mod_mat_mod_w_data; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_exe_mod_en_0; // @[pisa.scala 28:25]
  wire  proc_15_io_mod_exe_mod_en_1; // @[pisa.scala 28:25]
  wire [7:0] proc_15_io_mod_exe_mod_addr; // @[pisa.scala 28:25]
  wire [63:0] proc_15_io_mod_exe_mod_data_0; // @[pisa.scala 28:25]
  wire [63:0] proc_15_io_mod_exe_mod_data_1; // @[pisa.scala 28:25]
  Initializer init ( // @[pisa.scala 19:22]
    .clock(init_clock),
    .io_pipe_phv_in_data_0(init_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(init_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(init_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(init_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(init_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(init_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(init_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(init_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(init_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(init_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(init_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(init_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(init_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(init_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(init_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(init_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(init_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(init_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(init_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(init_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(init_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(init_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(init_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(init_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(init_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(init_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(init_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(init_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(init_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(init_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(init_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(init_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(init_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(init_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(init_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(init_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(init_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(init_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(init_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(init_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(init_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(init_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(init_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(init_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(init_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(init_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(init_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(init_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(init_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(init_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(init_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(init_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(init_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(init_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(init_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(init_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(init_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(init_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(init_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(init_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(init_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(init_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(init_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(init_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(init_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(init_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(init_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(init_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(init_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(init_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(init_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(init_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(init_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(init_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(init_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(init_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(init_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(init_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(init_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(init_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(init_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(init_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(init_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(init_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(init_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(init_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(init_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(init_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(init_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(init_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(init_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(init_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(init_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(init_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(init_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(init_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(init_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(init_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(init_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(init_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(init_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(init_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(init_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(init_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(init_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(init_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(init_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(init_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(init_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(init_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(init_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(init_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(init_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(init_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(init_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(init_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(init_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(init_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(init_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(init_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(init_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(init_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(init_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(init_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(init_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(init_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(init_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(init_io_pipe_phv_in_data_127),
    .io_pipe_phv_out_data_0(init_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(init_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(init_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(init_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(init_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(init_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(init_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(init_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(init_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(init_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(init_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(init_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(init_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(init_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(init_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(init_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(init_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(init_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(init_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(init_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(init_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(init_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(init_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(init_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(init_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(init_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(init_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(init_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(init_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(init_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(init_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(init_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(init_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(init_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(init_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(init_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(init_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(init_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(init_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(init_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(init_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(init_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(init_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(init_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(init_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(init_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(init_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(init_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(init_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(init_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(init_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(init_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(init_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(init_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(init_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(init_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(init_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(init_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(init_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(init_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(init_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(init_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(init_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(init_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(init_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(init_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(init_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(init_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(init_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(init_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(init_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(init_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(init_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(init_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(init_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(init_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(init_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(init_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(init_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(init_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(init_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(init_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(init_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(init_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(init_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(init_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(init_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(init_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(init_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(init_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(init_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(init_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(init_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(init_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(init_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(init_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(init_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(init_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(init_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(init_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(init_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(init_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(init_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(init_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(init_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(init_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(init_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(init_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(init_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(init_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(init_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(init_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(init_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(init_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(init_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(init_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(init_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(init_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(init_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(init_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(init_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(init_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(init_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(init_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(init_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(init_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(init_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(init_io_pipe_phv_out_data_127)
  );
  ParserPISA PAR ( // @[pisa.scala 23:21]
    .clock(PAR_clock),
    .io_pipe_phv_in_data_0(PAR_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(PAR_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(PAR_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(PAR_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(PAR_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(PAR_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(PAR_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(PAR_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(PAR_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(PAR_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(PAR_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(PAR_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(PAR_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(PAR_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(PAR_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(PAR_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(PAR_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(PAR_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(PAR_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(PAR_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(PAR_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(PAR_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(PAR_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(PAR_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(PAR_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(PAR_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(PAR_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(PAR_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(PAR_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(PAR_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(PAR_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(PAR_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(PAR_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(PAR_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(PAR_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(PAR_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(PAR_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(PAR_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(PAR_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(PAR_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(PAR_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(PAR_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(PAR_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(PAR_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(PAR_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(PAR_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(PAR_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(PAR_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(PAR_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(PAR_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(PAR_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(PAR_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(PAR_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(PAR_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(PAR_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(PAR_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(PAR_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(PAR_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(PAR_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(PAR_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(PAR_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(PAR_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(PAR_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(PAR_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(PAR_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(PAR_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(PAR_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(PAR_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(PAR_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(PAR_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(PAR_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(PAR_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(PAR_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(PAR_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(PAR_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(PAR_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(PAR_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(PAR_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(PAR_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(PAR_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(PAR_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(PAR_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(PAR_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(PAR_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(PAR_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(PAR_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(PAR_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(PAR_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(PAR_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(PAR_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(PAR_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(PAR_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(PAR_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(PAR_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(PAR_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(PAR_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(PAR_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(PAR_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(PAR_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(PAR_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(PAR_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(PAR_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(PAR_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(PAR_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(PAR_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(PAR_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(PAR_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(PAR_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(PAR_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(PAR_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(PAR_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(PAR_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(PAR_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(PAR_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(PAR_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(PAR_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(PAR_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(PAR_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(PAR_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(PAR_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(PAR_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(PAR_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(PAR_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(PAR_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(PAR_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(PAR_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(PAR_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(PAR_io_pipe_phv_in_data_127),
    .io_pipe_phv_out_data_0(PAR_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(PAR_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(PAR_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(PAR_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(PAR_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(PAR_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(PAR_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(PAR_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(PAR_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(PAR_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(PAR_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(PAR_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(PAR_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(PAR_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(PAR_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(PAR_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(PAR_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(PAR_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(PAR_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(PAR_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(PAR_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(PAR_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(PAR_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(PAR_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(PAR_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(PAR_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(PAR_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(PAR_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(PAR_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(PAR_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(PAR_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(PAR_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(PAR_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(PAR_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(PAR_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(PAR_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(PAR_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(PAR_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(PAR_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(PAR_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(PAR_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(PAR_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(PAR_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(PAR_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(PAR_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(PAR_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(PAR_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(PAR_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(PAR_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(PAR_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(PAR_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(PAR_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(PAR_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(PAR_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(PAR_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(PAR_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(PAR_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(PAR_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(PAR_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(PAR_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(PAR_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(PAR_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(PAR_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(PAR_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(PAR_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(PAR_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(PAR_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(PAR_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(PAR_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(PAR_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(PAR_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(PAR_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(PAR_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(PAR_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(PAR_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(PAR_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(PAR_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(PAR_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(PAR_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(PAR_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(PAR_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(PAR_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(PAR_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(PAR_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(PAR_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(PAR_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(PAR_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(PAR_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(PAR_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(PAR_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(PAR_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(PAR_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(PAR_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(PAR_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(PAR_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(PAR_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(PAR_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(PAR_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(PAR_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(PAR_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(PAR_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(PAR_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(PAR_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(PAR_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(PAR_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(PAR_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(PAR_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(PAR_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(PAR_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(PAR_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(PAR_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(PAR_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(PAR_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(PAR_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(PAR_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(PAR_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(PAR_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(PAR_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(PAR_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(PAR_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(PAR_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(PAR_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(PAR_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(PAR_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(PAR_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(PAR_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(PAR_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(PAR_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(PAR_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(PAR_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(PAR_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(PAR_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(PAR_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(PAR_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(PAR_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(PAR_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(PAR_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(PAR_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(PAR_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(PAR_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(PAR_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(PAR_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(PAR_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(PAR_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(PAR_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(PAR_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(PAR_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(PAR_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(PAR_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(PAR_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(PAR_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(PAR_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(PAR_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(PAR_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(PAR_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(PAR_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(PAR_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(PAR_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(PAR_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(PAR_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(PAR_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(PAR_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(PAR_io_pipe_phv_out_valid),
    .io_mod_en(PAR_io_mod_en),
    .io_mod_last_mau_id_mod(PAR_io_mod_last_mau_id_mod),
    .io_mod_last_mau_id(PAR_io_mod_last_mau_id),
    .io_mod_cs(PAR_io_mod_cs),
    .io_mod_module_mod_state_id_mod(PAR_io_mod_module_mod_state_id_mod),
    .io_mod_module_mod_state_id(PAR_io_mod_module_mod_state_id),
    .io_mod_module_mod_sram_w_cs(PAR_io_mod_module_mod_sram_w_cs),
    .io_mod_module_mod_sram_w_en(PAR_io_mod_module_mod_sram_w_en),
    .io_mod_module_mod_sram_w_addr(PAR_io_mod_module_mod_sram_w_addr),
    .io_mod_module_mod_sram_w_data(PAR_io_mod_module_mod_sram_w_data)
  );
  ProcessorPISA proc_0 ( // @[pisa.scala 28:25]
    .clock(proc_0_clock),
    .io_pipe_phv_in_data_0(proc_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_0_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_0_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_0_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_0_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_0_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_0_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_0_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_0_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_0_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_0_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_0_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_0_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_0_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_0_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_0_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_0_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_0_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_0_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_0_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_0_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_0_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_0_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_0_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_0_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_0_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_0_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_1 ( // @[pisa.scala 28:25]
    .clock(proc_1_clock),
    .io_pipe_phv_in_data_0(proc_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_1_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_1_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_1_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_1_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_1_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_1_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_1_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_1_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_1_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_1_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_1_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_1_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_1_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_1_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_1_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_1_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_1_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_1_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_1_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_1_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_1_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_1_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_1_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_1_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_1_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_1_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_2 ( // @[pisa.scala 28:25]
    .clock(proc_2_clock),
    .io_pipe_phv_in_data_0(proc_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_2_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_2_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_2_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_2_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_2_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_2_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_2_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_2_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_2_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_2_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_2_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_2_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_2_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_2_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_2_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_2_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_2_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_2_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_2_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_2_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_2_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_2_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_2_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_2_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_2_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_2_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_3 ( // @[pisa.scala 28:25]
    .clock(proc_3_clock),
    .io_pipe_phv_in_data_0(proc_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_3_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_3_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_3_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_3_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_3_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_3_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_3_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_3_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_3_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_3_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_3_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_3_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_3_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_3_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_3_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_3_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_3_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_3_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_3_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_3_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_3_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_3_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_3_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_3_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_3_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_3_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_4 ( // @[pisa.scala 28:25]
    .clock(proc_4_clock),
    .io_pipe_phv_in_data_0(proc_4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_4_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_4_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_4_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_4_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_4_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_4_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_4_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_4_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_4_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_4_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_4_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_4_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_4_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_4_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_4_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_4_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_4_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_4_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_4_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_4_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_4_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_4_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_4_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_4_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_4_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_4_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_5 ( // @[pisa.scala 28:25]
    .clock(proc_5_clock),
    .io_pipe_phv_in_data_0(proc_5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_5_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_5_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_5_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_5_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_5_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_5_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_5_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_5_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_5_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_5_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_5_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_5_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_5_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_5_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_5_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_5_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_5_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_5_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_5_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_5_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_5_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_5_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_5_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_5_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_5_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_5_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_6 ( // @[pisa.scala 28:25]
    .clock(proc_6_clock),
    .io_pipe_phv_in_data_0(proc_6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_6_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_6_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_6_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_6_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_6_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_6_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_6_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_6_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_6_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_6_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_6_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_6_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_6_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_6_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_6_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_6_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_6_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_6_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_6_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_6_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_6_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_6_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_6_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_6_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_6_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_6_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_7 ( // @[pisa.scala 28:25]
    .clock(proc_7_clock),
    .io_pipe_phv_in_data_0(proc_7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_7_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_7_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_7_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_7_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_7_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_7_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_7_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_7_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_7_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_7_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_7_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_7_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_7_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_7_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_7_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_7_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_7_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_7_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_7_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_7_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_7_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_7_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_7_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_7_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_7_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_7_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_8 ( // @[pisa.scala 28:25]
    .clock(proc_8_clock),
    .io_pipe_phv_in_data_0(proc_8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_8_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_8_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_8_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_8_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_8_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_8_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_8_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_8_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_8_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_8_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_8_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_8_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_8_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_8_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_8_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_8_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_8_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_8_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_8_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_8_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_8_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_8_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_8_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_8_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_8_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_8_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_9 ( // @[pisa.scala 28:25]
    .clock(proc_9_clock),
    .io_pipe_phv_in_data_0(proc_9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_9_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_9_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_9_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_9_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_9_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_9_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_9_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_9_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_9_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_9_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_9_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_9_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_9_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_9_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_9_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_9_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_9_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_9_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_9_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_9_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_9_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_9_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_9_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_9_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_9_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_9_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_9_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_9_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_9_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_9_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_9_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_9_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_9_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_9_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_9_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_9_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_9_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_9_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_9_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_9_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_9_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_9_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_9_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_9_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_9_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_9_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_9_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_9_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_9_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_9_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_9_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_9_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_9_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_9_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_9_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_9_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_9_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_9_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_9_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_9_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_9_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_9_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_9_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_9_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_9_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_9_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_9_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_9_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_9_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_9_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_9_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_9_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_9_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_9_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_9_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_9_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_9_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_9_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_9_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_9_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_9_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_9_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_9_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_9_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_9_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_9_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_9_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_9_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_9_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_9_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_9_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_9_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_9_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_9_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_9_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_9_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_9_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_9_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_9_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_9_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_9_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_9_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_9_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_9_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_9_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_9_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_9_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_9_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_9_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_9_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_9_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_9_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_9_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_9_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_9_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_9_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_9_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_9_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_9_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_9_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_9_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_9_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_9_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_9_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_9_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_9_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_9_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_9_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_9_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_9_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_9_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_9_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_9_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_9_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_9_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_9_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_9_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_9_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_9_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_9_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_9_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_9_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_9_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_9_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_9_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_9_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_9_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_9_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_9_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_9_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_9_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_9_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_9_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_9_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_10 ( // @[pisa.scala 28:25]
    .clock(proc_10_clock),
    .io_pipe_phv_in_data_0(proc_10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_10_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_10_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_10_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_10_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_10_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_10_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_10_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_10_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_10_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_10_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_10_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_10_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_10_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_10_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_10_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_10_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_10_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_10_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_10_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_10_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_10_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_10_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_10_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_10_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_10_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_10_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_10_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_10_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_10_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_10_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_10_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_10_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_10_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_10_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_10_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_10_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_10_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_10_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_10_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_10_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_10_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_10_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_10_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_10_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_10_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_10_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_10_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_10_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_10_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_10_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_10_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_10_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_10_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_10_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_10_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_10_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_10_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_10_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_10_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_10_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_10_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_10_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_10_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_10_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_10_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_10_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_10_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_10_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_10_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_10_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_10_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_10_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_10_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_10_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_10_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_10_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_10_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_10_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_10_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_10_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_10_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_10_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_10_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_10_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_10_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_10_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_10_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_10_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_10_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_10_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_10_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_10_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_10_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_10_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_10_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_10_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_10_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_10_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_10_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_10_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_10_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_10_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_10_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_10_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_10_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_10_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_10_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_10_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_10_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_10_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_10_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_10_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_10_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_10_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_10_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_10_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_10_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_10_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_10_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_10_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_10_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_10_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_10_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_10_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_10_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_10_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_10_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_10_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_10_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_10_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_10_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_10_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_10_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_10_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_10_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_10_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_10_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_10_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_10_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_10_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_10_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_10_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_10_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_10_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_10_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_10_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_10_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_10_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_10_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_10_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_10_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_10_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_10_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_10_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_11 ( // @[pisa.scala 28:25]
    .clock(proc_11_clock),
    .io_pipe_phv_in_data_0(proc_11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_11_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_11_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_11_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_11_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_11_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_11_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_11_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_11_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_11_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_11_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_11_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_11_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_11_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_11_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_11_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_11_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_11_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_11_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_11_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_11_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_11_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_11_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_11_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_11_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_11_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_11_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_11_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_11_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_11_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_11_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_11_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_11_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_11_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_11_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_11_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_11_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_11_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_11_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_11_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_11_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_11_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_11_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_11_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_11_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_11_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_11_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_11_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_11_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_11_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_11_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_11_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_11_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_11_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_11_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_11_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_11_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_11_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_11_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_11_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_11_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_11_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_11_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_11_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_11_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_11_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_11_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_11_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_11_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_11_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_11_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_11_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_11_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_11_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_11_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_11_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_11_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_11_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_11_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_11_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_11_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_11_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_11_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_11_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_11_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_11_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_11_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_11_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_11_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_11_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_11_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_11_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_11_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_11_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_11_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_11_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_11_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_11_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_11_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_11_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_11_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_11_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_11_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_11_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_11_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_11_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_11_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_11_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_11_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_11_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_11_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_11_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_11_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_11_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_11_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_11_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_11_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_11_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_11_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_11_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_11_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_11_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_11_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_11_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_11_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_11_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_11_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_11_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_11_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_11_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_11_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_11_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_11_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_11_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_11_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_11_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_11_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_11_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_11_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_11_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_11_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_11_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_11_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_11_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_11_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_11_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_11_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_11_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_11_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_11_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_11_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_11_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_11_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_11_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_11_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_12 ( // @[pisa.scala 28:25]
    .clock(proc_12_clock),
    .io_pipe_phv_in_data_0(proc_12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_12_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_12_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_12_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_12_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_12_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_12_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_12_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_12_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_12_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_12_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_12_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_12_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_12_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_12_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_12_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_12_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_12_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_12_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_12_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_12_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_12_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_12_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_12_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_12_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_12_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_12_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_12_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_12_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_12_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_12_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_12_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_12_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_12_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_12_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_12_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_12_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_12_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_12_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_12_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_12_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_12_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_12_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_12_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_12_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_12_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_12_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_12_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_12_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_12_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_12_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_12_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_12_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_12_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_12_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_12_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_12_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_12_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_12_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_12_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_12_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_12_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_12_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_12_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_12_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_12_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_12_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_12_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_12_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_12_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_12_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_12_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_12_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_12_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_12_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_12_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_12_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_12_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_12_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_12_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_12_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_12_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_12_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_12_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_12_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_12_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_12_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_12_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_12_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_12_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_12_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_12_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_12_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_12_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_12_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_12_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_12_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_12_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_12_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_12_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_12_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_12_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_12_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_12_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_12_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_12_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_12_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_12_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_12_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_12_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_12_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_12_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_12_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_12_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_12_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_12_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_12_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_12_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_12_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_12_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_12_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_12_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_12_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_12_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_12_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_12_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_12_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_12_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_12_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_12_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_12_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_12_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_12_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_12_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_12_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_12_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_12_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_12_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_12_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_12_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_12_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_12_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_12_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_12_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_12_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_12_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_12_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_12_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_12_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_12_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_12_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_12_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_12_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_12_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_12_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_12_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_13 ( // @[pisa.scala 28:25]
    .clock(proc_13_clock),
    .io_pipe_phv_in_data_0(proc_13_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_13_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_13_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_13_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_13_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_13_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_13_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_13_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_13_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_13_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_13_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_13_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_13_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_13_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_13_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_13_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_13_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_13_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_13_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_13_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_13_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_13_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_13_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_13_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_13_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_13_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_13_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_13_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_13_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_13_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_13_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_13_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_13_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_13_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_13_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_13_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_13_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_13_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_13_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_13_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_13_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_13_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_13_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_13_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_13_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_13_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_13_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_13_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_13_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_13_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_13_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_13_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_13_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_13_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_13_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_13_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_13_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_13_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_13_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_13_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_13_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_13_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_13_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_13_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_13_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_13_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_13_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_13_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_13_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_13_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_13_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_13_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_13_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_13_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_13_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_13_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_13_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_13_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_13_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_13_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_13_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_13_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_13_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_13_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_13_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_13_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_13_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_13_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_13_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_13_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_13_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_13_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_13_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_13_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_13_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_13_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_13_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_13_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_13_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_13_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_13_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_13_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_13_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_13_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_13_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_13_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_13_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_13_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_13_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_13_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_13_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_13_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_13_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_13_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_13_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_13_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_13_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_13_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_13_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_13_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_13_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_13_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_13_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_13_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_13_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_13_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_13_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_13_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_13_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_13_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_13_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_13_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_13_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_13_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_13_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_13_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_13_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_13_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_13_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_13_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_13_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_13_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_13_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_13_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_13_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_13_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_13_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_13_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_13_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_13_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_13_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_13_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_13_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_13_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_13_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_13_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_13_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_13_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_13_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_13_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_13_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_13_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_13_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_13_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_13_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_13_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_13_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_13_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_13_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_13_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_13_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_13_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_13_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_13_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_13_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_13_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_13_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_13_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_13_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_13_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_13_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_13_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_13_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_13_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_13_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_13_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_13_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_13_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_13_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_13_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_13_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_13_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_13_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_13_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_13_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_13_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_13_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_13_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_13_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_13_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_13_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_13_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_13_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_13_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_13_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_13_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_13_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_13_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_13_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_13_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_13_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_13_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_13_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_13_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_13_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_13_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_13_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_13_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_13_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_13_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_13_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_13_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_13_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_13_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_13_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_13_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_13_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_13_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_13_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_13_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_13_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_13_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_13_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_13_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_13_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_13_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_13_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_13_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_13_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_13_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_13_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_13_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_13_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_13_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_13_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_13_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_13_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_13_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_13_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_13_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_13_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_13_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_13_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_13_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_13_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_13_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_13_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_13_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_13_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_13_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_13_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_13_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_13_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_13_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_13_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_13_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_13_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_13_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_13_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_13_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_13_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_13_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_13_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_13_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_13_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_13_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_13_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_13_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_13_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_13_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_13_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_13_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_13_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_13_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_13_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_13_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_13_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_13_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_13_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_13_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_13_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_13_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_13_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_13_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_13_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_13_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_13_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_13_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_13_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_13_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_13_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_13_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_13_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_13_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_13_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_13_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_13_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_13_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_13_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_13_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_13_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_13_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_13_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_13_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_13_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_13_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_13_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_13_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_13_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_13_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_13_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_13_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_13_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_13_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_13_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_13_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_13_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_13_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_13_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_13_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_13_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_13_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_13_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_13_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_13_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_13_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_13_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_13_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_13_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_13_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_13_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_13_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_13_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_13_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_13_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_13_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_13_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_13_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_13_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_13_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_13_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_14 ( // @[pisa.scala 28:25]
    .clock(proc_14_clock),
    .io_pipe_phv_in_data_0(proc_14_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_14_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_14_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_14_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_14_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_14_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_14_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_14_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_14_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_14_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_14_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_14_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_14_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_14_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_14_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_14_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_14_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_14_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_14_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_14_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_14_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_14_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_14_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_14_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_14_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_14_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_14_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_14_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_14_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_14_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_14_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_14_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_14_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_14_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_14_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_14_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_14_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_14_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_14_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_14_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_14_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_14_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_14_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_14_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_14_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_14_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_14_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_14_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_14_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_14_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_14_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_14_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_14_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_14_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_14_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_14_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_14_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_14_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_14_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_14_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_14_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_14_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_14_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_14_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_14_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_14_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_14_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_14_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_14_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_14_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_14_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_14_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_14_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_14_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_14_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_14_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_14_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_14_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_14_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_14_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_14_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_14_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_14_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_14_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_14_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_14_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_14_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_14_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_14_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_14_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_14_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_14_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_14_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_14_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_14_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_14_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_14_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_14_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_14_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_14_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_14_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_14_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_14_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_14_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_14_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_14_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_14_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_14_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_14_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_14_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_14_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_14_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_14_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_14_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_14_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_14_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_14_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_14_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_14_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_14_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_14_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_14_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_14_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_14_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_14_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_14_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_14_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_14_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_14_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_14_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_14_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_14_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_14_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_14_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_14_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_14_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_14_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_14_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_14_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_14_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_14_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_14_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_14_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_14_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_14_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_14_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_14_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_14_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_14_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_14_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_14_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_14_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_14_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_14_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_14_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_14_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_14_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_14_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_14_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_14_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_14_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_14_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_14_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_14_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_14_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_14_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_14_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_14_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_14_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_14_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_14_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_14_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_14_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_14_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_14_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_14_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_14_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_14_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_14_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_14_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_14_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_14_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_14_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_14_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_14_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_14_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_14_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_14_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_14_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_14_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_14_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_14_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_14_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_14_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_14_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_14_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_14_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_14_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_14_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_14_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_14_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_14_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_14_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_14_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_14_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_14_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_14_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_14_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_14_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_14_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_14_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_14_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_14_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_14_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_14_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_14_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_14_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_14_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_14_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_14_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_14_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_14_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_14_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_14_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_14_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_14_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_14_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_14_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_14_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_14_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_14_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_14_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_14_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_14_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_14_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_14_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_14_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_14_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_14_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_14_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_14_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_14_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_14_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_14_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_14_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_14_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_14_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_14_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_14_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_14_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_14_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_14_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_14_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_14_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_14_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_14_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_14_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_14_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_14_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_14_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_14_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_14_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_14_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_14_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_14_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_14_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_14_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_14_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_14_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_14_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_14_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_14_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_14_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_14_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_14_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_14_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_14_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_14_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_14_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_14_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_14_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_14_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_14_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_14_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_14_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_14_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_14_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_14_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_14_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_14_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_14_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_14_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_14_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_14_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_14_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_14_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_14_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_14_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_14_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_14_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_14_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_14_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_14_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_14_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_14_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_14_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_14_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_14_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_14_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_14_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_14_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_14_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_14_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_14_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_14_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_14_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_14_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_14_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_14_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_14_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_14_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_14_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_14_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_14_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_14_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_14_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_14_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_14_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_14_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_14_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_14_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_14_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_14_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_14_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_14_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_14_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_14_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_14_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_14_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_14_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_14_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_14_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_14_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_14_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_14_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_14_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_14_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_14_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_14_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_14_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_14_io_mod_exe_mod_data_1)
  );
  ProcessorPISA proc_15 ( // @[pisa.scala 28:25]
    .clock(proc_15_clock),
    .io_pipe_phv_in_data_0(proc_15_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(proc_15_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(proc_15_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(proc_15_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(proc_15_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(proc_15_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(proc_15_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(proc_15_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(proc_15_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(proc_15_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(proc_15_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(proc_15_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(proc_15_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(proc_15_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(proc_15_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(proc_15_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(proc_15_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(proc_15_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(proc_15_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(proc_15_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(proc_15_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(proc_15_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(proc_15_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(proc_15_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(proc_15_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(proc_15_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(proc_15_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(proc_15_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(proc_15_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(proc_15_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(proc_15_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(proc_15_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(proc_15_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(proc_15_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(proc_15_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(proc_15_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(proc_15_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(proc_15_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(proc_15_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(proc_15_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(proc_15_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(proc_15_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(proc_15_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(proc_15_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(proc_15_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(proc_15_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(proc_15_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(proc_15_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(proc_15_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(proc_15_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(proc_15_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(proc_15_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(proc_15_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(proc_15_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(proc_15_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(proc_15_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(proc_15_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(proc_15_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(proc_15_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(proc_15_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(proc_15_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(proc_15_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(proc_15_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(proc_15_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(proc_15_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(proc_15_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(proc_15_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(proc_15_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(proc_15_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(proc_15_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(proc_15_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(proc_15_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(proc_15_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(proc_15_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(proc_15_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(proc_15_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(proc_15_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(proc_15_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(proc_15_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(proc_15_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(proc_15_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(proc_15_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(proc_15_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(proc_15_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(proc_15_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(proc_15_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(proc_15_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(proc_15_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(proc_15_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(proc_15_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(proc_15_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(proc_15_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(proc_15_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(proc_15_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(proc_15_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(proc_15_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(proc_15_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(proc_15_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(proc_15_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(proc_15_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(proc_15_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(proc_15_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(proc_15_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(proc_15_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(proc_15_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(proc_15_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(proc_15_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(proc_15_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(proc_15_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(proc_15_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(proc_15_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(proc_15_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(proc_15_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(proc_15_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(proc_15_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(proc_15_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(proc_15_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(proc_15_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(proc_15_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(proc_15_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(proc_15_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(proc_15_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(proc_15_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(proc_15_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(proc_15_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(proc_15_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(proc_15_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(proc_15_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(proc_15_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(proc_15_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(proc_15_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(proc_15_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(proc_15_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(proc_15_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(proc_15_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(proc_15_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(proc_15_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(proc_15_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(proc_15_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(proc_15_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(proc_15_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(proc_15_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(proc_15_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(proc_15_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(proc_15_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(proc_15_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(proc_15_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(proc_15_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(proc_15_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(proc_15_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(proc_15_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(proc_15_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(proc_15_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(proc_15_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(proc_15_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(proc_15_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(proc_15_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(proc_15_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(proc_15_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(proc_15_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_next_processor_id(proc_15_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(proc_15_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(proc_15_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(proc_15_io_pipe_phv_in_valid),
    .io_pipe_phv_out_data_0(proc_15_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(proc_15_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(proc_15_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(proc_15_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(proc_15_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(proc_15_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(proc_15_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(proc_15_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(proc_15_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(proc_15_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(proc_15_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(proc_15_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(proc_15_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(proc_15_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(proc_15_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(proc_15_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(proc_15_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(proc_15_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(proc_15_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(proc_15_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(proc_15_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(proc_15_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(proc_15_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(proc_15_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(proc_15_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(proc_15_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(proc_15_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(proc_15_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(proc_15_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(proc_15_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(proc_15_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(proc_15_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(proc_15_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(proc_15_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(proc_15_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(proc_15_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(proc_15_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(proc_15_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(proc_15_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(proc_15_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(proc_15_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(proc_15_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(proc_15_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(proc_15_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(proc_15_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(proc_15_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(proc_15_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(proc_15_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(proc_15_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(proc_15_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(proc_15_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(proc_15_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(proc_15_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(proc_15_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(proc_15_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(proc_15_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(proc_15_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(proc_15_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(proc_15_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(proc_15_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(proc_15_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(proc_15_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(proc_15_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(proc_15_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(proc_15_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(proc_15_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(proc_15_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(proc_15_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(proc_15_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(proc_15_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(proc_15_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(proc_15_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(proc_15_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(proc_15_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(proc_15_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(proc_15_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(proc_15_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(proc_15_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(proc_15_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(proc_15_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(proc_15_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(proc_15_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(proc_15_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(proc_15_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(proc_15_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(proc_15_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(proc_15_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(proc_15_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(proc_15_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(proc_15_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(proc_15_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(proc_15_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(proc_15_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(proc_15_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(proc_15_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(proc_15_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(proc_15_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(proc_15_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(proc_15_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(proc_15_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(proc_15_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(proc_15_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(proc_15_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(proc_15_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(proc_15_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(proc_15_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(proc_15_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(proc_15_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(proc_15_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(proc_15_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(proc_15_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(proc_15_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(proc_15_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(proc_15_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(proc_15_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(proc_15_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(proc_15_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(proc_15_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(proc_15_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(proc_15_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(proc_15_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(proc_15_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(proc_15_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(proc_15_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(proc_15_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(proc_15_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(proc_15_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(proc_15_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(proc_15_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(proc_15_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(proc_15_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(proc_15_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(proc_15_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(proc_15_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(proc_15_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(proc_15_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(proc_15_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(proc_15_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(proc_15_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(proc_15_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(proc_15_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(proc_15_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(proc_15_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(proc_15_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(proc_15_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(proc_15_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(proc_15_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(proc_15_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(proc_15_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(proc_15_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(proc_15_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(proc_15_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(proc_15_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(proc_15_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(proc_15_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(proc_15_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(proc_15_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(proc_15_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(proc_15_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(proc_15_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_next_processor_id(proc_15_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(proc_15_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(proc_15_io_pipe_phv_out_valid),
    .io_mod_mat_mod_en(proc_15_io_mod_mat_mod_en),
    .io_mod_mat_mod_config_id(proc_15_io_mod_mat_mod_config_id),
    .io_mod_mat_mod_key_mod_en(proc_15_io_mod_mat_mod_key_mod_en),
    .io_mod_mat_mod_key_mod_group_index(proc_15_io_mod_mat_mod_key_mod_group_index),
    .io_mod_mat_mod_key_mod_group_config(proc_15_io_mod_mat_mod_key_mod_group_config),
    .io_mod_mat_mod_key_mod_group_mask_0(proc_15_io_mod_mat_mod_key_mod_group_mask_0),
    .io_mod_mat_mod_key_mod_group_mask_1(proc_15_io_mod_mat_mod_key_mod_group_mask_1),
    .io_mod_mat_mod_key_mod_group_mask_2(proc_15_io_mod_mat_mod_key_mod_group_mask_2),
    .io_mod_mat_mod_key_mod_group_mask_3(proc_15_io_mod_mat_mod_key_mod_group_mask_3),
    .io_mod_mat_mod_key_mod_group_id_0(proc_15_io_mod_mat_mod_key_mod_group_id_0),
    .io_mod_mat_mod_key_mod_group_id_1(proc_15_io_mod_mat_mod_key_mod_group_id_1),
    .io_mod_mat_mod_key_mod_group_id_2(proc_15_io_mod_mat_mod_key_mod_group_id_2),
    .io_mod_mat_mod_key_mod_group_id_3(proc_15_io_mod_mat_mod_key_mod_group_id_3),
    .io_mod_mat_mod_table_mod_table_depth(proc_15_io_mod_mat_mod_table_mod_table_depth),
    .io_mod_mat_mod_table_mod_table_width(proc_15_io_mod_mat_mod_table_mod_table_width),
    .io_mod_mat_mod_w_en(proc_15_io_mod_mat_mod_w_en),
    .io_mod_mat_mod_w_sram_id(proc_15_io_mod_mat_mod_w_sram_id),
    .io_mod_mat_mod_w_addr(proc_15_io_mod_mat_mod_w_addr),
    .io_mod_mat_mod_w_data(proc_15_io_mod_mat_mod_w_data),
    .io_mod_exe_mod_en_0(proc_15_io_mod_exe_mod_en_0),
    .io_mod_exe_mod_en_1(proc_15_io_mod_exe_mod_en_1),
    .io_mod_exe_mod_addr(proc_15_io_mod_exe_mod_addr),
    .io_mod_exe_mod_data_0(proc_15_io_mod_exe_mod_data_0),
    .io_mod_exe_mod_data_1(proc_15_io_mod_exe_mod_data_1)
  );
  assign io_pipe_phv_out_data_0 = proc_15_io_pipe_phv_out_data_0; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_1 = proc_15_io_pipe_phv_out_data_1; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_2 = proc_15_io_pipe_phv_out_data_2; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_3 = proc_15_io_pipe_phv_out_data_3; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_4 = proc_15_io_pipe_phv_out_data_4; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_5 = proc_15_io_pipe_phv_out_data_5; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_6 = proc_15_io_pipe_phv_out_data_6; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_7 = proc_15_io_pipe_phv_out_data_7; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_8 = proc_15_io_pipe_phv_out_data_8; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_9 = proc_15_io_pipe_phv_out_data_9; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_10 = proc_15_io_pipe_phv_out_data_10; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_11 = proc_15_io_pipe_phv_out_data_11; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_12 = proc_15_io_pipe_phv_out_data_12; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_13 = proc_15_io_pipe_phv_out_data_13; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_14 = proc_15_io_pipe_phv_out_data_14; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_15 = proc_15_io_pipe_phv_out_data_15; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_16 = proc_15_io_pipe_phv_out_data_16; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_17 = proc_15_io_pipe_phv_out_data_17; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_18 = proc_15_io_pipe_phv_out_data_18; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_19 = proc_15_io_pipe_phv_out_data_19; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_20 = proc_15_io_pipe_phv_out_data_20; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_21 = proc_15_io_pipe_phv_out_data_21; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_22 = proc_15_io_pipe_phv_out_data_22; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_23 = proc_15_io_pipe_phv_out_data_23; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_24 = proc_15_io_pipe_phv_out_data_24; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_25 = proc_15_io_pipe_phv_out_data_25; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_26 = proc_15_io_pipe_phv_out_data_26; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_27 = proc_15_io_pipe_phv_out_data_27; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_28 = proc_15_io_pipe_phv_out_data_28; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_29 = proc_15_io_pipe_phv_out_data_29; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_30 = proc_15_io_pipe_phv_out_data_30; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_31 = proc_15_io_pipe_phv_out_data_31; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_32 = proc_15_io_pipe_phv_out_data_32; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_33 = proc_15_io_pipe_phv_out_data_33; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_34 = proc_15_io_pipe_phv_out_data_34; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_35 = proc_15_io_pipe_phv_out_data_35; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_36 = proc_15_io_pipe_phv_out_data_36; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_37 = proc_15_io_pipe_phv_out_data_37; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_38 = proc_15_io_pipe_phv_out_data_38; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_39 = proc_15_io_pipe_phv_out_data_39; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_40 = proc_15_io_pipe_phv_out_data_40; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_41 = proc_15_io_pipe_phv_out_data_41; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_42 = proc_15_io_pipe_phv_out_data_42; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_43 = proc_15_io_pipe_phv_out_data_43; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_44 = proc_15_io_pipe_phv_out_data_44; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_45 = proc_15_io_pipe_phv_out_data_45; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_46 = proc_15_io_pipe_phv_out_data_46; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_47 = proc_15_io_pipe_phv_out_data_47; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_48 = proc_15_io_pipe_phv_out_data_48; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_49 = proc_15_io_pipe_phv_out_data_49; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_50 = proc_15_io_pipe_phv_out_data_50; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_51 = proc_15_io_pipe_phv_out_data_51; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_52 = proc_15_io_pipe_phv_out_data_52; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_53 = proc_15_io_pipe_phv_out_data_53; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_54 = proc_15_io_pipe_phv_out_data_54; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_55 = proc_15_io_pipe_phv_out_data_55; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_56 = proc_15_io_pipe_phv_out_data_56; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_57 = proc_15_io_pipe_phv_out_data_57; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_58 = proc_15_io_pipe_phv_out_data_58; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_59 = proc_15_io_pipe_phv_out_data_59; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_60 = proc_15_io_pipe_phv_out_data_60; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_61 = proc_15_io_pipe_phv_out_data_61; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_62 = proc_15_io_pipe_phv_out_data_62; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_63 = proc_15_io_pipe_phv_out_data_63; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_64 = proc_15_io_pipe_phv_out_data_64; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_65 = proc_15_io_pipe_phv_out_data_65; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_66 = proc_15_io_pipe_phv_out_data_66; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_67 = proc_15_io_pipe_phv_out_data_67; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_68 = proc_15_io_pipe_phv_out_data_68; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_69 = proc_15_io_pipe_phv_out_data_69; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_70 = proc_15_io_pipe_phv_out_data_70; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_71 = proc_15_io_pipe_phv_out_data_71; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_72 = proc_15_io_pipe_phv_out_data_72; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_73 = proc_15_io_pipe_phv_out_data_73; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_74 = proc_15_io_pipe_phv_out_data_74; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_75 = proc_15_io_pipe_phv_out_data_75; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_76 = proc_15_io_pipe_phv_out_data_76; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_77 = proc_15_io_pipe_phv_out_data_77; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_78 = proc_15_io_pipe_phv_out_data_78; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_79 = proc_15_io_pipe_phv_out_data_79; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_80 = proc_15_io_pipe_phv_out_data_80; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_81 = proc_15_io_pipe_phv_out_data_81; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_82 = proc_15_io_pipe_phv_out_data_82; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_83 = proc_15_io_pipe_phv_out_data_83; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_84 = proc_15_io_pipe_phv_out_data_84; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_85 = proc_15_io_pipe_phv_out_data_85; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_86 = proc_15_io_pipe_phv_out_data_86; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_87 = proc_15_io_pipe_phv_out_data_87; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_88 = proc_15_io_pipe_phv_out_data_88; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_89 = proc_15_io_pipe_phv_out_data_89; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_90 = proc_15_io_pipe_phv_out_data_90; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_91 = proc_15_io_pipe_phv_out_data_91; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_92 = proc_15_io_pipe_phv_out_data_92; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_93 = proc_15_io_pipe_phv_out_data_93; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_94 = proc_15_io_pipe_phv_out_data_94; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_95 = proc_15_io_pipe_phv_out_data_95; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_96 = proc_15_io_pipe_phv_out_data_96; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_97 = proc_15_io_pipe_phv_out_data_97; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_98 = proc_15_io_pipe_phv_out_data_98; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_99 = proc_15_io_pipe_phv_out_data_99; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_100 = proc_15_io_pipe_phv_out_data_100; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_101 = proc_15_io_pipe_phv_out_data_101; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_102 = proc_15_io_pipe_phv_out_data_102; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_103 = proc_15_io_pipe_phv_out_data_103; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_104 = proc_15_io_pipe_phv_out_data_104; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_105 = proc_15_io_pipe_phv_out_data_105; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_106 = proc_15_io_pipe_phv_out_data_106; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_107 = proc_15_io_pipe_phv_out_data_107; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_108 = proc_15_io_pipe_phv_out_data_108; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_109 = proc_15_io_pipe_phv_out_data_109; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_110 = proc_15_io_pipe_phv_out_data_110; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_111 = proc_15_io_pipe_phv_out_data_111; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_112 = proc_15_io_pipe_phv_out_data_112; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_113 = proc_15_io_pipe_phv_out_data_113; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_114 = proc_15_io_pipe_phv_out_data_114; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_115 = proc_15_io_pipe_phv_out_data_115; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_116 = proc_15_io_pipe_phv_out_data_116; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_117 = proc_15_io_pipe_phv_out_data_117; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_118 = proc_15_io_pipe_phv_out_data_118; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_119 = proc_15_io_pipe_phv_out_data_119; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_120 = proc_15_io_pipe_phv_out_data_120; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_121 = proc_15_io_pipe_phv_out_data_121; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_122 = proc_15_io_pipe_phv_out_data_122; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_123 = proc_15_io_pipe_phv_out_data_123; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_124 = proc_15_io_pipe_phv_out_data_124; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_125 = proc_15_io_pipe_phv_out_data_125; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_126 = proc_15_io_pipe_phv_out_data_126; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_127 = proc_15_io_pipe_phv_out_data_127; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_128 = proc_15_io_pipe_phv_out_data_128; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_129 = proc_15_io_pipe_phv_out_data_129; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_130 = proc_15_io_pipe_phv_out_data_130; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_131 = proc_15_io_pipe_phv_out_data_131; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_132 = proc_15_io_pipe_phv_out_data_132; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_133 = proc_15_io_pipe_phv_out_data_133; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_134 = proc_15_io_pipe_phv_out_data_134; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_135 = proc_15_io_pipe_phv_out_data_135; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_136 = proc_15_io_pipe_phv_out_data_136; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_137 = proc_15_io_pipe_phv_out_data_137; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_138 = proc_15_io_pipe_phv_out_data_138; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_139 = proc_15_io_pipe_phv_out_data_139; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_140 = proc_15_io_pipe_phv_out_data_140; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_141 = proc_15_io_pipe_phv_out_data_141; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_142 = proc_15_io_pipe_phv_out_data_142; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_143 = proc_15_io_pipe_phv_out_data_143; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_144 = proc_15_io_pipe_phv_out_data_144; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_145 = proc_15_io_pipe_phv_out_data_145; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_146 = proc_15_io_pipe_phv_out_data_146; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_147 = proc_15_io_pipe_phv_out_data_147; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_148 = proc_15_io_pipe_phv_out_data_148; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_149 = proc_15_io_pipe_phv_out_data_149; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_150 = proc_15_io_pipe_phv_out_data_150; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_151 = proc_15_io_pipe_phv_out_data_151; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_152 = proc_15_io_pipe_phv_out_data_152; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_153 = proc_15_io_pipe_phv_out_data_153; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_154 = proc_15_io_pipe_phv_out_data_154; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_155 = proc_15_io_pipe_phv_out_data_155; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_156 = proc_15_io_pipe_phv_out_data_156; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_157 = proc_15_io_pipe_phv_out_data_157; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_158 = proc_15_io_pipe_phv_out_data_158; // @[pisa.scala 42:52]
  assign io_pipe_phv_out_data_159 = proc_15_io_pipe_phv_out_data_159; // @[pisa.scala 42:52]
  assign init_clock = clock;
  assign init_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[pisa.scala 20:25]
  assign init_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[pisa.scala 20:25]
  assign PAR_clock = clock;
  assign PAR_io_pipe_phv_in_data_0 = init_io_pipe_phv_out_data_0; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_1 = init_io_pipe_phv_out_data_1; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_2 = init_io_pipe_phv_out_data_2; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_3 = init_io_pipe_phv_out_data_3; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_4 = init_io_pipe_phv_out_data_4; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_5 = init_io_pipe_phv_out_data_5; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_6 = init_io_pipe_phv_out_data_6; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_7 = init_io_pipe_phv_out_data_7; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_8 = init_io_pipe_phv_out_data_8; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_9 = init_io_pipe_phv_out_data_9; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_10 = init_io_pipe_phv_out_data_10; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_11 = init_io_pipe_phv_out_data_11; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_12 = init_io_pipe_phv_out_data_12; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_13 = init_io_pipe_phv_out_data_13; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_14 = init_io_pipe_phv_out_data_14; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_15 = init_io_pipe_phv_out_data_15; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_16 = init_io_pipe_phv_out_data_16; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_17 = init_io_pipe_phv_out_data_17; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_18 = init_io_pipe_phv_out_data_18; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_19 = init_io_pipe_phv_out_data_19; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_20 = init_io_pipe_phv_out_data_20; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_21 = init_io_pipe_phv_out_data_21; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_22 = init_io_pipe_phv_out_data_22; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_23 = init_io_pipe_phv_out_data_23; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_24 = init_io_pipe_phv_out_data_24; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_25 = init_io_pipe_phv_out_data_25; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_26 = init_io_pipe_phv_out_data_26; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_27 = init_io_pipe_phv_out_data_27; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_28 = init_io_pipe_phv_out_data_28; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_29 = init_io_pipe_phv_out_data_29; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_30 = init_io_pipe_phv_out_data_30; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_31 = init_io_pipe_phv_out_data_31; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_32 = init_io_pipe_phv_out_data_32; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_33 = init_io_pipe_phv_out_data_33; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_34 = init_io_pipe_phv_out_data_34; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_35 = init_io_pipe_phv_out_data_35; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_36 = init_io_pipe_phv_out_data_36; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_37 = init_io_pipe_phv_out_data_37; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_38 = init_io_pipe_phv_out_data_38; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_39 = init_io_pipe_phv_out_data_39; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_40 = init_io_pipe_phv_out_data_40; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_41 = init_io_pipe_phv_out_data_41; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_42 = init_io_pipe_phv_out_data_42; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_43 = init_io_pipe_phv_out_data_43; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_44 = init_io_pipe_phv_out_data_44; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_45 = init_io_pipe_phv_out_data_45; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_46 = init_io_pipe_phv_out_data_46; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_47 = init_io_pipe_phv_out_data_47; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_48 = init_io_pipe_phv_out_data_48; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_49 = init_io_pipe_phv_out_data_49; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_50 = init_io_pipe_phv_out_data_50; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_51 = init_io_pipe_phv_out_data_51; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_52 = init_io_pipe_phv_out_data_52; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_53 = init_io_pipe_phv_out_data_53; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_54 = init_io_pipe_phv_out_data_54; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_55 = init_io_pipe_phv_out_data_55; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_56 = init_io_pipe_phv_out_data_56; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_57 = init_io_pipe_phv_out_data_57; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_58 = init_io_pipe_phv_out_data_58; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_59 = init_io_pipe_phv_out_data_59; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_60 = init_io_pipe_phv_out_data_60; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_61 = init_io_pipe_phv_out_data_61; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_62 = init_io_pipe_phv_out_data_62; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_63 = init_io_pipe_phv_out_data_63; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_64 = init_io_pipe_phv_out_data_64; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_65 = init_io_pipe_phv_out_data_65; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_66 = init_io_pipe_phv_out_data_66; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_67 = init_io_pipe_phv_out_data_67; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_68 = init_io_pipe_phv_out_data_68; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_69 = init_io_pipe_phv_out_data_69; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_70 = init_io_pipe_phv_out_data_70; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_71 = init_io_pipe_phv_out_data_71; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_72 = init_io_pipe_phv_out_data_72; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_73 = init_io_pipe_phv_out_data_73; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_74 = init_io_pipe_phv_out_data_74; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_75 = init_io_pipe_phv_out_data_75; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_76 = init_io_pipe_phv_out_data_76; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_77 = init_io_pipe_phv_out_data_77; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_78 = init_io_pipe_phv_out_data_78; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_79 = init_io_pipe_phv_out_data_79; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_80 = init_io_pipe_phv_out_data_80; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_81 = init_io_pipe_phv_out_data_81; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_82 = init_io_pipe_phv_out_data_82; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_83 = init_io_pipe_phv_out_data_83; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_84 = init_io_pipe_phv_out_data_84; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_85 = init_io_pipe_phv_out_data_85; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_86 = init_io_pipe_phv_out_data_86; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_87 = init_io_pipe_phv_out_data_87; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_88 = init_io_pipe_phv_out_data_88; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_89 = init_io_pipe_phv_out_data_89; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_90 = init_io_pipe_phv_out_data_90; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_91 = init_io_pipe_phv_out_data_91; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_92 = init_io_pipe_phv_out_data_92; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_93 = init_io_pipe_phv_out_data_93; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_94 = init_io_pipe_phv_out_data_94; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_95 = init_io_pipe_phv_out_data_95; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_96 = init_io_pipe_phv_out_data_96; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_97 = init_io_pipe_phv_out_data_97; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_98 = init_io_pipe_phv_out_data_98; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_99 = init_io_pipe_phv_out_data_99; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_100 = init_io_pipe_phv_out_data_100; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_101 = init_io_pipe_phv_out_data_101; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_102 = init_io_pipe_phv_out_data_102; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_103 = init_io_pipe_phv_out_data_103; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_104 = init_io_pipe_phv_out_data_104; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_105 = init_io_pipe_phv_out_data_105; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_106 = init_io_pipe_phv_out_data_106; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_107 = init_io_pipe_phv_out_data_107; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_108 = init_io_pipe_phv_out_data_108; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_109 = init_io_pipe_phv_out_data_109; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_110 = init_io_pipe_phv_out_data_110; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_111 = init_io_pipe_phv_out_data_111; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_112 = init_io_pipe_phv_out_data_112; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_113 = init_io_pipe_phv_out_data_113; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_114 = init_io_pipe_phv_out_data_114; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_115 = init_io_pipe_phv_out_data_115; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_116 = init_io_pipe_phv_out_data_116; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_117 = init_io_pipe_phv_out_data_117; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_118 = init_io_pipe_phv_out_data_118; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_119 = init_io_pipe_phv_out_data_119; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_120 = init_io_pipe_phv_out_data_120; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_121 = init_io_pipe_phv_out_data_121; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_122 = init_io_pipe_phv_out_data_122; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_123 = init_io_pipe_phv_out_data_123; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_124 = init_io_pipe_phv_out_data_124; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_125 = init_io_pipe_phv_out_data_125; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_126 = init_io_pipe_phv_out_data_126; // @[pisa.scala 24:24]
  assign PAR_io_pipe_phv_in_data_127 = init_io_pipe_phv_out_data_127; // @[pisa.scala 24:24]
  assign PAR_io_mod_en = io_mod_par_mod_en; // @[pisa.scala 25:16]
  assign PAR_io_mod_last_mau_id_mod = io_mod_par_mod_last_mau_id_mod; // @[pisa.scala 25:16]
  assign PAR_io_mod_last_mau_id = io_mod_par_mod_last_mau_id; // @[pisa.scala 25:16]
  assign PAR_io_mod_cs = io_mod_par_mod_cs; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_state_id_mod = io_mod_par_mod_module_mod_state_id_mod; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_state_id = io_mod_par_mod_module_mod_state_id; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_cs = io_mod_par_mod_module_mod_sram_w_cs; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_en = io_mod_par_mod_module_mod_sram_w_en; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_addr = io_mod_par_mod_module_mod_sram_w_addr; // @[pisa.scala 25:16]
  assign PAR_io_mod_module_mod_sram_w_data = io_mod_par_mod_module_mod_sram_w_data; // @[pisa.scala 25:16]
  assign proc_0_clock = clock;
  assign proc_0_io_pipe_phv_in_data_0 = PAR_io_pipe_phv_out_data_0; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_1 = PAR_io_pipe_phv_out_data_1; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_2 = PAR_io_pipe_phv_out_data_2; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_3 = PAR_io_pipe_phv_out_data_3; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_4 = PAR_io_pipe_phv_out_data_4; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_5 = PAR_io_pipe_phv_out_data_5; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_6 = PAR_io_pipe_phv_out_data_6; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_7 = PAR_io_pipe_phv_out_data_7; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_8 = PAR_io_pipe_phv_out_data_8; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_9 = PAR_io_pipe_phv_out_data_9; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_10 = PAR_io_pipe_phv_out_data_10; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_11 = PAR_io_pipe_phv_out_data_11; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_12 = PAR_io_pipe_phv_out_data_12; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_13 = PAR_io_pipe_phv_out_data_13; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_14 = PAR_io_pipe_phv_out_data_14; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_15 = PAR_io_pipe_phv_out_data_15; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_16 = PAR_io_pipe_phv_out_data_16; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_17 = PAR_io_pipe_phv_out_data_17; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_18 = PAR_io_pipe_phv_out_data_18; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_19 = PAR_io_pipe_phv_out_data_19; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_20 = PAR_io_pipe_phv_out_data_20; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_21 = PAR_io_pipe_phv_out_data_21; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_22 = PAR_io_pipe_phv_out_data_22; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_23 = PAR_io_pipe_phv_out_data_23; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_24 = PAR_io_pipe_phv_out_data_24; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_25 = PAR_io_pipe_phv_out_data_25; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_26 = PAR_io_pipe_phv_out_data_26; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_27 = PAR_io_pipe_phv_out_data_27; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_28 = PAR_io_pipe_phv_out_data_28; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_29 = PAR_io_pipe_phv_out_data_29; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_30 = PAR_io_pipe_phv_out_data_30; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_31 = PAR_io_pipe_phv_out_data_31; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_32 = PAR_io_pipe_phv_out_data_32; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_33 = PAR_io_pipe_phv_out_data_33; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_34 = PAR_io_pipe_phv_out_data_34; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_35 = PAR_io_pipe_phv_out_data_35; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_36 = PAR_io_pipe_phv_out_data_36; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_37 = PAR_io_pipe_phv_out_data_37; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_38 = PAR_io_pipe_phv_out_data_38; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_39 = PAR_io_pipe_phv_out_data_39; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_40 = PAR_io_pipe_phv_out_data_40; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_41 = PAR_io_pipe_phv_out_data_41; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_42 = PAR_io_pipe_phv_out_data_42; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_43 = PAR_io_pipe_phv_out_data_43; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_44 = PAR_io_pipe_phv_out_data_44; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_45 = PAR_io_pipe_phv_out_data_45; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_46 = PAR_io_pipe_phv_out_data_46; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_47 = PAR_io_pipe_phv_out_data_47; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_48 = PAR_io_pipe_phv_out_data_48; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_49 = PAR_io_pipe_phv_out_data_49; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_50 = PAR_io_pipe_phv_out_data_50; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_51 = PAR_io_pipe_phv_out_data_51; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_52 = PAR_io_pipe_phv_out_data_52; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_53 = PAR_io_pipe_phv_out_data_53; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_54 = PAR_io_pipe_phv_out_data_54; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_55 = PAR_io_pipe_phv_out_data_55; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_56 = PAR_io_pipe_phv_out_data_56; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_57 = PAR_io_pipe_phv_out_data_57; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_58 = PAR_io_pipe_phv_out_data_58; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_59 = PAR_io_pipe_phv_out_data_59; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_60 = PAR_io_pipe_phv_out_data_60; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_61 = PAR_io_pipe_phv_out_data_61; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_62 = PAR_io_pipe_phv_out_data_62; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_63 = PAR_io_pipe_phv_out_data_63; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_64 = PAR_io_pipe_phv_out_data_64; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_65 = PAR_io_pipe_phv_out_data_65; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_66 = PAR_io_pipe_phv_out_data_66; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_67 = PAR_io_pipe_phv_out_data_67; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_68 = PAR_io_pipe_phv_out_data_68; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_69 = PAR_io_pipe_phv_out_data_69; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_70 = PAR_io_pipe_phv_out_data_70; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_71 = PAR_io_pipe_phv_out_data_71; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_72 = PAR_io_pipe_phv_out_data_72; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_73 = PAR_io_pipe_phv_out_data_73; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_74 = PAR_io_pipe_phv_out_data_74; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_75 = PAR_io_pipe_phv_out_data_75; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_76 = PAR_io_pipe_phv_out_data_76; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_77 = PAR_io_pipe_phv_out_data_77; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_78 = PAR_io_pipe_phv_out_data_78; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_79 = PAR_io_pipe_phv_out_data_79; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_80 = PAR_io_pipe_phv_out_data_80; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_81 = PAR_io_pipe_phv_out_data_81; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_82 = PAR_io_pipe_phv_out_data_82; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_83 = PAR_io_pipe_phv_out_data_83; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_84 = PAR_io_pipe_phv_out_data_84; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_85 = PAR_io_pipe_phv_out_data_85; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_86 = PAR_io_pipe_phv_out_data_86; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_87 = PAR_io_pipe_phv_out_data_87; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_88 = PAR_io_pipe_phv_out_data_88; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_89 = PAR_io_pipe_phv_out_data_89; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_90 = PAR_io_pipe_phv_out_data_90; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_91 = PAR_io_pipe_phv_out_data_91; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_92 = PAR_io_pipe_phv_out_data_92; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_93 = PAR_io_pipe_phv_out_data_93; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_94 = PAR_io_pipe_phv_out_data_94; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_95 = PAR_io_pipe_phv_out_data_95; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_96 = PAR_io_pipe_phv_out_data_96; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_97 = PAR_io_pipe_phv_out_data_97; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_98 = PAR_io_pipe_phv_out_data_98; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_99 = PAR_io_pipe_phv_out_data_99; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_100 = PAR_io_pipe_phv_out_data_100; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_101 = PAR_io_pipe_phv_out_data_101; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_102 = PAR_io_pipe_phv_out_data_102; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_103 = PAR_io_pipe_phv_out_data_103; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_104 = PAR_io_pipe_phv_out_data_104; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_105 = PAR_io_pipe_phv_out_data_105; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_106 = PAR_io_pipe_phv_out_data_106; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_107 = PAR_io_pipe_phv_out_data_107; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_108 = PAR_io_pipe_phv_out_data_108; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_109 = PAR_io_pipe_phv_out_data_109; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_110 = PAR_io_pipe_phv_out_data_110; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_111 = PAR_io_pipe_phv_out_data_111; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_112 = PAR_io_pipe_phv_out_data_112; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_113 = PAR_io_pipe_phv_out_data_113; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_114 = PAR_io_pipe_phv_out_data_114; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_115 = PAR_io_pipe_phv_out_data_115; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_116 = PAR_io_pipe_phv_out_data_116; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_117 = PAR_io_pipe_phv_out_data_117; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_118 = PAR_io_pipe_phv_out_data_118; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_119 = PAR_io_pipe_phv_out_data_119; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_120 = PAR_io_pipe_phv_out_data_120; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_121 = PAR_io_pipe_phv_out_data_121; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_122 = PAR_io_pipe_phv_out_data_122; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_123 = PAR_io_pipe_phv_out_data_123; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_124 = PAR_io_pipe_phv_out_data_124; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_125 = PAR_io_pipe_phv_out_data_125; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_126 = PAR_io_pipe_phv_out_data_126; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_127 = PAR_io_pipe_phv_out_data_127; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_128 = PAR_io_pipe_phv_out_data_128; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_129 = PAR_io_pipe_phv_out_data_129; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_130 = PAR_io_pipe_phv_out_data_130; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_131 = PAR_io_pipe_phv_out_data_131; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_132 = PAR_io_pipe_phv_out_data_132; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_133 = PAR_io_pipe_phv_out_data_133; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_134 = PAR_io_pipe_phv_out_data_134; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_135 = PAR_io_pipe_phv_out_data_135; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_136 = PAR_io_pipe_phv_out_data_136; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_137 = PAR_io_pipe_phv_out_data_137; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_138 = PAR_io_pipe_phv_out_data_138; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_139 = PAR_io_pipe_phv_out_data_139; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_140 = PAR_io_pipe_phv_out_data_140; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_141 = PAR_io_pipe_phv_out_data_141; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_142 = PAR_io_pipe_phv_out_data_142; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_143 = PAR_io_pipe_phv_out_data_143; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_144 = PAR_io_pipe_phv_out_data_144; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_145 = PAR_io_pipe_phv_out_data_145; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_146 = PAR_io_pipe_phv_out_data_146; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_147 = PAR_io_pipe_phv_out_data_147; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_148 = PAR_io_pipe_phv_out_data_148; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_149 = PAR_io_pipe_phv_out_data_149; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_150 = PAR_io_pipe_phv_out_data_150; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_151 = PAR_io_pipe_phv_out_data_151; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_152 = PAR_io_pipe_phv_out_data_152; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_153 = PAR_io_pipe_phv_out_data_153; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_154 = PAR_io_pipe_phv_out_data_154; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_155 = PAR_io_pipe_phv_out_data_155; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_156 = PAR_io_pipe_phv_out_data_156; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_157 = PAR_io_pipe_phv_out_data_157; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_158 = PAR_io_pipe_phv_out_data_158; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_data_159 = PAR_io_pipe_phv_out_data_159; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_next_processor_id = PAR_io_pipe_phv_out_next_processor_id; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_next_config_id = PAR_io_pipe_phv_out_next_config_id; // @[pisa.scala 38:36]
  assign proc_0_io_pipe_phv_in_is_valid_processor = PAR_io_pipe_phv_out_valid; // @[pisa.scala 39:55]
  assign proc_0_io_pipe_phv_in_valid = PAR_io_pipe_phv_out_valid; // @[pisa.scala 38:36]
  assign proc_0_io_mod_mat_mod_en = io_mod_proc_mod_0_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_config_id = io_mod_proc_mod_0_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_0_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_0_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_0_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_0_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_0_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_0_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_0_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_en = io_mod_proc_mod_0_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_0_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_addr = io_mod_proc_mod_0_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_0_io_mod_mat_mod_w_data = io_mod_proc_mod_0_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_en_0 = io_mod_proc_mod_0_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_en_1 = io_mod_proc_mod_0_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_addr = io_mod_proc_mod_0_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_data_0 = io_mod_proc_mod_0_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_0_io_mod_exe_mod_data_1 = io_mod_proc_mod_0_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_1_clock = clock;
  assign proc_1_io_pipe_phv_in_data_0 = proc_0_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_1 = proc_0_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_2 = proc_0_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_3 = proc_0_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_4 = proc_0_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_5 = proc_0_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_6 = proc_0_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_7 = proc_0_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_8 = proc_0_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_9 = proc_0_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_10 = proc_0_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_11 = proc_0_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_12 = proc_0_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_13 = proc_0_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_14 = proc_0_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_15 = proc_0_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_16 = proc_0_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_17 = proc_0_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_18 = proc_0_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_19 = proc_0_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_20 = proc_0_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_21 = proc_0_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_22 = proc_0_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_23 = proc_0_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_24 = proc_0_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_25 = proc_0_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_26 = proc_0_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_27 = proc_0_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_28 = proc_0_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_29 = proc_0_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_30 = proc_0_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_31 = proc_0_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_32 = proc_0_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_33 = proc_0_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_34 = proc_0_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_35 = proc_0_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_36 = proc_0_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_37 = proc_0_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_38 = proc_0_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_39 = proc_0_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_40 = proc_0_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_41 = proc_0_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_42 = proc_0_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_43 = proc_0_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_44 = proc_0_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_45 = proc_0_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_46 = proc_0_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_47 = proc_0_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_48 = proc_0_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_49 = proc_0_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_50 = proc_0_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_51 = proc_0_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_52 = proc_0_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_53 = proc_0_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_54 = proc_0_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_55 = proc_0_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_56 = proc_0_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_57 = proc_0_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_58 = proc_0_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_59 = proc_0_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_60 = proc_0_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_61 = proc_0_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_62 = proc_0_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_63 = proc_0_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_64 = proc_0_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_65 = proc_0_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_66 = proc_0_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_67 = proc_0_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_68 = proc_0_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_69 = proc_0_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_70 = proc_0_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_71 = proc_0_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_72 = proc_0_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_73 = proc_0_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_74 = proc_0_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_75 = proc_0_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_76 = proc_0_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_77 = proc_0_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_78 = proc_0_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_79 = proc_0_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_80 = proc_0_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_81 = proc_0_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_82 = proc_0_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_83 = proc_0_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_84 = proc_0_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_85 = proc_0_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_86 = proc_0_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_87 = proc_0_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_88 = proc_0_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_89 = proc_0_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_90 = proc_0_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_91 = proc_0_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_92 = proc_0_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_93 = proc_0_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_94 = proc_0_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_95 = proc_0_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_96 = proc_0_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_97 = proc_0_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_98 = proc_0_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_99 = proc_0_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_100 = proc_0_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_101 = proc_0_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_102 = proc_0_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_103 = proc_0_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_104 = proc_0_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_105 = proc_0_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_106 = proc_0_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_107 = proc_0_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_108 = proc_0_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_109 = proc_0_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_110 = proc_0_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_111 = proc_0_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_112 = proc_0_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_113 = proc_0_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_114 = proc_0_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_115 = proc_0_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_116 = proc_0_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_117 = proc_0_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_118 = proc_0_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_119 = proc_0_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_120 = proc_0_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_121 = proc_0_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_122 = proc_0_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_123 = proc_0_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_124 = proc_0_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_125 = proc_0_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_126 = proc_0_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_127 = proc_0_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_128 = proc_0_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_129 = proc_0_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_130 = proc_0_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_131 = proc_0_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_132 = proc_0_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_133 = proc_0_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_134 = proc_0_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_135 = proc_0_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_136 = proc_0_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_137 = proc_0_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_138 = proc_0_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_139 = proc_0_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_140 = proc_0_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_141 = proc_0_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_142 = proc_0_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_143 = proc_0_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_144 = proc_0_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_145 = proc_0_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_146 = proc_0_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_147 = proc_0_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_148 = proc_0_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_149 = proc_0_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_150 = proc_0_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_151 = proc_0_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_152 = proc_0_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_153 = proc_0_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_154 = proc_0_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_155 = proc_0_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_156 = proc_0_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_157 = proc_0_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_158 = proc_0_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_data_159 = proc_0_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_next_processor_id = proc_0_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_next_config_id = proc_0_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_1_io_pipe_phv_in_is_valid_processor = 4'h1 == proc_0_io_pipe_phv_out_next_processor_id &
    proc_0_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_1_io_pipe_phv_in_valid = proc_0_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_1_io_mod_mat_mod_en = io_mod_proc_mod_1_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_config_id = io_mod_proc_mod_1_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_1_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_1_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_1_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_1_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_1_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_1_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_1_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_en = io_mod_proc_mod_1_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_1_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_addr = io_mod_proc_mod_1_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_1_io_mod_mat_mod_w_data = io_mod_proc_mod_1_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_en_0 = io_mod_proc_mod_1_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_en_1 = io_mod_proc_mod_1_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_addr = io_mod_proc_mod_1_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_data_0 = io_mod_proc_mod_1_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_1_io_mod_exe_mod_data_1 = io_mod_proc_mod_1_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_2_clock = clock;
  assign proc_2_io_pipe_phv_in_data_0 = proc_1_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_1 = proc_1_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_2 = proc_1_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_3 = proc_1_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_4 = proc_1_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_5 = proc_1_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_6 = proc_1_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_7 = proc_1_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_8 = proc_1_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_9 = proc_1_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_10 = proc_1_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_11 = proc_1_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_12 = proc_1_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_13 = proc_1_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_14 = proc_1_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_15 = proc_1_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_16 = proc_1_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_17 = proc_1_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_18 = proc_1_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_19 = proc_1_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_20 = proc_1_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_21 = proc_1_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_22 = proc_1_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_23 = proc_1_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_24 = proc_1_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_25 = proc_1_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_26 = proc_1_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_27 = proc_1_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_28 = proc_1_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_29 = proc_1_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_30 = proc_1_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_31 = proc_1_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_32 = proc_1_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_33 = proc_1_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_34 = proc_1_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_35 = proc_1_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_36 = proc_1_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_37 = proc_1_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_38 = proc_1_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_39 = proc_1_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_40 = proc_1_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_41 = proc_1_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_42 = proc_1_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_43 = proc_1_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_44 = proc_1_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_45 = proc_1_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_46 = proc_1_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_47 = proc_1_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_48 = proc_1_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_49 = proc_1_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_50 = proc_1_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_51 = proc_1_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_52 = proc_1_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_53 = proc_1_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_54 = proc_1_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_55 = proc_1_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_56 = proc_1_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_57 = proc_1_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_58 = proc_1_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_59 = proc_1_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_60 = proc_1_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_61 = proc_1_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_62 = proc_1_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_63 = proc_1_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_64 = proc_1_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_65 = proc_1_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_66 = proc_1_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_67 = proc_1_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_68 = proc_1_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_69 = proc_1_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_70 = proc_1_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_71 = proc_1_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_72 = proc_1_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_73 = proc_1_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_74 = proc_1_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_75 = proc_1_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_76 = proc_1_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_77 = proc_1_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_78 = proc_1_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_79 = proc_1_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_80 = proc_1_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_81 = proc_1_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_82 = proc_1_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_83 = proc_1_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_84 = proc_1_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_85 = proc_1_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_86 = proc_1_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_87 = proc_1_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_88 = proc_1_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_89 = proc_1_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_90 = proc_1_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_91 = proc_1_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_92 = proc_1_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_93 = proc_1_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_94 = proc_1_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_95 = proc_1_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_96 = proc_1_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_97 = proc_1_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_98 = proc_1_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_99 = proc_1_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_100 = proc_1_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_101 = proc_1_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_102 = proc_1_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_103 = proc_1_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_104 = proc_1_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_105 = proc_1_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_106 = proc_1_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_107 = proc_1_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_108 = proc_1_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_109 = proc_1_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_110 = proc_1_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_111 = proc_1_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_112 = proc_1_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_113 = proc_1_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_114 = proc_1_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_115 = proc_1_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_116 = proc_1_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_117 = proc_1_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_118 = proc_1_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_119 = proc_1_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_120 = proc_1_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_121 = proc_1_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_122 = proc_1_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_123 = proc_1_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_124 = proc_1_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_125 = proc_1_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_126 = proc_1_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_127 = proc_1_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_128 = proc_1_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_129 = proc_1_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_130 = proc_1_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_131 = proc_1_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_132 = proc_1_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_133 = proc_1_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_134 = proc_1_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_135 = proc_1_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_136 = proc_1_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_137 = proc_1_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_138 = proc_1_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_139 = proc_1_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_140 = proc_1_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_141 = proc_1_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_142 = proc_1_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_143 = proc_1_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_144 = proc_1_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_145 = proc_1_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_146 = proc_1_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_147 = proc_1_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_148 = proc_1_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_149 = proc_1_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_150 = proc_1_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_151 = proc_1_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_152 = proc_1_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_153 = proc_1_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_154 = proc_1_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_155 = proc_1_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_156 = proc_1_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_157 = proc_1_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_158 = proc_1_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_data_159 = proc_1_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_next_processor_id = proc_1_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_next_config_id = proc_1_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_2_io_pipe_phv_in_is_valid_processor = 4'h2 == proc_1_io_pipe_phv_out_next_processor_id &
    proc_1_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_2_io_pipe_phv_in_valid = proc_1_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_2_io_mod_mat_mod_en = io_mod_proc_mod_2_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_config_id = io_mod_proc_mod_2_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_2_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_2_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_2_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_2_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_2_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_2_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_2_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_en = io_mod_proc_mod_2_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_2_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_addr = io_mod_proc_mod_2_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_2_io_mod_mat_mod_w_data = io_mod_proc_mod_2_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_en_0 = io_mod_proc_mod_2_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_en_1 = io_mod_proc_mod_2_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_addr = io_mod_proc_mod_2_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_data_0 = io_mod_proc_mod_2_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_2_io_mod_exe_mod_data_1 = io_mod_proc_mod_2_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_3_clock = clock;
  assign proc_3_io_pipe_phv_in_data_0 = proc_2_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_1 = proc_2_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_2 = proc_2_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_3 = proc_2_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_4 = proc_2_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_5 = proc_2_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_6 = proc_2_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_7 = proc_2_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_8 = proc_2_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_9 = proc_2_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_10 = proc_2_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_11 = proc_2_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_12 = proc_2_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_13 = proc_2_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_14 = proc_2_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_15 = proc_2_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_16 = proc_2_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_17 = proc_2_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_18 = proc_2_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_19 = proc_2_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_20 = proc_2_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_21 = proc_2_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_22 = proc_2_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_23 = proc_2_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_24 = proc_2_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_25 = proc_2_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_26 = proc_2_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_27 = proc_2_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_28 = proc_2_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_29 = proc_2_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_30 = proc_2_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_31 = proc_2_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_32 = proc_2_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_33 = proc_2_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_34 = proc_2_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_35 = proc_2_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_36 = proc_2_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_37 = proc_2_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_38 = proc_2_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_39 = proc_2_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_40 = proc_2_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_41 = proc_2_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_42 = proc_2_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_43 = proc_2_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_44 = proc_2_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_45 = proc_2_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_46 = proc_2_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_47 = proc_2_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_48 = proc_2_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_49 = proc_2_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_50 = proc_2_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_51 = proc_2_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_52 = proc_2_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_53 = proc_2_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_54 = proc_2_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_55 = proc_2_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_56 = proc_2_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_57 = proc_2_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_58 = proc_2_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_59 = proc_2_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_60 = proc_2_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_61 = proc_2_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_62 = proc_2_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_63 = proc_2_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_64 = proc_2_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_65 = proc_2_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_66 = proc_2_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_67 = proc_2_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_68 = proc_2_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_69 = proc_2_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_70 = proc_2_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_71 = proc_2_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_72 = proc_2_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_73 = proc_2_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_74 = proc_2_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_75 = proc_2_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_76 = proc_2_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_77 = proc_2_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_78 = proc_2_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_79 = proc_2_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_80 = proc_2_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_81 = proc_2_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_82 = proc_2_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_83 = proc_2_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_84 = proc_2_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_85 = proc_2_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_86 = proc_2_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_87 = proc_2_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_88 = proc_2_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_89 = proc_2_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_90 = proc_2_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_91 = proc_2_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_92 = proc_2_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_93 = proc_2_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_94 = proc_2_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_95 = proc_2_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_96 = proc_2_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_97 = proc_2_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_98 = proc_2_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_99 = proc_2_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_100 = proc_2_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_101 = proc_2_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_102 = proc_2_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_103 = proc_2_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_104 = proc_2_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_105 = proc_2_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_106 = proc_2_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_107 = proc_2_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_108 = proc_2_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_109 = proc_2_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_110 = proc_2_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_111 = proc_2_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_112 = proc_2_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_113 = proc_2_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_114 = proc_2_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_115 = proc_2_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_116 = proc_2_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_117 = proc_2_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_118 = proc_2_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_119 = proc_2_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_120 = proc_2_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_121 = proc_2_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_122 = proc_2_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_123 = proc_2_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_124 = proc_2_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_125 = proc_2_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_126 = proc_2_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_127 = proc_2_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_128 = proc_2_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_129 = proc_2_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_130 = proc_2_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_131 = proc_2_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_132 = proc_2_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_133 = proc_2_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_134 = proc_2_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_135 = proc_2_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_136 = proc_2_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_137 = proc_2_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_138 = proc_2_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_139 = proc_2_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_140 = proc_2_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_141 = proc_2_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_142 = proc_2_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_143 = proc_2_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_144 = proc_2_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_145 = proc_2_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_146 = proc_2_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_147 = proc_2_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_148 = proc_2_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_149 = proc_2_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_150 = proc_2_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_151 = proc_2_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_152 = proc_2_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_153 = proc_2_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_154 = proc_2_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_155 = proc_2_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_156 = proc_2_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_157 = proc_2_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_158 = proc_2_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_data_159 = proc_2_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_next_processor_id = proc_2_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_next_config_id = proc_2_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_3_io_pipe_phv_in_is_valid_processor = 4'h3 == proc_2_io_pipe_phv_out_next_processor_id &
    proc_2_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_3_io_pipe_phv_in_valid = proc_2_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_3_io_mod_mat_mod_en = io_mod_proc_mod_3_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_config_id = io_mod_proc_mod_3_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_3_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_3_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_3_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_3_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_3_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_3_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_3_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_en = io_mod_proc_mod_3_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_3_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_addr = io_mod_proc_mod_3_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_3_io_mod_mat_mod_w_data = io_mod_proc_mod_3_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_en_0 = io_mod_proc_mod_3_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_en_1 = io_mod_proc_mod_3_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_addr = io_mod_proc_mod_3_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_data_0 = io_mod_proc_mod_3_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_3_io_mod_exe_mod_data_1 = io_mod_proc_mod_3_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_4_clock = clock;
  assign proc_4_io_pipe_phv_in_data_0 = proc_3_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_1 = proc_3_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_2 = proc_3_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_3 = proc_3_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_4 = proc_3_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_5 = proc_3_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_6 = proc_3_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_7 = proc_3_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_8 = proc_3_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_9 = proc_3_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_10 = proc_3_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_11 = proc_3_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_12 = proc_3_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_13 = proc_3_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_14 = proc_3_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_15 = proc_3_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_16 = proc_3_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_17 = proc_3_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_18 = proc_3_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_19 = proc_3_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_20 = proc_3_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_21 = proc_3_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_22 = proc_3_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_23 = proc_3_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_24 = proc_3_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_25 = proc_3_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_26 = proc_3_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_27 = proc_3_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_28 = proc_3_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_29 = proc_3_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_30 = proc_3_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_31 = proc_3_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_32 = proc_3_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_33 = proc_3_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_34 = proc_3_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_35 = proc_3_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_36 = proc_3_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_37 = proc_3_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_38 = proc_3_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_39 = proc_3_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_40 = proc_3_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_41 = proc_3_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_42 = proc_3_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_43 = proc_3_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_44 = proc_3_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_45 = proc_3_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_46 = proc_3_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_47 = proc_3_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_48 = proc_3_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_49 = proc_3_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_50 = proc_3_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_51 = proc_3_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_52 = proc_3_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_53 = proc_3_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_54 = proc_3_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_55 = proc_3_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_56 = proc_3_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_57 = proc_3_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_58 = proc_3_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_59 = proc_3_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_60 = proc_3_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_61 = proc_3_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_62 = proc_3_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_63 = proc_3_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_64 = proc_3_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_65 = proc_3_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_66 = proc_3_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_67 = proc_3_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_68 = proc_3_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_69 = proc_3_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_70 = proc_3_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_71 = proc_3_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_72 = proc_3_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_73 = proc_3_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_74 = proc_3_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_75 = proc_3_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_76 = proc_3_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_77 = proc_3_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_78 = proc_3_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_79 = proc_3_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_80 = proc_3_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_81 = proc_3_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_82 = proc_3_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_83 = proc_3_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_84 = proc_3_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_85 = proc_3_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_86 = proc_3_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_87 = proc_3_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_88 = proc_3_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_89 = proc_3_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_90 = proc_3_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_91 = proc_3_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_92 = proc_3_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_93 = proc_3_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_94 = proc_3_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_95 = proc_3_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_96 = proc_3_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_97 = proc_3_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_98 = proc_3_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_99 = proc_3_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_100 = proc_3_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_101 = proc_3_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_102 = proc_3_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_103 = proc_3_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_104 = proc_3_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_105 = proc_3_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_106 = proc_3_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_107 = proc_3_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_108 = proc_3_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_109 = proc_3_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_110 = proc_3_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_111 = proc_3_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_112 = proc_3_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_113 = proc_3_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_114 = proc_3_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_115 = proc_3_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_116 = proc_3_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_117 = proc_3_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_118 = proc_3_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_119 = proc_3_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_120 = proc_3_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_121 = proc_3_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_122 = proc_3_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_123 = proc_3_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_124 = proc_3_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_125 = proc_3_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_126 = proc_3_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_127 = proc_3_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_128 = proc_3_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_129 = proc_3_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_130 = proc_3_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_131 = proc_3_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_132 = proc_3_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_133 = proc_3_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_134 = proc_3_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_135 = proc_3_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_136 = proc_3_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_137 = proc_3_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_138 = proc_3_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_139 = proc_3_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_140 = proc_3_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_141 = proc_3_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_142 = proc_3_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_143 = proc_3_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_144 = proc_3_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_145 = proc_3_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_146 = proc_3_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_147 = proc_3_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_148 = proc_3_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_149 = proc_3_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_150 = proc_3_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_151 = proc_3_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_152 = proc_3_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_153 = proc_3_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_154 = proc_3_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_155 = proc_3_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_156 = proc_3_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_157 = proc_3_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_158 = proc_3_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_data_159 = proc_3_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_next_processor_id = proc_3_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_next_config_id = proc_3_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_4_io_pipe_phv_in_is_valid_processor = 4'h4 == proc_3_io_pipe_phv_out_next_processor_id &
    proc_3_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_4_io_pipe_phv_in_valid = proc_3_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_4_io_mod_mat_mod_en = io_mod_proc_mod_4_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_config_id = io_mod_proc_mod_4_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_4_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_4_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_4_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_4_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_4_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_4_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_4_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_en = io_mod_proc_mod_4_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_4_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_addr = io_mod_proc_mod_4_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_4_io_mod_mat_mod_w_data = io_mod_proc_mod_4_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_en_0 = io_mod_proc_mod_4_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_en_1 = io_mod_proc_mod_4_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_addr = io_mod_proc_mod_4_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_data_0 = io_mod_proc_mod_4_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_4_io_mod_exe_mod_data_1 = io_mod_proc_mod_4_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_5_clock = clock;
  assign proc_5_io_pipe_phv_in_data_0 = proc_4_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_1 = proc_4_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_2 = proc_4_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_3 = proc_4_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_4 = proc_4_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_5 = proc_4_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_6 = proc_4_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_7 = proc_4_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_8 = proc_4_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_9 = proc_4_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_10 = proc_4_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_11 = proc_4_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_12 = proc_4_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_13 = proc_4_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_14 = proc_4_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_15 = proc_4_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_16 = proc_4_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_17 = proc_4_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_18 = proc_4_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_19 = proc_4_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_20 = proc_4_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_21 = proc_4_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_22 = proc_4_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_23 = proc_4_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_24 = proc_4_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_25 = proc_4_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_26 = proc_4_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_27 = proc_4_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_28 = proc_4_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_29 = proc_4_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_30 = proc_4_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_31 = proc_4_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_32 = proc_4_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_33 = proc_4_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_34 = proc_4_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_35 = proc_4_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_36 = proc_4_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_37 = proc_4_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_38 = proc_4_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_39 = proc_4_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_40 = proc_4_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_41 = proc_4_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_42 = proc_4_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_43 = proc_4_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_44 = proc_4_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_45 = proc_4_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_46 = proc_4_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_47 = proc_4_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_48 = proc_4_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_49 = proc_4_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_50 = proc_4_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_51 = proc_4_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_52 = proc_4_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_53 = proc_4_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_54 = proc_4_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_55 = proc_4_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_56 = proc_4_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_57 = proc_4_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_58 = proc_4_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_59 = proc_4_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_60 = proc_4_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_61 = proc_4_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_62 = proc_4_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_63 = proc_4_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_64 = proc_4_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_65 = proc_4_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_66 = proc_4_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_67 = proc_4_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_68 = proc_4_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_69 = proc_4_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_70 = proc_4_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_71 = proc_4_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_72 = proc_4_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_73 = proc_4_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_74 = proc_4_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_75 = proc_4_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_76 = proc_4_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_77 = proc_4_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_78 = proc_4_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_79 = proc_4_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_80 = proc_4_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_81 = proc_4_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_82 = proc_4_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_83 = proc_4_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_84 = proc_4_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_85 = proc_4_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_86 = proc_4_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_87 = proc_4_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_88 = proc_4_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_89 = proc_4_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_90 = proc_4_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_91 = proc_4_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_92 = proc_4_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_93 = proc_4_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_94 = proc_4_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_95 = proc_4_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_96 = proc_4_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_97 = proc_4_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_98 = proc_4_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_99 = proc_4_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_100 = proc_4_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_101 = proc_4_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_102 = proc_4_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_103 = proc_4_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_104 = proc_4_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_105 = proc_4_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_106 = proc_4_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_107 = proc_4_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_108 = proc_4_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_109 = proc_4_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_110 = proc_4_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_111 = proc_4_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_112 = proc_4_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_113 = proc_4_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_114 = proc_4_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_115 = proc_4_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_116 = proc_4_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_117 = proc_4_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_118 = proc_4_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_119 = proc_4_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_120 = proc_4_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_121 = proc_4_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_122 = proc_4_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_123 = proc_4_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_124 = proc_4_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_125 = proc_4_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_126 = proc_4_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_127 = proc_4_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_128 = proc_4_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_129 = proc_4_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_130 = proc_4_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_131 = proc_4_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_132 = proc_4_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_133 = proc_4_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_134 = proc_4_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_135 = proc_4_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_136 = proc_4_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_137 = proc_4_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_138 = proc_4_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_139 = proc_4_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_140 = proc_4_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_141 = proc_4_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_142 = proc_4_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_143 = proc_4_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_144 = proc_4_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_145 = proc_4_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_146 = proc_4_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_147 = proc_4_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_148 = proc_4_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_149 = proc_4_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_150 = proc_4_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_151 = proc_4_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_152 = proc_4_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_153 = proc_4_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_154 = proc_4_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_155 = proc_4_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_156 = proc_4_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_157 = proc_4_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_158 = proc_4_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_data_159 = proc_4_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_next_processor_id = proc_4_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_next_config_id = proc_4_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_5_io_pipe_phv_in_is_valid_processor = 4'h5 == proc_4_io_pipe_phv_out_next_processor_id &
    proc_4_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_5_io_pipe_phv_in_valid = proc_4_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_5_io_mod_mat_mod_en = io_mod_proc_mod_5_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_config_id = io_mod_proc_mod_5_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_5_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_5_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_5_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_5_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_5_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_5_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_5_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_en = io_mod_proc_mod_5_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_5_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_addr = io_mod_proc_mod_5_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_5_io_mod_mat_mod_w_data = io_mod_proc_mod_5_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_en_0 = io_mod_proc_mod_5_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_en_1 = io_mod_proc_mod_5_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_addr = io_mod_proc_mod_5_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_data_0 = io_mod_proc_mod_5_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_5_io_mod_exe_mod_data_1 = io_mod_proc_mod_5_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_6_clock = clock;
  assign proc_6_io_pipe_phv_in_data_0 = proc_5_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_1 = proc_5_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_2 = proc_5_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_3 = proc_5_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_4 = proc_5_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_5 = proc_5_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_6 = proc_5_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_7 = proc_5_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_8 = proc_5_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_9 = proc_5_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_10 = proc_5_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_11 = proc_5_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_12 = proc_5_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_13 = proc_5_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_14 = proc_5_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_15 = proc_5_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_16 = proc_5_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_17 = proc_5_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_18 = proc_5_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_19 = proc_5_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_20 = proc_5_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_21 = proc_5_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_22 = proc_5_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_23 = proc_5_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_24 = proc_5_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_25 = proc_5_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_26 = proc_5_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_27 = proc_5_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_28 = proc_5_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_29 = proc_5_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_30 = proc_5_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_31 = proc_5_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_32 = proc_5_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_33 = proc_5_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_34 = proc_5_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_35 = proc_5_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_36 = proc_5_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_37 = proc_5_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_38 = proc_5_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_39 = proc_5_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_40 = proc_5_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_41 = proc_5_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_42 = proc_5_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_43 = proc_5_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_44 = proc_5_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_45 = proc_5_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_46 = proc_5_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_47 = proc_5_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_48 = proc_5_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_49 = proc_5_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_50 = proc_5_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_51 = proc_5_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_52 = proc_5_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_53 = proc_5_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_54 = proc_5_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_55 = proc_5_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_56 = proc_5_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_57 = proc_5_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_58 = proc_5_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_59 = proc_5_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_60 = proc_5_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_61 = proc_5_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_62 = proc_5_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_63 = proc_5_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_64 = proc_5_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_65 = proc_5_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_66 = proc_5_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_67 = proc_5_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_68 = proc_5_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_69 = proc_5_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_70 = proc_5_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_71 = proc_5_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_72 = proc_5_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_73 = proc_5_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_74 = proc_5_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_75 = proc_5_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_76 = proc_5_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_77 = proc_5_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_78 = proc_5_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_79 = proc_5_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_80 = proc_5_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_81 = proc_5_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_82 = proc_5_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_83 = proc_5_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_84 = proc_5_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_85 = proc_5_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_86 = proc_5_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_87 = proc_5_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_88 = proc_5_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_89 = proc_5_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_90 = proc_5_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_91 = proc_5_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_92 = proc_5_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_93 = proc_5_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_94 = proc_5_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_95 = proc_5_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_96 = proc_5_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_97 = proc_5_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_98 = proc_5_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_99 = proc_5_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_100 = proc_5_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_101 = proc_5_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_102 = proc_5_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_103 = proc_5_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_104 = proc_5_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_105 = proc_5_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_106 = proc_5_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_107 = proc_5_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_108 = proc_5_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_109 = proc_5_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_110 = proc_5_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_111 = proc_5_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_112 = proc_5_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_113 = proc_5_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_114 = proc_5_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_115 = proc_5_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_116 = proc_5_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_117 = proc_5_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_118 = proc_5_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_119 = proc_5_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_120 = proc_5_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_121 = proc_5_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_122 = proc_5_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_123 = proc_5_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_124 = proc_5_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_125 = proc_5_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_126 = proc_5_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_127 = proc_5_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_128 = proc_5_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_129 = proc_5_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_130 = proc_5_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_131 = proc_5_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_132 = proc_5_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_133 = proc_5_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_134 = proc_5_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_135 = proc_5_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_136 = proc_5_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_137 = proc_5_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_138 = proc_5_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_139 = proc_5_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_140 = proc_5_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_141 = proc_5_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_142 = proc_5_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_143 = proc_5_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_144 = proc_5_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_145 = proc_5_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_146 = proc_5_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_147 = proc_5_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_148 = proc_5_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_149 = proc_5_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_150 = proc_5_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_151 = proc_5_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_152 = proc_5_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_153 = proc_5_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_154 = proc_5_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_155 = proc_5_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_156 = proc_5_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_157 = proc_5_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_158 = proc_5_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_data_159 = proc_5_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_next_processor_id = proc_5_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_next_config_id = proc_5_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_6_io_pipe_phv_in_is_valid_processor = 4'h6 == proc_5_io_pipe_phv_out_next_processor_id &
    proc_5_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_6_io_pipe_phv_in_valid = proc_5_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_6_io_mod_mat_mod_en = io_mod_proc_mod_6_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_config_id = io_mod_proc_mod_6_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_6_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_6_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_6_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_6_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_6_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_6_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_6_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_en = io_mod_proc_mod_6_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_6_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_addr = io_mod_proc_mod_6_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_6_io_mod_mat_mod_w_data = io_mod_proc_mod_6_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_en_0 = io_mod_proc_mod_6_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_en_1 = io_mod_proc_mod_6_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_addr = io_mod_proc_mod_6_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_data_0 = io_mod_proc_mod_6_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_6_io_mod_exe_mod_data_1 = io_mod_proc_mod_6_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_7_clock = clock;
  assign proc_7_io_pipe_phv_in_data_0 = proc_6_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_1 = proc_6_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_2 = proc_6_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_3 = proc_6_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_4 = proc_6_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_5 = proc_6_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_6 = proc_6_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_7 = proc_6_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_8 = proc_6_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_9 = proc_6_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_10 = proc_6_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_11 = proc_6_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_12 = proc_6_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_13 = proc_6_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_14 = proc_6_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_15 = proc_6_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_16 = proc_6_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_17 = proc_6_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_18 = proc_6_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_19 = proc_6_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_20 = proc_6_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_21 = proc_6_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_22 = proc_6_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_23 = proc_6_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_24 = proc_6_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_25 = proc_6_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_26 = proc_6_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_27 = proc_6_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_28 = proc_6_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_29 = proc_6_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_30 = proc_6_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_31 = proc_6_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_32 = proc_6_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_33 = proc_6_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_34 = proc_6_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_35 = proc_6_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_36 = proc_6_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_37 = proc_6_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_38 = proc_6_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_39 = proc_6_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_40 = proc_6_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_41 = proc_6_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_42 = proc_6_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_43 = proc_6_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_44 = proc_6_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_45 = proc_6_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_46 = proc_6_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_47 = proc_6_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_48 = proc_6_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_49 = proc_6_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_50 = proc_6_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_51 = proc_6_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_52 = proc_6_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_53 = proc_6_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_54 = proc_6_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_55 = proc_6_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_56 = proc_6_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_57 = proc_6_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_58 = proc_6_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_59 = proc_6_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_60 = proc_6_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_61 = proc_6_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_62 = proc_6_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_63 = proc_6_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_64 = proc_6_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_65 = proc_6_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_66 = proc_6_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_67 = proc_6_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_68 = proc_6_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_69 = proc_6_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_70 = proc_6_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_71 = proc_6_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_72 = proc_6_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_73 = proc_6_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_74 = proc_6_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_75 = proc_6_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_76 = proc_6_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_77 = proc_6_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_78 = proc_6_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_79 = proc_6_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_80 = proc_6_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_81 = proc_6_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_82 = proc_6_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_83 = proc_6_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_84 = proc_6_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_85 = proc_6_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_86 = proc_6_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_87 = proc_6_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_88 = proc_6_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_89 = proc_6_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_90 = proc_6_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_91 = proc_6_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_92 = proc_6_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_93 = proc_6_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_94 = proc_6_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_95 = proc_6_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_96 = proc_6_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_97 = proc_6_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_98 = proc_6_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_99 = proc_6_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_100 = proc_6_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_101 = proc_6_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_102 = proc_6_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_103 = proc_6_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_104 = proc_6_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_105 = proc_6_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_106 = proc_6_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_107 = proc_6_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_108 = proc_6_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_109 = proc_6_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_110 = proc_6_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_111 = proc_6_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_112 = proc_6_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_113 = proc_6_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_114 = proc_6_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_115 = proc_6_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_116 = proc_6_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_117 = proc_6_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_118 = proc_6_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_119 = proc_6_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_120 = proc_6_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_121 = proc_6_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_122 = proc_6_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_123 = proc_6_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_124 = proc_6_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_125 = proc_6_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_126 = proc_6_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_127 = proc_6_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_128 = proc_6_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_129 = proc_6_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_130 = proc_6_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_131 = proc_6_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_132 = proc_6_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_133 = proc_6_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_134 = proc_6_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_135 = proc_6_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_136 = proc_6_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_137 = proc_6_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_138 = proc_6_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_139 = proc_6_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_140 = proc_6_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_141 = proc_6_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_142 = proc_6_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_143 = proc_6_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_144 = proc_6_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_145 = proc_6_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_146 = proc_6_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_147 = proc_6_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_148 = proc_6_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_149 = proc_6_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_150 = proc_6_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_151 = proc_6_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_152 = proc_6_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_153 = proc_6_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_154 = proc_6_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_155 = proc_6_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_156 = proc_6_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_157 = proc_6_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_158 = proc_6_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_data_159 = proc_6_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_next_processor_id = proc_6_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_next_config_id = proc_6_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_7_io_pipe_phv_in_is_valid_processor = 4'h7 == proc_6_io_pipe_phv_out_next_processor_id &
    proc_6_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_7_io_pipe_phv_in_valid = proc_6_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_7_io_mod_mat_mod_en = io_mod_proc_mod_7_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_config_id = io_mod_proc_mod_7_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_7_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_7_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_7_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_7_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_7_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_7_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_7_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_en = io_mod_proc_mod_7_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_7_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_addr = io_mod_proc_mod_7_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_7_io_mod_mat_mod_w_data = io_mod_proc_mod_7_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_en_0 = io_mod_proc_mod_7_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_en_1 = io_mod_proc_mod_7_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_addr = io_mod_proc_mod_7_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_data_0 = io_mod_proc_mod_7_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_7_io_mod_exe_mod_data_1 = io_mod_proc_mod_7_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_8_clock = clock;
  assign proc_8_io_pipe_phv_in_data_0 = proc_7_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_1 = proc_7_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_2 = proc_7_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_3 = proc_7_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_4 = proc_7_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_5 = proc_7_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_6 = proc_7_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_7 = proc_7_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_8 = proc_7_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_9 = proc_7_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_10 = proc_7_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_11 = proc_7_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_12 = proc_7_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_13 = proc_7_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_14 = proc_7_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_15 = proc_7_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_16 = proc_7_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_17 = proc_7_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_18 = proc_7_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_19 = proc_7_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_20 = proc_7_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_21 = proc_7_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_22 = proc_7_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_23 = proc_7_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_24 = proc_7_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_25 = proc_7_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_26 = proc_7_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_27 = proc_7_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_28 = proc_7_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_29 = proc_7_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_30 = proc_7_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_31 = proc_7_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_32 = proc_7_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_33 = proc_7_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_34 = proc_7_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_35 = proc_7_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_36 = proc_7_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_37 = proc_7_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_38 = proc_7_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_39 = proc_7_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_40 = proc_7_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_41 = proc_7_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_42 = proc_7_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_43 = proc_7_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_44 = proc_7_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_45 = proc_7_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_46 = proc_7_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_47 = proc_7_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_48 = proc_7_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_49 = proc_7_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_50 = proc_7_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_51 = proc_7_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_52 = proc_7_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_53 = proc_7_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_54 = proc_7_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_55 = proc_7_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_56 = proc_7_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_57 = proc_7_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_58 = proc_7_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_59 = proc_7_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_60 = proc_7_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_61 = proc_7_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_62 = proc_7_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_63 = proc_7_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_64 = proc_7_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_65 = proc_7_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_66 = proc_7_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_67 = proc_7_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_68 = proc_7_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_69 = proc_7_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_70 = proc_7_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_71 = proc_7_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_72 = proc_7_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_73 = proc_7_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_74 = proc_7_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_75 = proc_7_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_76 = proc_7_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_77 = proc_7_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_78 = proc_7_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_79 = proc_7_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_80 = proc_7_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_81 = proc_7_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_82 = proc_7_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_83 = proc_7_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_84 = proc_7_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_85 = proc_7_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_86 = proc_7_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_87 = proc_7_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_88 = proc_7_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_89 = proc_7_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_90 = proc_7_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_91 = proc_7_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_92 = proc_7_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_93 = proc_7_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_94 = proc_7_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_95 = proc_7_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_96 = proc_7_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_97 = proc_7_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_98 = proc_7_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_99 = proc_7_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_100 = proc_7_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_101 = proc_7_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_102 = proc_7_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_103 = proc_7_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_104 = proc_7_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_105 = proc_7_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_106 = proc_7_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_107 = proc_7_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_108 = proc_7_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_109 = proc_7_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_110 = proc_7_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_111 = proc_7_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_112 = proc_7_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_113 = proc_7_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_114 = proc_7_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_115 = proc_7_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_116 = proc_7_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_117 = proc_7_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_118 = proc_7_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_119 = proc_7_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_120 = proc_7_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_121 = proc_7_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_122 = proc_7_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_123 = proc_7_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_124 = proc_7_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_125 = proc_7_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_126 = proc_7_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_127 = proc_7_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_128 = proc_7_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_129 = proc_7_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_130 = proc_7_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_131 = proc_7_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_132 = proc_7_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_133 = proc_7_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_134 = proc_7_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_135 = proc_7_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_136 = proc_7_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_137 = proc_7_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_138 = proc_7_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_139 = proc_7_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_140 = proc_7_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_141 = proc_7_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_142 = proc_7_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_143 = proc_7_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_144 = proc_7_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_145 = proc_7_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_146 = proc_7_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_147 = proc_7_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_148 = proc_7_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_149 = proc_7_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_150 = proc_7_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_151 = proc_7_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_152 = proc_7_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_153 = proc_7_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_154 = proc_7_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_155 = proc_7_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_156 = proc_7_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_157 = proc_7_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_158 = proc_7_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_data_159 = proc_7_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_next_processor_id = proc_7_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_next_config_id = proc_7_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_8_io_pipe_phv_in_is_valid_processor = 4'h8 == proc_7_io_pipe_phv_out_next_processor_id &
    proc_7_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_8_io_pipe_phv_in_valid = proc_7_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_8_io_mod_mat_mod_en = io_mod_proc_mod_8_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_config_id = io_mod_proc_mod_8_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_8_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_8_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_8_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_8_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_8_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_8_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_8_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_en = io_mod_proc_mod_8_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_8_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_addr = io_mod_proc_mod_8_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_8_io_mod_mat_mod_w_data = io_mod_proc_mod_8_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_en_0 = io_mod_proc_mod_8_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_en_1 = io_mod_proc_mod_8_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_addr = io_mod_proc_mod_8_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_data_0 = io_mod_proc_mod_8_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_8_io_mod_exe_mod_data_1 = io_mod_proc_mod_8_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_9_clock = clock;
  assign proc_9_io_pipe_phv_in_data_0 = proc_8_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_1 = proc_8_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_2 = proc_8_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_3 = proc_8_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_4 = proc_8_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_5 = proc_8_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_6 = proc_8_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_7 = proc_8_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_8 = proc_8_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_9 = proc_8_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_10 = proc_8_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_11 = proc_8_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_12 = proc_8_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_13 = proc_8_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_14 = proc_8_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_15 = proc_8_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_16 = proc_8_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_17 = proc_8_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_18 = proc_8_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_19 = proc_8_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_20 = proc_8_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_21 = proc_8_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_22 = proc_8_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_23 = proc_8_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_24 = proc_8_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_25 = proc_8_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_26 = proc_8_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_27 = proc_8_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_28 = proc_8_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_29 = proc_8_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_30 = proc_8_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_31 = proc_8_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_32 = proc_8_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_33 = proc_8_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_34 = proc_8_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_35 = proc_8_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_36 = proc_8_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_37 = proc_8_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_38 = proc_8_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_39 = proc_8_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_40 = proc_8_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_41 = proc_8_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_42 = proc_8_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_43 = proc_8_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_44 = proc_8_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_45 = proc_8_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_46 = proc_8_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_47 = proc_8_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_48 = proc_8_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_49 = proc_8_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_50 = proc_8_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_51 = proc_8_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_52 = proc_8_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_53 = proc_8_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_54 = proc_8_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_55 = proc_8_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_56 = proc_8_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_57 = proc_8_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_58 = proc_8_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_59 = proc_8_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_60 = proc_8_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_61 = proc_8_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_62 = proc_8_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_63 = proc_8_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_64 = proc_8_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_65 = proc_8_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_66 = proc_8_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_67 = proc_8_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_68 = proc_8_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_69 = proc_8_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_70 = proc_8_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_71 = proc_8_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_72 = proc_8_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_73 = proc_8_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_74 = proc_8_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_75 = proc_8_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_76 = proc_8_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_77 = proc_8_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_78 = proc_8_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_79 = proc_8_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_80 = proc_8_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_81 = proc_8_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_82 = proc_8_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_83 = proc_8_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_84 = proc_8_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_85 = proc_8_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_86 = proc_8_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_87 = proc_8_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_88 = proc_8_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_89 = proc_8_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_90 = proc_8_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_91 = proc_8_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_92 = proc_8_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_93 = proc_8_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_94 = proc_8_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_95 = proc_8_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_96 = proc_8_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_97 = proc_8_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_98 = proc_8_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_99 = proc_8_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_100 = proc_8_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_101 = proc_8_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_102 = proc_8_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_103 = proc_8_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_104 = proc_8_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_105 = proc_8_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_106 = proc_8_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_107 = proc_8_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_108 = proc_8_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_109 = proc_8_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_110 = proc_8_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_111 = proc_8_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_112 = proc_8_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_113 = proc_8_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_114 = proc_8_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_115 = proc_8_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_116 = proc_8_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_117 = proc_8_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_118 = proc_8_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_119 = proc_8_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_120 = proc_8_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_121 = proc_8_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_122 = proc_8_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_123 = proc_8_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_124 = proc_8_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_125 = proc_8_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_126 = proc_8_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_127 = proc_8_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_128 = proc_8_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_129 = proc_8_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_130 = proc_8_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_131 = proc_8_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_132 = proc_8_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_133 = proc_8_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_134 = proc_8_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_135 = proc_8_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_136 = proc_8_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_137 = proc_8_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_138 = proc_8_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_139 = proc_8_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_140 = proc_8_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_141 = proc_8_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_142 = proc_8_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_143 = proc_8_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_144 = proc_8_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_145 = proc_8_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_146 = proc_8_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_147 = proc_8_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_148 = proc_8_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_149 = proc_8_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_150 = proc_8_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_151 = proc_8_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_152 = proc_8_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_153 = proc_8_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_154 = proc_8_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_155 = proc_8_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_156 = proc_8_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_157 = proc_8_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_158 = proc_8_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_data_159 = proc_8_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_next_processor_id = proc_8_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_next_config_id = proc_8_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_9_io_pipe_phv_in_is_valid_processor = 4'h9 == proc_8_io_pipe_phv_out_next_processor_id &
    proc_8_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_9_io_pipe_phv_in_valid = proc_8_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_9_io_mod_mat_mod_en = io_mod_proc_mod_9_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_config_id = io_mod_proc_mod_9_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_9_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_9_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_9_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_9_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_9_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_9_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_9_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_en = io_mod_proc_mod_9_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_9_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_addr = io_mod_proc_mod_9_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_9_io_mod_mat_mod_w_data = io_mod_proc_mod_9_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_en_0 = io_mod_proc_mod_9_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_en_1 = io_mod_proc_mod_9_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_addr = io_mod_proc_mod_9_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_data_0 = io_mod_proc_mod_9_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_9_io_mod_exe_mod_data_1 = io_mod_proc_mod_9_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_10_clock = clock;
  assign proc_10_io_pipe_phv_in_data_0 = proc_9_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_1 = proc_9_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_2 = proc_9_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_3 = proc_9_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_4 = proc_9_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_5 = proc_9_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_6 = proc_9_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_7 = proc_9_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_8 = proc_9_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_9 = proc_9_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_10 = proc_9_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_11 = proc_9_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_12 = proc_9_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_13 = proc_9_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_14 = proc_9_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_15 = proc_9_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_16 = proc_9_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_17 = proc_9_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_18 = proc_9_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_19 = proc_9_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_20 = proc_9_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_21 = proc_9_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_22 = proc_9_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_23 = proc_9_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_24 = proc_9_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_25 = proc_9_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_26 = proc_9_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_27 = proc_9_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_28 = proc_9_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_29 = proc_9_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_30 = proc_9_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_31 = proc_9_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_32 = proc_9_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_33 = proc_9_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_34 = proc_9_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_35 = proc_9_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_36 = proc_9_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_37 = proc_9_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_38 = proc_9_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_39 = proc_9_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_40 = proc_9_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_41 = proc_9_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_42 = proc_9_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_43 = proc_9_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_44 = proc_9_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_45 = proc_9_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_46 = proc_9_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_47 = proc_9_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_48 = proc_9_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_49 = proc_9_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_50 = proc_9_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_51 = proc_9_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_52 = proc_9_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_53 = proc_9_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_54 = proc_9_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_55 = proc_9_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_56 = proc_9_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_57 = proc_9_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_58 = proc_9_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_59 = proc_9_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_60 = proc_9_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_61 = proc_9_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_62 = proc_9_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_63 = proc_9_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_64 = proc_9_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_65 = proc_9_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_66 = proc_9_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_67 = proc_9_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_68 = proc_9_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_69 = proc_9_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_70 = proc_9_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_71 = proc_9_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_72 = proc_9_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_73 = proc_9_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_74 = proc_9_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_75 = proc_9_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_76 = proc_9_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_77 = proc_9_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_78 = proc_9_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_79 = proc_9_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_80 = proc_9_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_81 = proc_9_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_82 = proc_9_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_83 = proc_9_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_84 = proc_9_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_85 = proc_9_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_86 = proc_9_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_87 = proc_9_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_88 = proc_9_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_89 = proc_9_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_90 = proc_9_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_91 = proc_9_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_92 = proc_9_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_93 = proc_9_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_94 = proc_9_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_95 = proc_9_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_96 = proc_9_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_97 = proc_9_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_98 = proc_9_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_99 = proc_9_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_100 = proc_9_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_101 = proc_9_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_102 = proc_9_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_103 = proc_9_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_104 = proc_9_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_105 = proc_9_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_106 = proc_9_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_107 = proc_9_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_108 = proc_9_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_109 = proc_9_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_110 = proc_9_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_111 = proc_9_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_112 = proc_9_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_113 = proc_9_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_114 = proc_9_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_115 = proc_9_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_116 = proc_9_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_117 = proc_9_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_118 = proc_9_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_119 = proc_9_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_120 = proc_9_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_121 = proc_9_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_122 = proc_9_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_123 = proc_9_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_124 = proc_9_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_125 = proc_9_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_126 = proc_9_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_127 = proc_9_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_128 = proc_9_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_129 = proc_9_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_130 = proc_9_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_131 = proc_9_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_132 = proc_9_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_133 = proc_9_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_134 = proc_9_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_135 = proc_9_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_136 = proc_9_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_137 = proc_9_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_138 = proc_9_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_139 = proc_9_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_140 = proc_9_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_141 = proc_9_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_142 = proc_9_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_143 = proc_9_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_144 = proc_9_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_145 = proc_9_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_146 = proc_9_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_147 = proc_9_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_148 = proc_9_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_149 = proc_9_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_150 = proc_9_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_151 = proc_9_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_152 = proc_9_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_153 = proc_9_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_154 = proc_9_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_155 = proc_9_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_156 = proc_9_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_157 = proc_9_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_158 = proc_9_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_data_159 = proc_9_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_next_processor_id = proc_9_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_next_config_id = proc_9_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_10_io_pipe_phv_in_is_valid_processor = 4'ha == proc_9_io_pipe_phv_out_next_processor_id &
    proc_9_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_10_io_pipe_phv_in_valid = proc_9_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_10_io_mod_mat_mod_en = io_mod_proc_mod_10_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_config_id = io_mod_proc_mod_10_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_10_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_10_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_10_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_10_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_10_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_10_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_10_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_en = io_mod_proc_mod_10_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_10_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_addr = io_mod_proc_mod_10_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_10_io_mod_mat_mod_w_data = io_mod_proc_mod_10_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_en_0 = io_mod_proc_mod_10_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_en_1 = io_mod_proc_mod_10_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_addr = io_mod_proc_mod_10_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_data_0 = io_mod_proc_mod_10_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_10_io_mod_exe_mod_data_1 = io_mod_proc_mod_10_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_11_clock = clock;
  assign proc_11_io_pipe_phv_in_data_0 = proc_10_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_1 = proc_10_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_2 = proc_10_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_3 = proc_10_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_4 = proc_10_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_5 = proc_10_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_6 = proc_10_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_7 = proc_10_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_8 = proc_10_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_9 = proc_10_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_10 = proc_10_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_11 = proc_10_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_12 = proc_10_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_13 = proc_10_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_14 = proc_10_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_15 = proc_10_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_16 = proc_10_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_17 = proc_10_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_18 = proc_10_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_19 = proc_10_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_20 = proc_10_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_21 = proc_10_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_22 = proc_10_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_23 = proc_10_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_24 = proc_10_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_25 = proc_10_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_26 = proc_10_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_27 = proc_10_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_28 = proc_10_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_29 = proc_10_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_30 = proc_10_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_31 = proc_10_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_32 = proc_10_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_33 = proc_10_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_34 = proc_10_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_35 = proc_10_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_36 = proc_10_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_37 = proc_10_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_38 = proc_10_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_39 = proc_10_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_40 = proc_10_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_41 = proc_10_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_42 = proc_10_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_43 = proc_10_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_44 = proc_10_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_45 = proc_10_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_46 = proc_10_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_47 = proc_10_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_48 = proc_10_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_49 = proc_10_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_50 = proc_10_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_51 = proc_10_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_52 = proc_10_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_53 = proc_10_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_54 = proc_10_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_55 = proc_10_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_56 = proc_10_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_57 = proc_10_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_58 = proc_10_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_59 = proc_10_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_60 = proc_10_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_61 = proc_10_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_62 = proc_10_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_63 = proc_10_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_64 = proc_10_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_65 = proc_10_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_66 = proc_10_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_67 = proc_10_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_68 = proc_10_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_69 = proc_10_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_70 = proc_10_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_71 = proc_10_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_72 = proc_10_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_73 = proc_10_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_74 = proc_10_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_75 = proc_10_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_76 = proc_10_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_77 = proc_10_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_78 = proc_10_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_79 = proc_10_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_80 = proc_10_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_81 = proc_10_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_82 = proc_10_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_83 = proc_10_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_84 = proc_10_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_85 = proc_10_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_86 = proc_10_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_87 = proc_10_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_88 = proc_10_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_89 = proc_10_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_90 = proc_10_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_91 = proc_10_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_92 = proc_10_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_93 = proc_10_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_94 = proc_10_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_95 = proc_10_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_96 = proc_10_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_97 = proc_10_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_98 = proc_10_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_99 = proc_10_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_100 = proc_10_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_101 = proc_10_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_102 = proc_10_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_103 = proc_10_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_104 = proc_10_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_105 = proc_10_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_106 = proc_10_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_107 = proc_10_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_108 = proc_10_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_109 = proc_10_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_110 = proc_10_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_111 = proc_10_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_112 = proc_10_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_113 = proc_10_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_114 = proc_10_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_115 = proc_10_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_116 = proc_10_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_117 = proc_10_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_118 = proc_10_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_119 = proc_10_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_120 = proc_10_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_121 = proc_10_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_122 = proc_10_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_123 = proc_10_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_124 = proc_10_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_125 = proc_10_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_126 = proc_10_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_127 = proc_10_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_128 = proc_10_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_129 = proc_10_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_130 = proc_10_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_131 = proc_10_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_132 = proc_10_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_133 = proc_10_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_134 = proc_10_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_135 = proc_10_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_136 = proc_10_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_137 = proc_10_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_138 = proc_10_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_139 = proc_10_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_140 = proc_10_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_141 = proc_10_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_142 = proc_10_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_143 = proc_10_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_144 = proc_10_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_145 = proc_10_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_146 = proc_10_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_147 = proc_10_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_148 = proc_10_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_149 = proc_10_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_150 = proc_10_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_151 = proc_10_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_152 = proc_10_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_153 = proc_10_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_154 = proc_10_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_155 = proc_10_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_156 = proc_10_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_157 = proc_10_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_158 = proc_10_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_data_159 = proc_10_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_next_processor_id = proc_10_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_next_config_id = proc_10_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_11_io_pipe_phv_in_is_valid_processor = 4'hb == proc_10_io_pipe_phv_out_next_processor_id &
    proc_10_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_11_io_pipe_phv_in_valid = proc_10_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_11_io_mod_mat_mod_en = io_mod_proc_mod_11_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_config_id = io_mod_proc_mod_11_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_11_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_11_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_11_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_11_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_11_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_11_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_11_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_en = io_mod_proc_mod_11_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_11_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_addr = io_mod_proc_mod_11_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_11_io_mod_mat_mod_w_data = io_mod_proc_mod_11_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_en_0 = io_mod_proc_mod_11_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_en_1 = io_mod_proc_mod_11_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_addr = io_mod_proc_mod_11_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_data_0 = io_mod_proc_mod_11_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_11_io_mod_exe_mod_data_1 = io_mod_proc_mod_11_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_12_clock = clock;
  assign proc_12_io_pipe_phv_in_data_0 = proc_11_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_1 = proc_11_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_2 = proc_11_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_3 = proc_11_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_4 = proc_11_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_5 = proc_11_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_6 = proc_11_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_7 = proc_11_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_8 = proc_11_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_9 = proc_11_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_10 = proc_11_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_11 = proc_11_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_12 = proc_11_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_13 = proc_11_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_14 = proc_11_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_15 = proc_11_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_16 = proc_11_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_17 = proc_11_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_18 = proc_11_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_19 = proc_11_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_20 = proc_11_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_21 = proc_11_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_22 = proc_11_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_23 = proc_11_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_24 = proc_11_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_25 = proc_11_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_26 = proc_11_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_27 = proc_11_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_28 = proc_11_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_29 = proc_11_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_30 = proc_11_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_31 = proc_11_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_32 = proc_11_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_33 = proc_11_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_34 = proc_11_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_35 = proc_11_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_36 = proc_11_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_37 = proc_11_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_38 = proc_11_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_39 = proc_11_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_40 = proc_11_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_41 = proc_11_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_42 = proc_11_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_43 = proc_11_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_44 = proc_11_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_45 = proc_11_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_46 = proc_11_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_47 = proc_11_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_48 = proc_11_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_49 = proc_11_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_50 = proc_11_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_51 = proc_11_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_52 = proc_11_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_53 = proc_11_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_54 = proc_11_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_55 = proc_11_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_56 = proc_11_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_57 = proc_11_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_58 = proc_11_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_59 = proc_11_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_60 = proc_11_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_61 = proc_11_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_62 = proc_11_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_63 = proc_11_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_64 = proc_11_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_65 = proc_11_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_66 = proc_11_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_67 = proc_11_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_68 = proc_11_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_69 = proc_11_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_70 = proc_11_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_71 = proc_11_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_72 = proc_11_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_73 = proc_11_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_74 = proc_11_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_75 = proc_11_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_76 = proc_11_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_77 = proc_11_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_78 = proc_11_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_79 = proc_11_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_80 = proc_11_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_81 = proc_11_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_82 = proc_11_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_83 = proc_11_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_84 = proc_11_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_85 = proc_11_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_86 = proc_11_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_87 = proc_11_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_88 = proc_11_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_89 = proc_11_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_90 = proc_11_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_91 = proc_11_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_92 = proc_11_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_93 = proc_11_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_94 = proc_11_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_95 = proc_11_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_96 = proc_11_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_97 = proc_11_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_98 = proc_11_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_99 = proc_11_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_100 = proc_11_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_101 = proc_11_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_102 = proc_11_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_103 = proc_11_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_104 = proc_11_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_105 = proc_11_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_106 = proc_11_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_107 = proc_11_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_108 = proc_11_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_109 = proc_11_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_110 = proc_11_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_111 = proc_11_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_112 = proc_11_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_113 = proc_11_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_114 = proc_11_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_115 = proc_11_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_116 = proc_11_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_117 = proc_11_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_118 = proc_11_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_119 = proc_11_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_120 = proc_11_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_121 = proc_11_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_122 = proc_11_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_123 = proc_11_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_124 = proc_11_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_125 = proc_11_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_126 = proc_11_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_127 = proc_11_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_128 = proc_11_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_129 = proc_11_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_130 = proc_11_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_131 = proc_11_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_132 = proc_11_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_133 = proc_11_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_134 = proc_11_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_135 = proc_11_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_136 = proc_11_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_137 = proc_11_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_138 = proc_11_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_139 = proc_11_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_140 = proc_11_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_141 = proc_11_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_142 = proc_11_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_143 = proc_11_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_144 = proc_11_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_145 = proc_11_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_146 = proc_11_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_147 = proc_11_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_148 = proc_11_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_149 = proc_11_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_150 = proc_11_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_151 = proc_11_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_152 = proc_11_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_153 = proc_11_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_154 = proc_11_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_155 = proc_11_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_156 = proc_11_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_157 = proc_11_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_158 = proc_11_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_data_159 = proc_11_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_next_processor_id = proc_11_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_next_config_id = proc_11_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_12_io_pipe_phv_in_is_valid_processor = 4'hc == proc_11_io_pipe_phv_out_next_processor_id &
    proc_11_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_12_io_pipe_phv_in_valid = proc_11_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_12_io_mod_mat_mod_en = io_mod_proc_mod_12_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_config_id = io_mod_proc_mod_12_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_12_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_12_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_12_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_12_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_12_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_12_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_12_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_12_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_12_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_12_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_12_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_12_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_12_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_w_en = io_mod_proc_mod_12_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_12_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_w_addr = io_mod_proc_mod_12_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_12_io_mod_mat_mod_w_data = io_mod_proc_mod_12_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_12_io_mod_exe_mod_en_0 = io_mod_proc_mod_12_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_12_io_mod_exe_mod_en_1 = io_mod_proc_mod_12_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_12_io_mod_exe_mod_addr = io_mod_proc_mod_12_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_12_io_mod_exe_mod_data_0 = io_mod_proc_mod_12_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_12_io_mod_exe_mod_data_1 = io_mod_proc_mod_12_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_13_clock = clock;
  assign proc_13_io_pipe_phv_in_data_0 = proc_12_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_1 = proc_12_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_2 = proc_12_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_3 = proc_12_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_4 = proc_12_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_5 = proc_12_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_6 = proc_12_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_7 = proc_12_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_8 = proc_12_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_9 = proc_12_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_10 = proc_12_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_11 = proc_12_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_12 = proc_12_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_13 = proc_12_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_14 = proc_12_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_15 = proc_12_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_16 = proc_12_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_17 = proc_12_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_18 = proc_12_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_19 = proc_12_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_20 = proc_12_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_21 = proc_12_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_22 = proc_12_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_23 = proc_12_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_24 = proc_12_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_25 = proc_12_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_26 = proc_12_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_27 = proc_12_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_28 = proc_12_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_29 = proc_12_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_30 = proc_12_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_31 = proc_12_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_32 = proc_12_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_33 = proc_12_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_34 = proc_12_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_35 = proc_12_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_36 = proc_12_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_37 = proc_12_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_38 = proc_12_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_39 = proc_12_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_40 = proc_12_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_41 = proc_12_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_42 = proc_12_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_43 = proc_12_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_44 = proc_12_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_45 = proc_12_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_46 = proc_12_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_47 = proc_12_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_48 = proc_12_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_49 = proc_12_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_50 = proc_12_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_51 = proc_12_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_52 = proc_12_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_53 = proc_12_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_54 = proc_12_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_55 = proc_12_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_56 = proc_12_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_57 = proc_12_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_58 = proc_12_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_59 = proc_12_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_60 = proc_12_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_61 = proc_12_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_62 = proc_12_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_63 = proc_12_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_64 = proc_12_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_65 = proc_12_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_66 = proc_12_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_67 = proc_12_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_68 = proc_12_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_69 = proc_12_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_70 = proc_12_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_71 = proc_12_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_72 = proc_12_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_73 = proc_12_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_74 = proc_12_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_75 = proc_12_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_76 = proc_12_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_77 = proc_12_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_78 = proc_12_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_79 = proc_12_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_80 = proc_12_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_81 = proc_12_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_82 = proc_12_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_83 = proc_12_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_84 = proc_12_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_85 = proc_12_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_86 = proc_12_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_87 = proc_12_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_88 = proc_12_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_89 = proc_12_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_90 = proc_12_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_91 = proc_12_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_92 = proc_12_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_93 = proc_12_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_94 = proc_12_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_95 = proc_12_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_96 = proc_12_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_97 = proc_12_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_98 = proc_12_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_99 = proc_12_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_100 = proc_12_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_101 = proc_12_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_102 = proc_12_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_103 = proc_12_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_104 = proc_12_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_105 = proc_12_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_106 = proc_12_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_107 = proc_12_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_108 = proc_12_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_109 = proc_12_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_110 = proc_12_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_111 = proc_12_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_112 = proc_12_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_113 = proc_12_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_114 = proc_12_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_115 = proc_12_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_116 = proc_12_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_117 = proc_12_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_118 = proc_12_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_119 = proc_12_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_120 = proc_12_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_121 = proc_12_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_122 = proc_12_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_123 = proc_12_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_124 = proc_12_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_125 = proc_12_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_126 = proc_12_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_127 = proc_12_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_128 = proc_12_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_129 = proc_12_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_130 = proc_12_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_131 = proc_12_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_132 = proc_12_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_133 = proc_12_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_134 = proc_12_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_135 = proc_12_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_136 = proc_12_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_137 = proc_12_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_138 = proc_12_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_139 = proc_12_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_140 = proc_12_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_141 = proc_12_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_142 = proc_12_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_143 = proc_12_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_144 = proc_12_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_145 = proc_12_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_146 = proc_12_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_147 = proc_12_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_148 = proc_12_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_149 = proc_12_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_150 = proc_12_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_151 = proc_12_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_152 = proc_12_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_153 = proc_12_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_154 = proc_12_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_155 = proc_12_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_156 = proc_12_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_157 = proc_12_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_158 = proc_12_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_data_159 = proc_12_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_next_processor_id = proc_12_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_next_config_id = proc_12_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_13_io_pipe_phv_in_is_valid_processor = 4'hd == proc_12_io_pipe_phv_out_next_processor_id &
    proc_12_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_13_io_pipe_phv_in_valid = proc_12_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_13_io_mod_mat_mod_en = io_mod_proc_mod_13_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_config_id = io_mod_proc_mod_13_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_13_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_13_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_13_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_13_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_13_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_13_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_13_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_13_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_13_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_13_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_13_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_13_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_13_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_w_en = io_mod_proc_mod_13_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_13_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_w_addr = io_mod_proc_mod_13_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_13_io_mod_mat_mod_w_data = io_mod_proc_mod_13_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_13_io_mod_exe_mod_en_0 = io_mod_proc_mod_13_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_13_io_mod_exe_mod_en_1 = io_mod_proc_mod_13_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_13_io_mod_exe_mod_addr = io_mod_proc_mod_13_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_13_io_mod_exe_mod_data_0 = io_mod_proc_mod_13_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_13_io_mod_exe_mod_data_1 = io_mod_proc_mod_13_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_14_clock = clock;
  assign proc_14_io_pipe_phv_in_data_0 = proc_13_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_1 = proc_13_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_2 = proc_13_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_3 = proc_13_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_4 = proc_13_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_5 = proc_13_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_6 = proc_13_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_7 = proc_13_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_8 = proc_13_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_9 = proc_13_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_10 = proc_13_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_11 = proc_13_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_12 = proc_13_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_13 = proc_13_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_14 = proc_13_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_15 = proc_13_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_16 = proc_13_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_17 = proc_13_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_18 = proc_13_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_19 = proc_13_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_20 = proc_13_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_21 = proc_13_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_22 = proc_13_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_23 = proc_13_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_24 = proc_13_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_25 = proc_13_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_26 = proc_13_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_27 = proc_13_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_28 = proc_13_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_29 = proc_13_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_30 = proc_13_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_31 = proc_13_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_32 = proc_13_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_33 = proc_13_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_34 = proc_13_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_35 = proc_13_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_36 = proc_13_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_37 = proc_13_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_38 = proc_13_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_39 = proc_13_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_40 = proc_13_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_41 = proc_13_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_42 = proc_13_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_43 = proc_13_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_44 = proc_13_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_45 = proc_13_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_46 = proc_13_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_47 = proc_13_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_48 = proc_13_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_49 = proc_13_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_50 = proc_13_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_51 = proc_13_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_52 = proc_13_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_53 = proc_13_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_54 = proc_13_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_55 = proc_13_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_56 = proc_13_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_57 = proc_13_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_58 = proc_13_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_59 = proc_13_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_60 = proc_13_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_61 = proc_13_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_62 = proc_13_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_63 = proc_13_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_64 = proc_13_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_65 = proc_13_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_66 = proc_13_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_67 = proc_13_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_68 = proc_13_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_69 = proc_13_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_70 = proc_13_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_71 = proc_13_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_72 = proc_13_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_73 = proc_13_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_74 = proc_13_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_75 = proc_13_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_76 = proc_13_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_77 = proc_13_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_78 = proc_13_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_79 = proc_13_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_80 = proc_13_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_81 = proc_13_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_82 = proc_13_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_83 = proc_13_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_84 = proc_13_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_85 = proc_13_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_86 = proc_13_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_87 = proc_13_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_88 = proc_13_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_89 = proc_13_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_90 = proc_13_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_91 = proc_13_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_92 = proc_13_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_93 = proc_13_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_94 = proc_13_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_95 = proc_13_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_96 = proc_13_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_97 = proc_13_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_98 = proc_13_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_99 = proc_13_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_100 = proc_13_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_101 = proc_13_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_102 = proc_13_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_103 = proc_13_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_104 = proc_13_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_105 = proc_13_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_106 = proc_13_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_107 = proc_13_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_108 = proc_13_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_109 = proc_13_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_110 = proc_13_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_111 = proc_13_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_112 = proc_13_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_113 = proc_13_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_114 = proc_13_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_115 = proc_13_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_116 = proc_13_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_117 = proc_13_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_118 = proc_13_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_119 = proc_13_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_120 = proc_13_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_121 = proc_13_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_122 = proc_13_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_123 = proc_13_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_124 = proc_13_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_125 = proc_13_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_126 = proc_13_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_127 = proc_13_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_128 = proc_13_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_129 = proc_13_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_130 = proc_13_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_131 = proc_13_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_132 = proc_13_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_133 = proc_13_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_134 = proc_13_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_135 = proc_13_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_136 = proc_13_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_137 = proc_13_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_138 = proc_13_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_139 = proc_13_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_140 = proc_13_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_141 = proc_13_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_142 = proc_13_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_143 = proc_13_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_144 = proc_13_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_145 = proc_13_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_146 = proc_13_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_147 = proc_13_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_148 = proc_13_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_149 = proc_13_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_150 = proc_13_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_151 = proc_13_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_152 = proc_13_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_153 = proc_13_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_154 = proc_13_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_155 = proc_13_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_156 = proc_13_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_157 = proc_13_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_158 = proc_13_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_data_159 = proc_13_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_next_processor_id = proc_13_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_next_config_id = proc_13_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_14_io_pipe_phv_in_is_valid_processor = 4'he == proc_13_io_pipe_phv_out_next_processor_id &
    proc_13_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_14_io_pipe_phv_in_valid = proc_13_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_14_io_mod_mat_mod_en = io_mod_proc_mod_14_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_config_id = io_mod_proc_mod_14_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_14_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_14_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_14_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_14_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_14_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_14_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_14_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_14_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_14_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_14_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_14_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_14_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_14_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_w_en = io_mod_proc_mod_14_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_14_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_w_addr = io_mod_proc_mod_14_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_14_io_mod_mat_mod_w_data = io_mod_proc_mod_14_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_14_io_mod_exe_mod_en_0 = io_mod_proc_mod_14_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_14_io_mod_exe_mod_en_1 = io_mod_proc_mod_14_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_14_io_mod_exe_mod_addr = io_mod_proc_mod_14_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_14_io_mod_exe_mod_data_0 = io_mod_proc_mod_14_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_14_io_mod_exe_mod_data_1 = io_mod_proc_mod_14_exe_mod_data_1; // @[pisa.scala 29:20]
  assign proc_15_clock = clock;
  assign proc_15_io_pipe_phv_in_data_0 = proc_14_io_pipe_phv_out_data_0; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_1 = proc_14_io_pipe_phv_out_data_1; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_2 = proc_14_io_pipe_phv_out_data_2; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_3 = proc_14_io_pipe_phv_out_data_3; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_4 = proc_14_io_pipe_phv_out_data_4; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_5 = proc_14_io_pipe_phv_out_data_5; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_6 = proc_14_io_pipe_phv_out_data_6; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_7 = proc_14_io_pipe_phv_out_data_7; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_8 = proc_14_io_pipe_phv_out_data_8; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_9 = proc_14_io_pipe_phv_out_data_9; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_10 = proc_14_io_pipe_phv_out_data_10; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_11 = proc_14_io_pipe_phv_out_data_11; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_12 = proc_14_io_pipe_phv_out_data_12; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_13 = proc_14_io_pipe_phv_out_data_13; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_14 = proc_14_io_pipe_phv_out_data_14; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_15 = proc_14_io_pipe_phv_out_data_15; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_16 = proc_14_io_pipe_phv_out_data_16; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_17 = proc_14_io_pipe_phv_out_data_17; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_18 = proc_14_io_pipe_phv_out_data_18; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_19 = proc_14_io_pipe_phv_out_data_19; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_20 = proc_14_io_pipe_phv_out_data_20; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_21 = proc_14_io_pipe_phv_out_data_21; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_22 = proc_14_io_pipe_phv_out_data_22; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_23 = proc_14_io_pipe_phv_out_data_23; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_24 = proc_14_io_pipe_phv_out_data_24; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_25 = proc_14_io_pipe_phv_out_data_25; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_26 = proc_14_io_pipe_phv_out_data_26; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_27 = proc_14_io_pipe_phv_out_data_27; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_28 = proc_14_io_pipe_phv_out_data_28; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_29 = proc_14_io_pipe_phv_out_data_29; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_30 = proc_14_io_pipe_phv_out_data_30; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_31 = proc_14_io_pipe_phv_out_data_31; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_32 = proc_14_io_pipe_phv_out_data_32; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_33 = proc_14_io_pipe_phv_out_data_33; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_34 = proc_14_io_pipe_phv_out_data_34; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_35 = proc_14_io_pipe_phv_out_data_35; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_36 = proc_14_io_pipe_phv_out_data_36; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_37 = proc_14_io_pipe_phv_out_data_37; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_38 = proc_14_io_pipe_phv_out_data_38; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_39 = proc_14_io_pipe_phv_out_data_39; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_40 = proc_14_io_pipe_phv_out_data_40; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_41 = proc_14_io_pipe_phv_out_data_41; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_42 = proc_14_io_pipe_phv_out_data_42; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_43 = proc_14_io_pipe_phv_out_data_43; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_44 = proc_14_io_pipe_phv_out_data_44; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_45 = proc_14_io_pipe_phv_out_data_45; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_46 = proc_14_io_pipe_phv_out_data_46; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_47 = proc_14_io_pipe_phv_out_data_47; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_48 = proc_14_io_pipe_phv_out_data_48; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_49 = proc_14_io_pipe_phv_out_data_49; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_50 = proc_14_io_pipe_phv_out_data_50; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_51 = proc_14_io_pipe_phv_out_data_51; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_52 = proc_14_io_pipe_phv_out_data_52; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_53 = proc_14_io_pipe_phv_out_data_53; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_54 = proc_14_io_pipe_phv_out_data_54; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_55 = proc_14_io_pipe_phv_out_data_55; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_56 = proc_14_io_pipe_phv_out_data_56; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_57 = proc_14_io_pipe_phv_out_data_57; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_58 = proc_14_io_pipe_phv_out_data_58; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_59 = proc_14_io_pipe_phv_out_data_59; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_60 = proc_14_io_pipe_phv_out_data_60; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_61 = proc_14_io_pipe_phv_out_data_61; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_62 = proc_14_io_pipe_phv_out_data_62; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_63 = proc_14_io_pipe_phv_out_data_63; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_64 = proc_14_io_pipe_phv_out_data_64; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_65 = proc_14_io_pipe_phv_out_data_65; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_66 = proc_14_io_pipe_phv_out_data_66; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_67 = proc_14_io_pipe_phv_out_data_67; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_68 = proc_14_io_pipe_phv_out_data_68; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_69 = proc_14_io_pipe_phv_out_data_69; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_70 = proc_14_io_pipe_phv_out_data_70; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_71 = proc_14_io_pipe_phv_out_data_71; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_72 = proc_14_io_pipe_phv_out_data_72; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_73 = proc_14_io_pipe_phv_out_data_73; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_74 = proc_14_io_pipe_phv_out_data_74; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_75 = proc_14_io_pipe_phv_out_data_75; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_76 = proc_14_io_pipe_phv_out_data_76; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_77 = proc_14_io_pipe_phv_out_data_77; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_78 = proc_14_io_pipe_phv_out_data_78; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_79 = proc_14_io_pipe_phv_out_data_79; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_80 = proc_14_io_pipe_phv_out_data_80; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_81 = proc_14_io_pipe_phv_out_data_81; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_82 = proc_14_io_pipe_phv_out_data_82; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_83 = proc_14_io_pipe_phv_out_data_83; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_84 = proc_14_io_pipe_phv_out_data_84; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_85 = proc_14_io_pipe_phv_out_data_85; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_86 = proc_14_io_pipe_phv_out_data_86; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_87 = proc_14_io_pipe_phv_out_data_87; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_88 = proc_14_io_pipe_phv_out_data_88; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_89 = proc_14_io_pipe_phv_out_data_89; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_90 = proc_14_io_pipe_phv_out_data_90; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_91 = proc_14_io_pipe_phv_out_data_91; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_92 = proc_14_io_pipe_phv_out_data_92; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_93 = proc_14_io_pipe_phv_out_data_93; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_94 = proc_14_io_pipe_phv_out_data_94; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_95 = proc_14_io_pipe_phv_out_data_95; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_96 = proc_14_io_pipe_phv_out_data_96; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_97 = proc_14_io_pipe_phv_out_data_97; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_98 = proc_14_io_pipe_phv_out_data_98; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_99 = proc_14_io_pipe_phv_out_data_99; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_100 = proc_14_io_pipe_phv_out_data_100; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_101 = proc_14_io_pipe_phv_out_data_101; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_102 = proc_14_io_pipe_phv_out_data_102; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_103 = proc_14_io_pipe_phv_out_data_103; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_104 = proc_14_io_pipe_phv_out_data_104; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_105 = proc_14_io_pipe_phv_out_data_105; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_106 = proc_14_io_pipe_phv_out_data_106; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_107 = proc_14_io_pipe_phv_out_data_107; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_108 = proc_14_io_pipe_phv_out_data_108; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_109 = proc_14_io_pipe_phv_out_data_109; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_110 = proc_14_io_pipe_phv_out_data_110; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_111 = proc_14_io_pipe_phv_out_data_111; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_112 = proc_14_io_pipe_phv_out_data_112; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_113 = proc_14_io_pipe_phv_out_data_113; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_114 = proc_14_io_pipe_phv_out_data_114; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_115 = proc_14_io_pipe_phv_out_data_115; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_116 = proc_14_io_pipe_phv_out_data_116; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_117 = proc_14_io_pipe_phv_out_data_117; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_118 = proc_14_io_pipe_phv_out_data_118; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_119 = proc_14_io_pipe_phv_out_data_119; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_120 = proc_14_io_pipe_phv_out_data_120; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_121 = proc_14_io_pipe_phv_out_data_121; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_122 = proc_14_io_pipe_phv_out_data_122; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_123 = proc_14_io_pipe_phv_out_data_123; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_124 = proc_14_io_pipe_phv_out_data_124; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_125 = proc_14_io_pipe_phv_out_data_125; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_126 = proc_14_io_pipe_phv_out_data_126; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_127 = proc_14_io_pipe_phv_out_data_127; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_128 = proc_14_io_pipe_phv_out_data_128; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_129 = proc_14_io_pipe_phv_out_data_129; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_130 = proc_14_io_pipe_phv_out_data_130; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_131 = proc_14_io_pipe_phv_out_data_131; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_132 = proc_14_io_pipe_phv_out_data_132; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_133 = proc_14_io_pipe_phv_out_data_133; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_134 = proc_14_io_pipe_phv_out_data_134; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_135 = proc_14_io_pipe_phv_out_data_135; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_136 = proc_14_io_pipe_phv_out_data_136; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_137 = proc_14_io_pipe_phv_out_data_137; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_138 = proc_14_io_pipe_phv_out_data_138; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_139 = proc_14_io_pipe_phv_out_data_139; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_140 = proc_14_io_pipe_phv_out_data_140; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_141 = proc_14_io_pipe_phv_out_data_141; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_142 = proc_14_io_pipe_phv_out_data_142; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_143 = proc_14_io_pipe_phv_out_data_143; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_144 = proc_14_io_pipe_phv_out_data_144; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_145 = proc_14_io_pipe_phv_out_data_145; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_146 = proc_14_io_pipe_phv_out_data_146; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_147 = proc_14_io_pipe_phv_out_data_147; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_148 = proc_14_io_pipe_phv_out_data_148; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_149 = proc_14_io_pipe_phv_out_data_149; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_150 = proc_14_io_pipe_phv_out_data_150; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_151 = proc_14_io_pipe_phv_out_data_151; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_152 = proc_14_io_pipe_phv_out_data_152; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_153 = proc_14_io_pipe_phv_out_data_153; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_154 = proc_14_io_pipe_phv_out_data_154; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_155 = proc_14_io_pipe_phv_out_data_155; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_156 = proc_14_io_pipe_phv_out_data_156; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_157 = proc_14_io_pipe_phv_out_data_157; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_158 = proc_14_io_pipe_phv_out_data_158; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_data_159 = proc_14_io_pipe_phv_out_data_159; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_next_processor_id = proc_14_io_pipe_phv_out_next_processor_id; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_next_config_id = proc_14_io_pipe_phv_out_next_config_id; // @[pisa.scala 35:36]
  assign proc_15_io_pipe_phv_in_is_valid_processor = 4'hf == proc_14_io_pipe_phv_out_next_processor_id &
    proc_14_io_pipe_phv_out_valid; // @[pisa.scala 36:110]
  assign proc_15_io_pipe_phv_in_valid = proc_14_io_pipe_phv_out_valid; // @[pisa.scala 35:36]
  assign proc_15_io_mod_mat_mod_en = io_mod_proc_mod_15_mat_mod_en; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_config_id = io_mod_proc_mod_15_mat_mod_config_id; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_en = io_mod_proc_mod_15_mat_mod_key_mod_en; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_index = io_mod_proc_mod_15_mat_mod_key_mod_group_index; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_config = io_mod_proc_mod_15_mat_mod_key_mod_group_config; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_mask_0 = io_mod_proc_mod_15_mat_mod_key_mod_group_mask_0; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_mask_1 = io_mod_proc_mod_15_mat_mod_key_mod_group_mask_1; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_mask_2 = io_mod_proc_mod_15_mat_mod_key_mod_group_mask_2; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_mask_3 = io_mod_proc_mod_15_mat_mod_key_mod_group_mask_3; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_id_0 = io_mod_proc_mod_15_mat_mod_key_mod_group_id_0; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_id_1 = io_mod_proc_mod_15_mat_mod_key_mod_group_id_1; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_id_2 = io_mod_proc_mod_15_mat_mod_key_mod_group_id_2; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_key_mod_group_id_3 = io_mod_proc_mod_15_mat_mod_key_mod_group_id_3; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_table_mod_table_depth = io_mod_proc_mod_15_mat_mod_table_mod_table_depth; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_table_mod_table_width = io_mod_proc_mod_15_mat_mod_table_mod_table_width; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_w_en = io_mod_proc_mod_15_mat_mod_w_en; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_w_sram_id = io_mod_proc_mod_15_mat_mod_w_sram_id; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_w_addr = io_mod_proc_mod_15_mat_mod_w_addr; // @[pisa.scala 29:20]
  assign proc_15_io_mod_mat_mod_w_data = io_mod_proc_mod_15_mat_mod_w_data; // @[pisa.scala 29:20]
  assign proc_15_io_mod_exe_mod_en_0 = io_mod_proc_mod_15_exe_mod_en_0; // @[pisa.scala 29:20]
  assign proc_15_io_mod_exe_mod_en_1 = io_mod_proc_mod_15_exe_mod_en_1; // @[pisa.scala 29:20]
  assign proc_15_io_mod_exe_mod_addr = io_mod_proc_mod_15_exe_mod_addr; // @[pisa.scala 29:20]
  assign proc_15_io_mod_exe_mod_data_0 = io_mod_proc_mod_15_exe_mod_data_0; // @[pisa.scala 29:20]
  assign proc_15_io_mod_exe_mod_data_1 = io_mod_proc_mod_15_exe_mod_data_1; // @[pisa.scala 29:20]
endmodule
