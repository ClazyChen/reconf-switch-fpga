module Executor(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [2:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [2:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input         io_hit,
  input  [63:0] io_match_value,
  input         io_action_mod_en_0,
  input         io_action_mod_en_1,
  input  [7:0]  io_action_mod_addr,
  input  [63:0] io_action_mod_data_0,
  input  [63:0] io_action_mod_data_1
);
  wire  pipe1_clock; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[executor.scala 489:23]
  wire [2:0] pipe1_io_pipe_phv_in_next_processor_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 489:23]
  wire [2:0] pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[executor.scala 489:23]
  wire  pipe1_io_hit; // @[executor.scala 489:23]
  wire [63:0] pipe1_io_match_value; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_0; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_2; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_3; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_4; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_5; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_6; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_0; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_1; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_2; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_3; // @[executor.scala 489:23]
  wire  pipe1_io_action_mod_en_0; // @[executor.scala 489:23]
  wire  pipe1_io_action_mod_en_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_action_mod_addr; // @[executor.scala 489:23]
  wire [63:0] pipe1_io_action_mod_data_0; // @[executor.scala 489:23]
  wire [63:0] pipe1_io_action_mod_data_1; // @[executor.scala 489:23]
  wire  pipe2_clock; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[executor.scala 490:23]
  wire [2:0] pipe2_io_pipe_phv_in_next_processor_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 490:23]
  wire [2:0] pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_6; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_0; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_1; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_2; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_6; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_0; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_1; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_2; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_3; // @[executor.scala 490:23]
  wire  pipe3_clock; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_160; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_161; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_162; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_163; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_164; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_165; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_166; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_167; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_168; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_169; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_170; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_171; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_172; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_173; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_174; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_175; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_176; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_177; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_178; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_179; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_180; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_181; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_182; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_183; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_184; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_185; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_186; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_187; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_188; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_189; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_190; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_191; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_192; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_193; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_194; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_195; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_196; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_197; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_198; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_199; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_200; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_201; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_202; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_203; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_204; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_205; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_206; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_207; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_208; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_209; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_210; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_211; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_212; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_213; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_214; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_215; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_216; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_217; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_218; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_219; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_220; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_221; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_222; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_223; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_224; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_225; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_226; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_227; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_228; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_229; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_230; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_231; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_232; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_233; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_234; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_235; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_236; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_237; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_238; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_239; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_240; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_241; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_242; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_243; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_244; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_245; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_246; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_247; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_248; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_249; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_250; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_251; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_252; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_253; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_254; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_255; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[executor.scala 491:23]
  wire [2:0] pipe3_io_pipe_phv_in_next_processor_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_160; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_161; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_162; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_163; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_164; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_165; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_166; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_167; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_168; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_169; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_170; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_171; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_172; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_173; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_174; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_175; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_176; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_177; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_178; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_179; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_180; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_181; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_182; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_183; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_184; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_185; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_186; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_187; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_188; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_189; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_190; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_191; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_192; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_193; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_194; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_195; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_196; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_197; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_198; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_199; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_200; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_201; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_202; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_203; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_204; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_205; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_206; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_207; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_208; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_209; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_210; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_211; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_212; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_213; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_214; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_215; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_216; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_217; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_218; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_219; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_220; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_221; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_222; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_223; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_224; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_225; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_226; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_227; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_228; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_229; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_230; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_231; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_232; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_233; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_234; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_235; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_236; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_237; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_238; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_239; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_240; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_241; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_242; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_243; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_244; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_245; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_246; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_247; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_248; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_249; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_250; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_251; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_252; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_253; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_254; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_255; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 491:23]
  wire [2:0] pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_4; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_5; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_6; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_0; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_1; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_2; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_3; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_0; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_1; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_2; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_3; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_0; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_1; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_2; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_3; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_0; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_1; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_2; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_3; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_0; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_1; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_2; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_3; // @[executor.scala 491:23]
  wire  pipe4_clock; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_160; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_161; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_162; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_163; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_164; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_165; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_166; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_167; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_168; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_169; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_170; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_171; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_172; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_173; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_174; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_175; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_176; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_177; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_178; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_179; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_180; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_181; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_182; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_183; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_184; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_185; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_186; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_187; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_188; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_189; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_190; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_191; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_192; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_193; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_194; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_195; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_196; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_197; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_198; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_199; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_200; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_201; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_202; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_203; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_204; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_205; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_206; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_207; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_208; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_209; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_210; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_211; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_212; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_213; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_214; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_215; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_216; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_217; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_218; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_219; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_220; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_221; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_222; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_223; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_224; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_225; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_226; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_227; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_228; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_229; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_230; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_231; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_232; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_233; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_234; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_235; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_236; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_237; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_238; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_239; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_240; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_241; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_242; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_243; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_244; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_245; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_246; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_247; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_248; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_249; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_250; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_251; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_252; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_253; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_254; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_255; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[executor.scala 492:23]
  wire [2:0] pipe4_io_pipe_phv_in_next_processor_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_160; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_161; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_162; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_163; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_164; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_165; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_166; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_167; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_168; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_169; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_170; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_171; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_172; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_173; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_174; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_175; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_176; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_177; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_178; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_179; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_180; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_181; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_182; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_183; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_184; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_185; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_186; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_187; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_188; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_189; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_190; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_191; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_192; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_193; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_194; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_195; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_196; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_197; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_198; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_199; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_200; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_201; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_202; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_203; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_204; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_205; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_206; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_207; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_208; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_209; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_210; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_211; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_212; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_213; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_214; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_215; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_216; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_217; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_218; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_219; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_220; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_221; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_222; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_223; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_224; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_225; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_226; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_227; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_228; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_229; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_230; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_231; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_232; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_233; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_234; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_235; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_236; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_237; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_238; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_239; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_240; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_241; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_242; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_243; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_244; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_245; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_246; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_247; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_248; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_249; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_250; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_251; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_252; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_253; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_254; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_255; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 492:23]
  wire [2:0] pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_3; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_3; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_0; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_1; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_2; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_3; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_0; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_1; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_2; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_3; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_3; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_3; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_0; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_1; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_2; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_3; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_0; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_1; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_2; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_3; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_0; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_1; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_2; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_3; // @[executor.scala 492:23]
  wire  pipe5_clock; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_96; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_97; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_98; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_99; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_100; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_101; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_102; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_103; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_104; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_105; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_106; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_107; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_108; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_109; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_110; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_111; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_112; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_113; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_114; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_115; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_116; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_117; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_118; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_119; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_120; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_121; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_122; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_123; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_124; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_125; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_126; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_127; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_128; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_129; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_130; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_131; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_132; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_133; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_134; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_135; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_136; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_137; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_138; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_139; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_140; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_141; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_142; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_143; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_144; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_145; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_146; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_147; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_148; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_149; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_150; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_151; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_152; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_153; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_154; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_155; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_156; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_157; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_158; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_159; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_160; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_161; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_162; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_163; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_164; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_165; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_166; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_167; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_168; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_169; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_170; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_171; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_172; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_173; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_174; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_175; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_176; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_177; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_178; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_179; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_180; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_181; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_182; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_183; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_184; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_185; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_186; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_187; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_188; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_189; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_190; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_191; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_192; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_193; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_194; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_195; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_196; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_197; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_198; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_199; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_200; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_201; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_202; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_203; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_204; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_205; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_206; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_207; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_208; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_209; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_210; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_211; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_212; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_213; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_214; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_215; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_216; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_217; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_218; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_219; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_220; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_221; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_222; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_223; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_224; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_225; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_226; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_227; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_228; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_229; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_230; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_231; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_232; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_233; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_234; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_235; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_236; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_237; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_238; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_239; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_240; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_241; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_242; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_243; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_244; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_245; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_246; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_247; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_248; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_249; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_250; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_251; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_252; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_253; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_254; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_255; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[executor.scala 493:23]
  wire [2:0] pipe5_io_pipe_phv_in_next_processor_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_96; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_97; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_98; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_99; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_100; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_101; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_102; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_103; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_104; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_105; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_106; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_107; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_108; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_109; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_110; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_111; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_112; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_113; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_114; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_115; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_116; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_117; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_118; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_119; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_120; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_121; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_122; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_123; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_124; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_125; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_126; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_127; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_128; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_129; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_130; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_131; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_132; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_133; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_134; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_135; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_136; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_137; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_138; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_139; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_140; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_141; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_142; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_143; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_144; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_145; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_146; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_147; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_148; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_149; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_150; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_151; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_152; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_153; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_154; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_155; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_156; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_157; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_158; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_159; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_160; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_161; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_162; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_163; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_164; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_165; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_166; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_167; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_168; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_169; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_170; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_171; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_172; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_173; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_174; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_175; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_176; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_177; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_178; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_179; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_180; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_181; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_182; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_183; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_184; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_185; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_186; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_187; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_188; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_189; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_190; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_191; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_192; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_193; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_194; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_195; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_196; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_197; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_198; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_199; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_200; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_201; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_202; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_203; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_204; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_205; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_206; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_207; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_208; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_209; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_210; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_211; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_212; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_213; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_214; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_215; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_216; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_217; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_218; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_219; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_220; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_221; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_222; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_223; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_224; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_225; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_226; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_227; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_228; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_229; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_230; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_231; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_232; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_233; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_234; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_235; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_236; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_237; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_238; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_239; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_240; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_241; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_242; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_243; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_244; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_245; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_246; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_247; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_248; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_249; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_250; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_251; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_252; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_253; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_254; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_255; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 493:23]
  wire [2:0] pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_3; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_3; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_0; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_1; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_2; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_3; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_0; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_1; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_2; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_3; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_0; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_1; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_2; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_3; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_3; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_3; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_0; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_1; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_2; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_3; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_0; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_1; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_2; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_3; // @[executor.scala 493:23]
  wire  pipe6_clock; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_96; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_97; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_98; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_99; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_100; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_101; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_102; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_103; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_104; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_105; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_106; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_107; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_108; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_109; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_110; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_111; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_112; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_113; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_114; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_115; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_116; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_117; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_118; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_119; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_120; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_121; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_122; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_123; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_124; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_125; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_126; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_127; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_128; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_129; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_130; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_131; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_132; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_133; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_134; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_135; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_136; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_137; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_138; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_139; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_140; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_141; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_142; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_143; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_144; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_145; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_146; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_147; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_148; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_149; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_150; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_151; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_152; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_153; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_154; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_155; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_156; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_157; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_158; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_159; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_160; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_161; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_162; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_163; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_164; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_165; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_166; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_167; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_168; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_169; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_170; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_171; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_172; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_173; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_174; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_175; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_176; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_177; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_178; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_179; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_180; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_181; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_182; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_183; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_184; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_185; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_186; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_187; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_188; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_189; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_190; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_191; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_192; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_193; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_194; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_195; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_196; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_197; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_198; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_199; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_200; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_201; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_202; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_203; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_204; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_205; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_206; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_207; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_208; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_209; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_210; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_211; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_212; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_213; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_214; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_215; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_216; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_217; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_218; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_219; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_220; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_221; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_222; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_223; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_224; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_225; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_226; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_227; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_228; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_229; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_230; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_231; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_232; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_233; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_234; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_235; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_236; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_237; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_238; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_239; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_240; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_241; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_242; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_243; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_244; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_245; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_246; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_247; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_248; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_249; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_250; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_251; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_252; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_253; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_254; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_255; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[executor.scala 494:23]
  wire [2:0] pipe6_io_pipe_phv_in_next_processor_id; // @[executor.scala 494:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[executor.scala 494:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_96; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_97; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_98; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_99; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_100; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_101; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_102; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_103; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_104; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_105; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_106; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_107; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_108; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_109; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_110; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_111; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_112; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_113; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_114; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_115; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_116; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_117; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_118; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_119; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_120; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_121; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_122; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_123; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_124; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_125; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_126; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_127; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_128; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_129; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_130; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_131; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_132; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_133; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_134; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_135; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_136; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_137; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_138; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_139; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_140; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_141; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_142; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_143; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_144; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_145; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_146; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_147; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_148; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_149; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_150; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_151; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_152; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_153; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_154; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_155; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_156; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_157; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_158; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_159; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_160; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_161; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_162; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_163; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_164; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_165; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_166; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_167; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_168; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_169; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_170; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_171; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_172; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_173; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_174; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_175; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_176; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_177; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_178; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_179; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_180; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_181; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_182; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_183; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_184; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_185; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_186; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_187; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_188; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_189; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_190; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_191; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_192; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_193; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_194; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_195; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_196; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_197; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_198; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_199; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_200; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_201; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_202; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_203; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_204; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_205; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_206; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_207; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_208; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_209; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_210; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_211; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_212; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_213; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_214; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_215; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_216; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_217; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_218; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_219; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_220; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_221; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_222; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_223; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_224; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_225; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_226; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_227; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_228; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_229; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_230; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_231; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_232; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_233; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_234; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_235; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_236; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_237; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_238; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_239; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_240; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_241; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_242; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_243; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_244; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_245; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_246; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_247; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_248; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_249; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_250; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_251; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_252; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_253; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_254; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_255; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 494:23]
  wire [2:0] pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 494:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_0; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_1; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_2; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_3; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_0; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_1; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_2; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_3; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_0; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_1; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_2; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_3; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_0; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_1; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_2; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_3; // @[executor.scala 494:23]
  ActionReader pipe1 ( // @[executor.scala 489:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_hit(pipe1_io_hit),
    .io_match_value(pipe1_io_match_value),
    .io_args_out_0(pipe1_io_args_out_0),
    .io_args_out_1(pipe1_io_args_out_1),
    .io_args_out_2(pipe1_io_args_out_2),
    .io_args_out_3(pipe1_io_args_out_3),
    .io_args_out_4(pipe1_io_args_out_4),
    .io_args_out_5(pipe1_io_args_out_5),
    .io_args_out_6(pipe1_io_args_out_6),
    .io_vliw_out_0(pipe1_io_vliw_out_0),
    .io_vliw_out_1(pipe1_io_vliw_out_1),
    .io_vliw_out_2(pipe1_io_vliw_out_2),
    .io_vliw_out_3(pipe1_io_vliw_out_3),
    .io_action_mod_en_0(pipe1_io_action_mod_en_0),
    .io_action_mod_en_1(pipe1_io_action_mod_en_1),
    .io_action_mod_addr(pipe1_io_action_mod_addr),
    .io_action_mod_data_0(pipe1_io_action_mod_data_0),
    .io_action_mod_data_1(pipe1_io_action_mod_data_1)
  );
  PrimitiveGetOffset pipe2 ( // @[executor.scala 490:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe2_io_args_in_0),
    .io_args_in_1(pipe2_io_args_in_1),
    .io_args_in_2(pipe2_io_args_in_2),
    .io_args_in_3(pipe2_io_args_in_3),
    .io_args_in_4(pipe2_io_args_in_4),
    .io_args_in_5(pipe2_io_args_in_5),
    .io_args_in_6(pipe2_io_args_in_6),
    .io_vliw_in_0(pipe2_io_vliw_in_0),
    .io_vliw_in_1(pipe2_io_vliw_in_1),
    .io_vliw_in_2(pipe2_io_vliw_in_2),
    .io_vliw_in_3(pipe2_io_vliw_in_3),
    .io_args_out_0(pipe2_io_args_out_0),
    .io_args_out_1(pipe2_io_args_out_1),
    .io_args_out_2(pipe2_io_args_out_2),
    .io_args_out_3(pipe2_io_args_out_3),
    .io_args_out_4(pipe2_io_args_out_4),
    .io_args_out_5(pipe2_io_args_out_5),
    .io_args_out_6(pipe2_io_args_out_6),
    .io_vliw_out_0(pipe2_io_vliw_out_0),
    .io_vliw_out_1(pipe2_io_vliw_out_1),
    .io_vliw_out_2(pipe2_io_vliw_out_2),
    .io_vliw_out_3(pipe2_io_vliw_out_3),
    .io_offset_out_0(pipe2_io_offset_out_0),
    .io_offset_out_1(pipe2_io_offset_out_1),
    .io_offset_out_2(pipe2_io_offset_out_2),
    .io_offset_out_3(pipe2_io_offset_out_3),
    .io_length_out_0(pipe2_io_length_out_0),
    .io_length_out_1(pipe2_io_length_out_1),
    .io_length_out_2(pipe2_io_length_out_2),
    .io_length_out_3(pipe2_io_length_out_3)
  );
  PrimitiveGetSource pipe3 ( // @[executor.scala 491:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe3_io_args_in_0),
    .io_args_in_1(pipe3_io_args_in_1),
    .io_args_in_2(pipe3_io_args_in_2),
    .io_args_in_3(pipe3_io_args_in_3),
    .io_args_in_4(pipe3_io_args_in_4),
    .io_args_in_5(pipe3_io_args_in_5),
    .io_args_in_6(pipe3_io_args_in_6),
    .io_vliw_in_0(pipe3_io_vliw_in_0),
    .io_vliw_in_1(pipe3_io_vliw_in_1),
    .io_vliw_in_2(pipe3_io_vliw_in_2),
    .io_vliw_in_3(pipe3_io_vliw_in_3),
    .io_offset_in_0(pipe3_io_offset_in_0),
    .io_offset_in_1(pipe3_io_offset_in_1),
    .io_offset_in_2(pipe3_io_offset_in_2),
    .io_offset_in_3(pipe3_io_offset_in_3),
    .io_length_in_0(pipe3_io_length_in_0),
    .io_length_in_1(pipe3_io_length_in_1),
    .io_length_in_2(pipe3_io_length_in_2),
    .io_length_in_3(pipe3_io_length_in_3),
    .io_vliw_out_0(pipe3_io_vliw_out_0),
    .io_vliw_out_1(pipe3_io_vliw_out_1),
    .io_vliw_out_2(pipe3_io_vliw_out_2),
    .io_vliw_out_3(pipe3_io_vliw_out_3),
    .io_field_out_0(pipe3_io_field_out_0),
    .io_field_out_1(pipe3_io_field_out_1),
    .io_field_out_2(pipe3_io_field_out_2),
    .io_field_out_3(pipe3_io_field_out_3),
    .io_mask_out_0(pipe3_io_mask_out_0),
    .io_mask_out_1(pipe3_io_mask_out_1),
    .io_mask_out_2(pipe3_io_mask_out_2),
    .io_mask_out_3(pipe3_io_mask_out_3),
    .io_bias_out_0(pipe3_io_bias_out_0),
    .io_bias_out_1(pipe3_io_bias_out_1),
    .io_bias_out_2(pipe3_io_bias_out_2),
    .io_bias_out_3(pipe3_io_bias_out_3)
  );
  PrimitiveShiftSource pipe4 ( // @[executor.scala 492:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_vliw_in_0(pipe4_io_vliw_in_0),
    .io_vliw_in_1(pipe4_io_vliw_in_1),
    .io_vliw_in_2(pipe4_io_vliw_in_2),
    .io_vliw_in_3(pipe4_io_vliw_in_3),
    .io_field_in_0(pipe4_io_field_in_0),
    .io_field_in_1(pipe4_io_field_in_1),
    .io_field_in_2(pipe4_io_field_in_2),
    .io_field_in_3(pipe4_io_field_in_3),
    .io_mask_in_0(pipe4_io_mask_in_0),
    .io_mask_in_1(pipe4_io_mask_in_1),
    .io_mask_in_2(pipe4_io_mask_in_2),
    .io_mask_in_3(pipe4_io_mask_in_3),
    .io_bias_in_0(pipe4_io_bias_in_0),
    .io_bias_in_1(pipe4_io_bias_in_1),
    .io_bias_in_2(pipe4_io_bias_in_2),
    .io_bias_in_3(pipe4_io_bias_in_3),
    .io_vliw_out_0(pipe4_io_vliw_out_0),
    .io_vliw_out_1(pipe4_io_vliw_out_1),
    .io_vliw_out_2(pipe4_io_vliw_out_2),
    .io_vliw_out_3(pipe4_io_vliw_out_3),
    .io_field_out_0(pipe4_io_field_out_0),
    .io_field_out_1(pipe4_io_field_out_1),
    .io_field_out_2(pipe4_io_field_out_2),
    .io_field_out_3(pipe4_io_field_out_3),
    .io_mask_out_0(pipe4_io_mask_out_0),
    .io_mask_out_1(pipe4_io_mask_out_1),
    .io_mask_out_2(pipe4_io_mask_out_2),
    .io_mask_out_3(pipe4_io_mask_out_3),
    .io_bias_out_0(pipe4_io_bias_out_0),
    .io_bias_out_1(pipe4_io_bias_out_1),
    .io_bias_out_2(pipe4_io_bias_out_2),
    .io_bias_out_3(pipe4_io_bias_out_3),
    .io_dst_offset_out_0(pipe4_io_dst_offset_out_0),
    .io_dst_offset_out_1(pipe4_io_dst_offset_out_1),
    .io_dst_offset_out_2(pipe4_io_dst_offset_out_2),
    .io_dst_offset_out_3(pipe4_io_dst_offset_out_3)
  );
  PrimitiveALU pipe5 ( // @[executor.scala 493:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe5_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe5_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe5_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe5_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe5_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe5_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe5_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe5_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe5_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe5_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe5_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe5_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe5_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe5_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe5_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe5_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe5_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe5_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe5_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe5_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe5_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe5_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe5_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe5_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe5_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe5_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe5_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe5_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe5_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe5_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe5_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe5_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe5_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe5_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe5_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe5_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe5_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe5_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe5_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe5_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe5_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe5_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe5_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe5_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe5_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe5_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe5_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe5_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe5_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe5_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe5_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe5_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe5_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe5_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe5_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe5_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe5_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe5_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe5_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe5_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe5_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe5_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe5_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe5_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe5_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe5_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe5_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe5_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe5_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe5_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe5_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe5_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe5_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe5_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe5_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe5_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe5_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe5_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe5_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe5_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe5_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe5_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe5_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe5_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe5_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe5_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe5_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe5_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe5_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe5_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe5_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe5_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe5_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe5_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe5_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe5_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe5_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe5_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe5_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe5_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe5_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe5_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe5_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe5_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe5_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe5_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe5_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe5_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe5_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe5_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe5_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe5_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe5_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe5_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe5_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe5_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe5_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe5_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe5_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe5_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe5_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe5_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe5_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe5_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe5_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe5_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe5_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe5_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe5_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe5_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe5_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe5_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe5_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe5_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe5_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe5_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe5_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe5_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe5_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe5_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe5_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe5_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe5_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe5_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe5_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe5_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe5_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe5_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe5_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe5_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe5_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe5_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe5_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe5_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe5_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe5_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe5_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe5_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe5_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe5_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe5_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe5_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe5_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe5_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe5_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe5_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe5_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe5_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe5_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe5_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe5_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe5_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe5_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe5_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe5_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe5_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe5_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe5_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe5_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe5_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe5_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe5_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe5_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe5_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe5_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe5_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe5_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe5_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe5_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe5_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe5_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe5_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_vliw_in_0(pipe5_io_vliw_in_0),
    .io_vliw_in_1(pipe5_io_vliw_in_1),
    .io_vliw_in_2(pipe5_io_vliw_in_2),
    .io_vliw_in_3(pipe5_io_vliw_in_3),
    .io_field_in_0(pipe5_io_field_in_0),
    .io_field_in_1(pipe5_io_field_in_1),
    .io_field_in_2(pipe5_io_field_in_2),
    .io_field_in_3(pipe5_io_field_in_3),
    .io_mask_in_0(pipe5_io_mask_in_0),
    .io_mask_in_1(pipe5_io_mask_in_1),
    .io_mask_in_2(pipe5_io_mask_in_2),
    .io_mask_in_3(pipe5_io_mask_in_3),
    .io_bias_in_0(pipe5_io_bias_in_0),
    .io_bias_in_1(pipe5_io_bias_in_1),
    .io_bias_in_2(pipe5_io_bias_in_2),
    .io_bias_in_3(pipe5_io_bias_in_3),
    .io_dst_offset_in_0(pipe5_io_dst_offset_in_0),
    .io_dst_offset_in_1(pipe5_io_dst_offset_in_1),
    .io_dst_offset_in_2(pipe5_io_dst_offset_in_2),
    .io_dst_offset_in_3(pipe5_io_dst_offset_in_3),
    .io_vliw_out_0(pipe5_io_vliw_out_0),
    .io_vliw_out_1(pipe5_io_vliw_out_1),
    .io_vliw_out_2(pipe5_io_vliw_out_2),
    .io_vliw_out_3(pipe5_io_vliw_out_3),
    .io_field_out_0(pipe5_io_field_out_0),
    .io_field_out_1(pipe5_io_field_out_1),
    .io_field_out_2(pipe5_io_field_out_2),
    .io_field_out_3(pipe5_io_field_out_3),
    .io_mask_out_0(pipe5_io_mask_out_0),
    .io_mask_out_1(pipe5_io_mask_out_1),
    .io_mask_out_2(pipe5_io_mask_out_2),
    .io_mask_out_3(pipe5_io_mask_out_3),
    .io_dst_offset_out_0(pipe5_io_dst_offset_out_0),
    .io_dst_offset_out_1(pipe5_io_dst_offset_out_1),
    .io_dst_offset_out_2(pipe5_io_dst_offset_out_2),
    .io_dst_offset_out_3(pipe5_io_dst_offset_out_3)
  );
  PrimitiveWriteBack pipe6 ( // @[executor.scala 494:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe6_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe6_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe6_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe6_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe6_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe6_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe6_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe6_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe6_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe6_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe6_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe6_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe6_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe6_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe6_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe6_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe6_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe6_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe6_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe6_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe6_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe6_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe6_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe6_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe6_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe6_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe6_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe6_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe6_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe6_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe6_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe6_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe6_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe6_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe6_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe6_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe6_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe6_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe6_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe6_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe6_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe6_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe6_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe6_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe6_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe6_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe6_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe6_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe6_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe6_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe6_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe6_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe6_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe6_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe6_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe6_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe6_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe6_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe6_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe6_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe6_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe6_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe6_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe6_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe6_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe6_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe6_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe6_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe6_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe6_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe6_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe6_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe6_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe6_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe6_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe6_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe6_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe6_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe6_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe6_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe6_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe6_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe6_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe6_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe6_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe6_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe6_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe6_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe6_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe6_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe6_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe6_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe6_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe6_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe6_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe6_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe6_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe6_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe6_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe6_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe6_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe6_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe6_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe6_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe6_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe6_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe6_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe6_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe6_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe6_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe6_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe6_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe6_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe6_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe6_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe6_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe6_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe6_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe6_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe6_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe6_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe6_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe6_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe6_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe6_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe6_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe6_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe6_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe6_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe6_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe6_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe6_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe6_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe6_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe6_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe6_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe6_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe6_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe6_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe6_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe6_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe6_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe6_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe6_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe6_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe6_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe6_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe6_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe6_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe6_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe6_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe6_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe6_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe6_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe6_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe6_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe6_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe6_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe6_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe6_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe6_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe6_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe6_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe6_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe6_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe6_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe6_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe6_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe6_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe6_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe6_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe6_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe6_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe6_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe6_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe6_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe6_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe6_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe6_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe6_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe6_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe6_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe6_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe6_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe6_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe6_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe6_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe6_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe6_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe6_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe6_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe6_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_vliw_in_0(pipe6_io_vliw_in_0),
    .io_vliw_in_1(pipe6_io_vliw_in_1),
    .io_vliw_in_2(pipe6_io_vliw_in_2),
    .io_vliw_in_3(pipe6_io_vliw_in_3),
    .io_field_in_0(pipe6_io_field_in_0),
    .io_field_in_1(pipe6_io_field_in_1),
    .io_field_in_2(pipe6_io_field_in_2),
    .io_field_in_3(pipe6_io_field_in_3),
    .io_mask_in_0(pipe6_io_mask_in_0),
    .io_mask_in_1(pipe6_io_mask_in_1),
    .io_mask_in_2(pipe6_io_mask_in_2),
    .io_mask_in_3(pipe6_io_mask_in_3),
    .io_dst_offset_in_0(pipe6_io_dst_offset_in_0),
    .io_dst_offset_in_1(pipe6_io_dst_offset_in_1),
    .io_dst_offset_in_2(pipe6_io_dst_offset_in_2),
    .io_dst_offset_in_3(pipe6_io_dst_offset_in_3)
  );
  assign io_pipe_phv_out_data_0 = pipe6_io_pipe_phv_out_data_0; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_1 = pipe6_io_pipe_phv_out_data_1; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_2 = pipe6_io_pipe_phv_out_data_2; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_3 = pipe6_io_pipe_phv_out_data_3; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_4 = pipe6_io_pipe_phv_out_data_4; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_5 = pipe6_io_pipe_phv_out_data_5; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_6 = pipe6_io_pipe_phv_out_data_6; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_7 = pipe6_io_pipe_phv_out_data_7; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_8 = pipe6_io_pipe_phv_out_data_8; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_9 = pipe6_io_pipe_phv_out_data_9; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_10 = pipe6_io_pipe_phv_out_data_10; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_11 = pipe6_io_pipe_phv_out_data_11; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_12 = pipe6_io_pipe_phv_out_data_12; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_13 = pipe6_io_pipe_phv_out_data_13; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_14 = pipe6_io_pipe_phv_out_data_14; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_15 = pipe6_io_pipe_phv_out_data_15; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_16 = pipe6_io_pipe_phv_out_data_16; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_17 = pipe6_io_pipe_phv_out_data_17; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_18 = pipe6_io_pipe_phv_out_data_18; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_19 = pipe6_io_pipe_phv_out_data_19; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_20 = pipe6_io_pipe_phv_out_data_20; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_21 = pipe6_io_pipe_phv_out_data_21; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_22 = pipe6_io_pipe_phv_out_data_22; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_23 = pipe6_io_pipe_phv_out_data_23; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_24 = pipe6_io_pipe_phv_out_data_24; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_25 = pipe6_io_pipe_phv_out_data_25; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_26 = pipe6_io_pipe_phv_out_data_26; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_27 = pipe6_io_pipe_phv_out_data_27; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_28 = pipe6_io_pipe_phv_out_data_28; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_29 = pipe6_io_pipe_phv_out_data_29; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_30 = pipe6_io_pipe_phv_out_data_30; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_31 = pipe6_io_pipe_phv_out_data_31; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_32 = pipe6_io_pipe_phv_out_data_32; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_33 = pipe6_io_pipe_phv_out_data_33; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_34 = pipe6_io_pipe_phv_out_data_34; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_35 = pipe6_io_pipe_phv_out_data_35; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_36 = pipe6_io_pipe_phv_out_data_36; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_37 = pipe6_io_pipe_phv_out_data_37; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_38 = pipe6_io_pipe_phv_out_data_38; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_39 = pipe6_io_pipe_phv_out_data_39; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_40 = pipe6_io_pipe_phv_out_data_40; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_41 = pipe6_io_pipe_phv_out_data_41; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_42 = pipe6_io_pipe_phv_out_data_42; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_43 = pipe6_io_pipe_phv_out_data_43; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_44 = pipe6_io_pipe_phv_out_data_44; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_45 = pipe6_io_pipe_phv_out_data_45; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_46 = pipe6_io_pipe_phv_out_data_46; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_47 = pipe6_io_pipe_phv_out_data_47; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_48 = pipe6_io_pipe_phv_out_data_48; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_49 = pipe6_io_pipe_phv_out_data_49; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_50 = pipe6_io_pipe_phv_out_data_50; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_51 = pipe6_io_pipe_phv_out_data_51; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_52 = pipe6_io_pipe_phv_out_data_52; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_53 = pipe6_io_pipe_phv_out_data_53; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_54 = pipe6_io_pipe_phv_out_data_54; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_55 = pipe6_io_pipe_phv_out_data_55; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_56 = pipe6_io_pipe_phv_out_data_56; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_57 = pipe6_io_pipe_phv_out_data_57; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_58 = pipe6_io_pipe_phv_out_data_58; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_59 = pipe6_io_pipe_phv_out_data_59; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_60 = pipe6_io_pipe_phv_out_data_60; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_61 = pipe6_io_pipe_phv_out_data_61; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_62 = pipe6_io_pipe_phv_out_data_62; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_63 = pipe6_io_pipe_phv_out_data_63; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_64 = pipe6_io_pipe_phv_out_data_64; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_65 = pipe6_io_pipe_phv_out_data_65; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_66 = pipe6_io_pipe_phv_out_data_66; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_67 = pipe6_io_pipe_phv_out_data_67; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_68 = pipe6_io_pipe_phv_out_data_68; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_69 = pipe6_io_pipe_phv_out_data_69; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_70 = pipe6_io_pipe_phv_out_data_70; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_71 = pipe6_io_pipe_phv_out_data_71; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_72 = pipe6_io_pipe_phv_out_data_72; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_73 = pipe6_io_pipe_phv_out_data_73; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_74 = pipe6_io_pipe_phv_out_data_74; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_75 = pipe6_io_pipe_phv_out_data_75; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_76 = pipe6_io_pipe_phv_out_data_76; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_77 = pipe6_io_pipe_phv_out_data_77; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_78 = pipe6_io_pipe_phv_out_data_78; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_79 = pipe6_io_pipe_phv_out_data_79; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_80 = pipe6_io_pipe_phv_out_data_80; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_81 = pipe6_io_pipe_phv_out_data_81; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_82 = pipe6_io_pipe_phv_out_data_82; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_83 = pipe6_io_pipe_phv_out_data_83; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_84 = pipe6_io_pipe_phv_out_data_84; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_85 = pipe6_io_pipe_phv_out_data_85; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_86 = pipe6_io_pipe_phv_out_data_86; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_87 = pipe6_io_pipe_phv_out_data_87; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_88 = pipe6_io_pipe_phv_out_data_88; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_89 = pipe6_io_pipe_phv_out_data_89; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_90 = pipe6_io_pipe_phv_out_data_90; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_91 = pipe6_io_pipe_phv_out_data_91; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_92 = pipe6_io_pipe_phv_out_data_92; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_93 = pipe6_io_pipe_phv_out_data_93; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_94 = pipe6_io_pipe_phv_out_data_94; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_95 = pipe6_io_pipe_phv_out_data_95; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_96 = pipe6_io_pipe_phv_out_data_96; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_97 = pipe6_io_pipe_phv_out_data_97; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_98 = pipe6_io_pipe_phv_out_data_98; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_99 = pipe6_io_pipe_phv_out_data_99; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_100 = pipe6_io_pipe_phv_out_data_100; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_101 = pipe6_io_pipe_phv_out_data_101; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_102 = pipe6_io_pipe_phv_out_data_102; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_103 = pipe6_io_pipe_phv_out_data_103; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_104 = pipe6_io_pipe_phv_out_data_104; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_105 = pipe6_io_pipe_phv_out_data_105; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_106 = pipe6_io_pipe_phv_out_data_106; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_107 = pipe6_io_pipe_phv_out_data_107; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_108 = pipe6_io_pipe_phv_out_data_108; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_109 = pipe6_io_pipe_phv_out_data_109; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_110 = pipe6_io_pipe_phv_out_data_110; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_111 = pipe6_io_pipe_phv_out_data_111; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_112 = pipe6_io_pipe_phv_out_data_112; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_113 = pipe6_io_pipe_phv_out_data_113; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_114 = pipe6_io_pipe_phv_out_data_114; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_115 = pipe6_io_pipe_phv_out_data_115; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_116 = pipe6_io_pipe_phv_out_data_116; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_117 = pipe6_io_pipe_phv_out_data_117; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_118 = pipe6_io_pipe_phv_out_data_118; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_119 = pipe6_io_pipe_phv_out_data_119; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_120 = pipe6_io_pipe_phv_out_data_120; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_121 = pipe6_io_pipe_phv_out_data_121; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_122 = pipe6_io_pipe_phv_out_data_122; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_123 = pipe6_io_pipe_phv_out_data_123; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_124 = pipe6_io_pipe_phv_out_data_124; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_125 = pipe6_io_pipe_phv_out_data_125; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_126 = pipe6_io_pipe_phv_out_data_126; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_127 = pipe6_io_pipe_phv_out_data_127; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_128 = pipe6_io_pipe_phv_out_data_128; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_129 = pipe6_io_pipe_phv_out_data_129; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_130 = pipe6_io_pipe_phv_out_data_130; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_131 = pipe6_io_pipe_phv_out_data_131; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_132 = pipe6_io_pipe_phv_out_data_132; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_133 = pipe6_io_pipe_phv_out_data_133; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_134 = pipe6_io_pipe_phv_out_data_134; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_135 = pipe6_io_pipe_phv_out_data_135; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_136 = pipe6_io_pipe_phv_out_data_136; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_137 = pipe6_io_pipe_phv_out_data_137; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_138 = pipe6_io_pipe_phv_out_data_138; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_139 = pipe6_io_pipe_phv_out_data_139; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_140 = pipe6_io_pipe_phv_out_data_140; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_141 = pipe6_io_pipe_phv_out_data_141; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_142 = pipe6_io_pipe_phv_out_data_142; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_143 = pipe6_io_pipe_phv_out_data_143; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_144 = pipe6_io_pipe_phv_out_data_144; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_145 = pipe6_io_pipe_phv_out_data_145; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_146 = pipe6_io_pipe_phv_out_data_146; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_147 = pipe6_io_pipe_phv_out_data_147; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_148 = pipe6_io_pipe_phv_out_data_148; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_149 = pipe6_io_pipe_phv_out_data_149; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_150 = pipe6_io_pipe_phv_out_data_150; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_151 = pipe6_io_pipe_phv_out_data_151; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_152 = pipe6_io_pipe_phv_out_data_152; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_153 = pipe6_io_pipe_phv_out_data_153; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_154 = pipe6_io_pipe_phv_out_data_154; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_155 = pipe6_io_pipe_phv_out_data_155; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_156 = pipe6_io_pipe_phv_out_data_156; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_157 = pipe6_io_pipe_phv_out_data_157; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_158 = pipe6_io_pipe_phv_out_data_158; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_159 = pipe6_io_pipe_phv_out_data_159; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_160 = pipe6_io_pipe_phv_out_data_160; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_161 = pipe6_io_pipe_phv_out_data_161; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_162 = pipe6_io_pipe_phv_out_data_162; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_163 = pipe6_io_pipe_phv_out_data_163; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_164 = pipe6_io_pipe_phv_out_data_164; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_165 = pipe6_io_pipe_phv_out_data_165; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_166 = pipe6_io_pipe_phv_out_data_166; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_167 = pipe6_io_pipe_phv_out_data_167; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_168 = pipe6_io_pipe_phv_out_data_168; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_169 = pipe6_io_pipe_phv_out_data_169; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_170 = pipe6_io_pipe_phv_out_data_170; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_171 = pipe6_io_pipe_phv_out_data_171; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_172 = pipe6_io_pipe_phv_out_data_172; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_173 = pipe6_io_pipe_phv_out_data_173; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_174 = pipe6_io_pipe_phv_out_data_174; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_175 = pipe6_io_pipe_phv_out_data_175; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_176 = pipe6_io_pipe_phv_out_data_176; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_177 = pipe6_io_pipe_phv_out_data_177; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_178 = pipe6_io_pipe_phv_out_data_178; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_179 = pipe6_io_pipe_phv_out_data_179; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_180 = pipe6_io_pipe_phv_out_data_180; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_181 = pipe6_io_pipe_phv_out_data_181; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_182 = pipe6_io_pipe_phv_out_data_182; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_183 = pipe6_io_pipe_phv_out_data_183; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_184 = pipe6_io_pipe_phv_out_data_184; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_185 = pipe6_io_pipe_phv_out_data_185; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_186 = pipe6_io_pipe_phv_out_data_186; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_187 = pipe6_io_pipe_phv_out_data_187; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_188 = pipe6_io_pipe_phv_out_data_188; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_189 = pipe6_io_pipe_phv_out_data_189; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_190 = pipe6_io_pipe_phv_out_data_190; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_191 = pipe6_io_pipe_phv_out_data_191; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_192 = pipe6_io_pipe_phv_out_data_192; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_193 = pipe6_io_pipe_phv_out_data_193; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_194 = pipe6_io_pipe_phv_out_data_194; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_195 = pipe6_io_pipe_phv_out_data_195; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_196 = pipe6_io_pipe_phv_out_data_196; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_197 = pipe6_io_pipe_phv_out_data_197; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_198 = pipe6_io_pipe_phv_out_data_198; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_199 = pipe6_io_pipe_phv_out_data_199; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_200 = pipe6_io_pipe_phv_out_data_200; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_201 = pipe6_io_pipe_phv_out_data_201; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_202 = pipe6_io_pipe_phv_out_data_202; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_203 = pipe6_io_pipe_phv_out_data_203; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_204 = pipe6_io_pipe_phv_out_data_204; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_205 = pipe6_io_pipe_phv_out_data_205; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_206 = pipe6_io_pipe_phv_out_data_206; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_207 = pipe6_io_pipe_phv_out_data_207; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_208 = pipe6_io_pipe_phv_out_data_208; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_209 = pipe6_io_pipe_phv_out_data_209; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_210 = pipe6_io_pipe_phv_out_data_210; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_211 = pipe6_io_pipe_phv_out_data_211; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_212 = pipe6_io_pipe_phv_out_data_212; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_213 = pipe6_io_pipe_phv_out_data_213; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_214 = pipe6_io_pipe_phv_out_data_214; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_215 = pipe6_io_pipe_phv_out_data_215; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_216 = pipe6_io_pipe_phv_out_data_216; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_217 = pipe6_io_pipe_phv_out_data_217; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_218 = pipe6_io_pipe_phv_out_data_218; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_219 = pipe6_io_pipe_phv_out_data_219; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_220 = pipe6_io_pipe_phv_out_data_220; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_221 = pipe6_io_pipe_phv_out_data_221; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_222 = pipe6_io_pipe_phv_out_data_222; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_223 = pipe6_io_pipe_phv_out_data_223; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_224 = pipe6_io_pipe_phv_out_data_224; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_225 = pipe6_io_pipe_phv_out_data_225; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_226 = pipe6_io_pipe_phv_out_data_226; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_227 = pipe6_io_pipe_phv_out_data_227; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_228 = pipe6_io_pipe_phv_out_data_228; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_229 = pipe6_io_pipe_phv_out_data_229; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_230 = pipe6_io_pipe_phv_out_data_230; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_231 = pipe6_io_pipe_phv_out_data_231; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_232 = pipe6_io_pipe_phv_out_data_232; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_233 = pipe6_io_pipe_phv_out_data_233; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_234 = pipe6_io_pipe_phv_out_data_234; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_235 = pipe6_io_pipe_phv_out_data_235; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_236 = pipe6_io_pipe_phv_out_data_236; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_237 = pipe6_io_pipe_phv_out_data_237; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_238 = pipe6_io_pipe_phv_out_data_238; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_239 = pipe6_io_pipe_phv_out_data_239; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_240 = pipe6_io_pipe_phv_out_data_240; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_241 = pipe6_io_pipe_phv_out_data_241; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_242 = pipe6_io_pipe_phv_out_data_242; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_243 = pipe6_io_pipe_phv_out_data_243; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_244 = pipe6_io_pipe_phv_out_data_244; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_245 = pipe6_io_pipe_phv_out_data_245; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_246 = pipe6_io_pipe_phv_out_data_246; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_247 = pipe6_io_pipe_phv_out_data_247; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_248 = pipe6_io_pipe_phv_out_data_248; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_249 = pipe6_io_pipe_phv_out_data_249; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_250 = pipe6_io_pipe_phv_out_data_250; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_251 = pipe6_io_pipe_phv_out_data_251; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_252 = pipe6_io_pipe_phv_out_data_252; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_253 = pipe6_io_pipe_phv_out_data_253; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_254 = pipe6_io_pipe_phv_out_data_254; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_255 = pipe6_io_pipe_phv_out_data_255; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_0 = pipe6_io_pipe_phv_out_header_0; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_1 = pipe6_io_pipe_phv_out_header_1; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_2 = pipe6_io_pipe_phv_out_header_2; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_3 = pipe6_io_pipe_phv_out_header_3; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_4 = pipe6_io_pipe_phv_out_header_4; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_5 = pipe6_io_pipe_phv_out_header_5; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_6 = pipe6_io_pipe_phv_out_header_6; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_7 = pipe6_io_pipe_phv_out_header_7; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_8 = pipe6_io_pipe_phv_out_header_8; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_9 = pipe6_io_pipe_phv_out_header_9; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_10 = pipe6_io_pipe_phv_out_header_10; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_11 = pipe6_io_pipe_phv_out_header_11; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_12 = pipe6_io_pipe_phv_out_header_12; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_13 = pipe6_io_pipe_phv_out_header_13; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_14 = pipe6_io_pipe_phv_out_header_14; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_15 = pipe6_io_pipe_phv_out_header_15; // @[executor.scala 530:27]
  assign io_pipe_phv_out_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 530:27]
  assign io_pipe_phv_out_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 530:27]
  assign io_pipe_phv_out_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 530:27]
  assign io_pipe_phv_out_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 530:27]
  assign io_pipe_phv_out_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[executor.scala 530:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[executor.scala 496:26]
  assign pipe1_io_hit = io_hit; // @[executor.scala 497:26]
  assign pipe1_io_match_value = io_match_value; // @[executor.scala 498:26]
  assign pipe1_io_action_mod_en_0 = io_action_mod_en_0; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_en_1 = io_action_mod_en_1; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_addr = io_action_mod_addr; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_data_0 = io_action_mod_data_0; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_data_1 = io_action_mod_data_1; // @[executor.scala 499:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[executor.scala 501:26]
  assign pipe2_io_args_in_0 = pipe1_io_args_out_0; // @[executor.scala 502:26]
  assign pipe2_io_args_in_1 = pipe1_io_args_out_1; // @[executor.scala 502:26]
  assign pipe2_io_args_in_2 = pipe1_io_args_out_2; // @[executor.scala 502:26]
  assign pipe2_io_args_in_3 = pipe1_io_args_out_3; // @[executor.scala 502:26]
  assign pipe2_io_args_in_4 = pipe1_io_args_out_4; // @[executor.scala 502:26]
  assign pipe2_io_args_in_5 = pipe1_io_args_out_5; // @[executor.scala 502:26]
  assign pipe2_io_args_in_6 = pipe1_io_args_out_6; // @[executor.scala 502:26]
  assign pipe2_io_vliw_in_0 = pipe1_io_vliw_out_0; // @[executor.scala 503:26]
  assign pipe2_io_vliw_in_1 = pipe1_io_vliw_out_1; // @[executor.scala 503:26]
  assign pipe2_io_vliw_in_2 = pipe1_io_vliw_out_2; // @[executor.scala 503:26]
  assign pipe2_io_vliw_in_3 = pipe1_io_vliw_out_3; // @[executor.scala 503:26]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[executor.scala 505:26]
  assign pipe3_io_args_in_0 = pipe2_io_args_out_0; // @[executor.scala 506:26]
  assign pipe3_io_args_in_1 = pipe2_io_args_out_1; // @[executor.scala 506:26]
  assign pipe3_io_args_in_2 = pipe2_io_args_out_2; // @[executor.scala 506:26]
  assign pipe3_io_args_in_3 = pipe2_io_args_out_3; // @[executor.scala 506:26]
  assign pipe3_io_args_in_4 = pipe2_io_args_out_4; // @[executor.scala 506:26]
  assign pipe3_io_args_in_5 = pipe2_io_args_out_5; // @[executor.scala 506:26]
  assign pipe3_io_args_in_6 = pipe2_io_args_out_6; // @[executor.scala 506:26]
  assign pipe3_io_vliw_in_0 = pipe2_io_vliw_out_0; // @[executor.scala 507:26]
  assign pipe3_io_vliw_in_1 = pipe2_io_vliw_out_1; // @[executor.scala 507:26]
  assign pipe3_io_vliw_in_2 = pipe2_io_vliw_out_2; // @[executor.scala 507:26]
  assign pipe3_io_vliw_in_3 = pipe2_io_vliw_out_3; // @[executor.scala 507:26]
  assign pipe3_io_offset_in_0 = pipe2_io_offset_out_0; // @[executor.scala 508:26]
  assign pipe3_io_offset_in_1 = pipe2_io_offset_out_1; // @[executor.scala 508:26]
  assign pipe3_io_offset_in_2 = pipe2_io_offset_out_2; // @[executor.scala 508:26]
  assign pipe3_io_offset_in_3 = pipe2_io_offset_out_3; // @[executor.scala 508:26]
  assign pipe3_io_length_in_0 = pipe2_io_length_out_0; // @[executor.scala 509:26]
  assign pipe3_io_length_in_1 = pipe2_io_length_out_1; // @[executor.scala 509:26]
  assign pipe3_io_length_in_2 = pipe2_io_length_out_2; // @[executor.scala 509:26]
  assign pipe3_io_length_in_3 = pipe2_io_length_out_3; // @[executor.scala 509:26]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_160 = pipe3_io_pipe_phv_out_data_160; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_161 = pipe3_io_pipe_phv_out_data_161; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_162 = pipe3_io_pipe_phv_out_data_162; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_163 = pipe3_io_pipe_phv_out_data_163; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_164 = pipe3_io_pipe_phv_out_data_164; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_165 = pipe3_io_pipe_phv_out_data_165; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_166 = pipe3_io_pipe_phv_out_data_166; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_167 = pipe3_io_pipe_phv_out_data_167; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_168 = pipe3_io_pipe_phv_out_data_168; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_169 = pipe3_io_pipe_phv_out_data_169; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_170 = pipe3_io_pipe_phv_out_data_170; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_171 = pipe3_io_pipe_phv_out_data_171; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_172 = pipe3_io_pipe_phv_out_data_172; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_173 = pipe3_io_pipe_phv_out_data_173; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_174 = pipe3_io_pipe_phv_out_data_174; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_175 = pipe3_io_pipe_phv_out_data_175; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_176 = pipe3_io_pipe_phv_out_data_176; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_177 = pipe3_io_pipe_phv_out_data_177; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_178 = pipe3_io_pipe_phv_out_data_178; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_179 = pipe3_io_pipe_phv_out_data_179; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_180 = pipe3_io_pipe_phv_out_data_180; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_181 = pipe3_io_pipe_phv_out_data_181; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_182 = pipe3_io_pipe_phv_out_data_182; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_183 = pipe3_io_pipe_phv_out_data_183; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_184 = pipe3_io_pipe_phv_out_data_184; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_185 = pipe3_io_pipe_phv_out_data_185; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_186 = pipe3_io_pipe_phv_out_data_186; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_187 = pipe3_io_pipe_phv_out_data_187; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_188 = pipe3_io_pipe_phv_out_data_188; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_189 = pipe3_io_pipe_phv_out_data_189; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_190 = pipe3_io_pipe_phv_out_data_190; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_191 = pipe3_io_pipe_phv_out_data_191; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_192 = pipe3_io_pipe_phv_out_data_192; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_193 = pipe3_io_pipe_phv_out_data_193; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_194 = pipe3_io_pipe_phv_out_data_194; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_195 = pipe3_io_pipe_phv_out_data_195; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_196 = pipe3_io_pipe_phv_out_data_196; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_197 = pipe3_io_pipe_phv_out_data_197; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_198 = pipe3_io_pipe_phv_out_data_198; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_199 = pipe3_io_pipe_phv_out_data_199; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_200 = pipe3_io_pipe_phv_out_data_200; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_201 = pipe3_io_pipe_phv_out_data_201; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_202 = pipe3_io_pipe_phv_out_data_202; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_203 = pipe3_io_pipe_phv_out_data_203; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_204 = pipe3_io_pipe_phv_out_data_204; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_205 = pipe3_io_pipe_phv_out_data_205; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_206 = pipe3_io_pipe_phv_out_data_206; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_207 = pipe3_io_pipe_phv_out_data_207; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_208 = pipe3_io_pipe_phv_out_data_208; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_209 = pipe3_io_pipe_phv_out_data_209; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_210 = pipe3_io_pipe_phv_out_data_210; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_211 = pipe3_io_pipe_phv_out_data_211; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_212 = pipe3_io_pipe_phv_out_data_212; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_213 = pipe3_io_pipe_phv_out_data_213; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_214 = pipe3_io_pipe_phv_out_data_214; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_215 = pipe3_io_pipe_phv_out_data_215; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_216 = pipe3_io_pipe_phv_out_data_216; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_217 = pipe3_io_pipe_phv_out_data_217; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_218 = pipe3_io_pipe_phv_out_data_218; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_219 = pipe3_io_pipe_phv_out_data_219; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_220 = pipe3_io_pipe_phv_out_data_220; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_221 = pipe3_io_pipe_phv_out_data_221; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_222 = pipe3_io_pipe_phv_out_data_222; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_223 = pipe3_io_pipe_phv_out_data_223; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_224 = pipe3_io_pipe_phv_out_data_224; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_225 = pipe3_io_pipe_phv_out_data_225; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_226 = pipe3_io_pipe_phv_out_data_226; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_227 = pipe3_io_pipe_phv_out_data_227; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_228 = pipe3_io_pipe_phv_out_data_228; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_229 = pipe3_io_pipe_phv_out_data_229; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_230 = pipe3_io_pipe_phv_out_data_230; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_231 = pipe3_io_pipe_phv_out_data_231; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_232 = pipe3_io_pipe_phv_out_data_232; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_233 = pipe3_io_pipe_phv_out_data_233; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_234 = pipe3_io_pipe_phv_out_data_234; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_235 = pipe3_io_pipe_phv_out_data_235; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_236 = pipe3_io_pipe_phv_out_data_236; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_237 = pipe3_io_pipe_phv_out_data_237; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_238 = pipe3_io_pipe_phv_out_data_238; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_239 = pipe3_io_pipe_phv_out_data_239; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_240 = pipe3_io_pipe_phv_out_data_240; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_241 = pipe3_io_pipe_phv_out_data_241; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_242 = pipe3_io_pipe_phv_out_data_242; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_243 = pipe3_io_pipe_phv_out_data_243; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_244 = pipe3_io_pipe_phv_out_data_244; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_245 = pipe3_io_pipe_phv_out_data_245; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_246 = pipe3_io_pipe_phv_out_data_246; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_247 = pipe3_io_pipe_phv_out_data_247; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_248 = pipe3_io_pipe_phv_out_data_248; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_249 = pipe3_io_pipe_phv_out_data_249; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_250 = pipe3_io_pipe_phv_out_data_250; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_251 = pipe3_io_pipe_phv_out_data_251; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_252 = pipe3_io_pipe_phv_out_data_252; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_253 = pipe3_io_pipe_phv_out_data_253; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_254 = pipe3_io_pipe_phv_out_data_254; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_255 = pipe3_io_pipe_phv_out_data_255; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[executor.scala 511:27]
  assign pipe4_io_vliw_in_0 = pipe3_io_vliw_out_0; // @[executor.scala 512:27]
  assign pipe4_io_vliw_in_1 = pipe3_io_vliw_out_1; // @[executor.scala 512:27]
  assign pipe4_io_vliw_in_2 = pipe3_io_vliw_out_2; // @[executor.scala 512:27]
  assign pipe4_io_vliw_in_3 = pipe3_io_vliw_out_3; // @[executor.scala 512:27]
  assign pipe4_io_field_in_0 = pipe3_io_field_out_0; // @[executor.scala 513:27]
  assign pipe4_io_field_in_1 = pipe3_io_field_out_1; // @[executor.scala 513:27]
  assign pipe4_io_field_in_2 = pipe3_io_field_out_2; // @[executor.scala 513:27]
  assign pipe4_io_field_in_3 = pipe3_io_field_out_3; // @[executor.scala 513:27]
  assign pipe4_io_mask_in_0 = pipe3_io_mask_out_0; // @[executor.scala 514:27]
  assign pipe4_io_mask_in_1 = pipe3_io_mask_out_1; // @[executor.scala 514:27]
  assign pipe4_io_mask_in_2 = pipe3_io_mask_out_2; // @[executor.scala 514:27]
  assign pipe4_io_mask_in_3 = pipe3_io_mask_out_3; // @[executor.scala 514:27]
  assign pipe4_io_bias_in_0 = pipe3_io_bias_out_0; // @[executor.scala 515:27]
  assign pipe4_io_bias_in_1 = pipe3_io_bias_out_1; // @[executor.scala 515:27]
  assign pipe4_io_bias_in_2 = pipe3_io_bias_out_2; // @[executor.scala 515:27]
  assign pipe4_io_bias_in_3 = pipe3_io_bias_out_3; // @[executor.scala 515:27]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_96 = pipe4_io_pipe_phv_out_data_96; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_97 = pipe4_io_pipe_phv_out_data_97; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_98 = pipe4_io_pipe_phv_out_data_98; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_99 = pipe4_io_pipe_phv_out_data_99; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_100 = pipe4_io_pipe_phv_out_data_100; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_101 = pipe4_io_pipe_phv_out_data_101; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_102 = pipe4_io_pipe_phv_out_data_102; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_103 = pipe4_io_pipe_phv_out_data_103; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_104 = pipe4_io_pipe_phv_out_data_104; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_105 = pipe4_io_pipe_phv_out_data_105; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_106 = pipe4_io_pipe_phv_out_data_106; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_107 = pipe4_io_pipe_phv_out_data_107; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_108 = pipe4_io_pipe_phv_out_data_108; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_109 = pipe4_io_pipe_phv_out_data_109; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_110 = pipe4_io_pipe_phv_out_data_110; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_111 = pipe4_io_pipe_phv_out_data_111; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_112 = pipe4_io_pipe_phv_out_data_112; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_113 = pipe4_io_pipe_phv_out_data_113; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_114 = pipe4_io_pipe_phv_out_data_114; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_115 = pipe4_io_pipe_phv_out_data_115; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_116 = pipe4_io_pipe_phv_out_data_116; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_117 = pipe4_io_pipe_phv_out_data_117; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_118 = pipe4_io_pipe_phv_out_data_118; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_119 = pipe4_io_pipe_phv_out_data_119; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_120 = pipe4_io_pipe_phv_out_data_120; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_121 = pipe4_io_pipe_phv_out_data_121; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_122 = pipe4_io_pipe_phv_out_data_122; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_123 = pipe4_io_pipe_phv_out_data_123; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_124 = pipe4_io_pipe_phv_out_data_124; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_125 = pipe4_io_pipe_phv_out_data_125; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_126 = pipe4_io_pipe_phv_out_data_126; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_127 = pipe4_io_pipe_phv_out_data_127; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_128 = pipe4_io_pipe_phv_out_data_128; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_129 = pipe4_io_pipe_phv_out_data_129; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_130 = pipe4_io_pipe_phv_out_data_130; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_131 = pipe4_io_pipe_phv_out_data_131; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_132 = pipe4_io_pipe_phv_out_data_132; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_133 = pipe4_io_pipe_phv_out_data_133; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_134 = pipe4_io_pipe_phv_out_data_134; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_135 = pipe4_io_pipe_phv_out_data_135; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_136 = pipe4_io_pipe_phv_out_data_136; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_137 = pipe4_io_pipe_phv_out_data_137; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_138 = pipe4_io_pipe_phv_out_data_138; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_139 = pipe4_io_pipe_phv_out_data_139; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_140 = pipe4_io_pipe_phv_out_data_140; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_141 = pipe4_io_pipe_phv_out_data_141; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_142 = pipe4_io_pipe_phv_out_data_142; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_143 = pipe4_io_pipe_phv_out_data_143; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_144 = pipe4_io_pipe_phv_out_data_144; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_145 = pipe4_io_pipe_phv_out_data_145; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_146 = pipe4_io_pipe_phv_out_data_146; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_147 = pipe4_io_pipe_phv_out_data_147; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_148 = pipe4_io_pipe_phv_out_data_148; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_149 = pipe4_io_pipe_phv_out_data_149; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_150 = pipe4_io_pipe_phv_out_data_150; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_151 = pipe4_io_pipe_phv_out_data_151; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_152 = pipe4_io_pipe_phv_out_data_152; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_153 = pipe4_io_pipe_phv_out_data_153; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_154 = pipe4_io_pipe_phv_out_data_154; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_155 = pipe4_io_pipe_phv_out_data_155; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_156 = pipe4_io_pipe_phv_out_data_156; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_157 = pipe4_io_pipe_phv_out_data_157; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_158 = pipe4_io_pipe_phv_out_data_158; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_159 = pipe4_io_pipe_phv_out_data_159; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_160 = pipe4_io_pipe_phv_out_data_160; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_161 = pipe4_io_pipe_phv_out_data_161; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_162 = pipe4_io_pipe_phv_out_data_162; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_163 = pipe4_io_pipe_phv_out_data_163; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_164 = pipe4_io_pipe_phv_out_data_164; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_165 = pipe4_io_pipe_phv_out_data_165; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_166 = pipe4_io_pipe_phv_out_data_166; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_167 = pipe4_io_pipe_phv_out_data_167; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_168 = pipe4_io_pipe_phv_out_data_168; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_169 = pipe4_io_pipe_phv_out_data_169; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_170 = pipe4_io_pipe_phv_out_data_170; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_171 = pipe4_io_pipe_phv_out_data_171; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_172 = pipe4_io_pipe_phv_out_data_172; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_173 = pipe4_io_pipe_phv_out_data_173; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_174 = pipe4_io_pipe_phv_out_data_174; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_175 = pipe4_io_pipe_phv_out_data_175; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_176 = pipe4_io_pipe_phv_out_data_176; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_177 = pipe4_io_pipe_phv_out_data_177; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_178 = pipe4_io_pipe_phv_out_data_178; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_179 = pipe4_io_pipe_phv_out_data_179; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_180 = pipe4_io_pipe_phv_out_data_180; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_181 = pipe4_io_pipe_phv_out_data_181; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_182 = pipe4_io_pipe_phv_out_data_182; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_183 = pipe4_io_pipe_phv_out_data_183; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_184 = pipe4_io_pipe_phv_out_data_184; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_185 = pipe4_io_pipe_phv_out_data_185; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_186 = pipe4_io_pipe_phv_out_data_186; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_187 = pipe4_io_pipe_phv_out_data_187; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_188 = pipe4_io_pipe_phv_out_data_188; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_189 = pipe4_io_pipe_phv_out_data_189; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_190 = pipe4_io_pipe_phv_out_data_190; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_191 = pipe4_io_pipe_phv_out_data_191; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_192 = pipe4_io_pipe_phv_out_data_192; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_193 = pipe4_io_pipe_phv_out_data_193; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_194 = pipe4_io_pipe_phv_out_data_194; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_195 = pipe4_io_pipe_phv_out_data_195; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_196 = pipe4_io_pipe_phv_out_data_196; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_197 = pipe4_io_pipe_phv_out_data_197; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_198 = pipe4_io_pipe_phv_out_data_198; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_199 = pipe4_io_pipe_phv_out_data_199; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_200 = pipe4_io_pipe_phv_out_data_200; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_201 = pipe4_io_pipe_phv_out_data_201; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_202 = pipe4_io_pipe_phv_out_data_202; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_203 = pipe4_io_pipe_phv_out_data_203; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_204 = pipe4_io_pipe_phv_out_data_204; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_205 = pipe4_io_pipe_phv_out_data_205; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_206 = pipe4_io_pipe_phv_out_data_206; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_207 = pipe4_io_pipe_phv_out_data_207; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_208 = pipe4_io_pipe_phv_out_data_208; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_209 = pipe4_io_pipe_phv_out_data_209; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_210 = pipe4_io_pipe_phv_out_data_210; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_211 = pipe4_io_pipe_phv_out_data_211; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_212 = pipe4_io_pipe_phv_out_data_212; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_213 = pipe4_io_pipe_phv_out_data_213; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_214 = pipe4_io_pipe_phv_out_data_214; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_215 = pipe4_io_pipe_phv_out_data_215; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_216 = pipe4_io_pipe_phv_out_data_216; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_217 = pipe4_io_pipe_phv_out_data_217; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_218 = pipe4_io_pipe_phv_out_data_218; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_219 = pipe4_io_pipe_phv_out_data_219; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_220 = pipe4_io_pipe_phv_out_data_220; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_221 = pipe4_io_pipe_phv_out_data_221; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_222 = pipe4_io_pipe_phv_out_data_222; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_223 = pipe4_io_pipe_phv_out_data_223; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_224 = pipe4_io_pipe_phv_out_data_224; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_225 = pipe4_io_pipe_phv_out_data_225; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_226 = pipe4_io_pipe_phv_out_data_226; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_227 = pipe4_io_pipe_phv_out_data_227; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_228 = pipe4_io_pipe_phv_out_data_228; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_229 = pipe4_io_pipe_phv_out_data_229; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_230 = pipe4_io_pipe_phv_out_data_230; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_231 = pipe4_io_pipe_phv_out_data_231; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_232 = pipe4_io_pipe_phv_out_data_232; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_233 = pipe4_io_pipe_phv_out_data_233; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_234 = pipe4_io_pipe_phv_out_data_234; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_235 = pipe4_io_pipe_phv_out_data_235; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_236 = pipe4_io_pipe_phv_out_data_236; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_237 = pipe4_io_pipe_phv_out_data_237; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_238 = pipe4_io_pipe_phv_out_data_238; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_239 = pipe4_io_pipe_phv_out_data_239; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_240 = pipe4_io_pipe_phv_out_data_240; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_241 = pipe4_io_pipe_phv_out_data_241; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_242 = pipe4_io_pipe_phv_out_data_242; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_243 = pipe4_io_pipe_phv_out_data_243; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_244 = pipe4_io_pipe_phv_out_data_244; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_245 = pipe4_io_pipe_phv_out_data_245; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_246 = pipe4_io_pipe_phv_out_data_246; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_247 = pipe4_io_pipe_phv_out_data_247; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_248 = pipe4_io_pipe_phv_out_data_248; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_249 = pipe4_io_pipe_phv_out_data_249; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_250 = pipe4_io_pipe_phv_out_data_250; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_251 = pipe4_io_pipe_phv_out_data_251; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_252 = pipe4_io_pipe_phv_out_data_252; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_253 = pipe4_io_pipe_phv_out_data_253; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_254 = pipe4_io_pipe_phv_out_data_254; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_255 = pipe4_io_pipe_phv_out_data_255; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[executor.scala 517:26]
  assign pipe5_io_vliw_in_0 = pipe4_io_vliw_out_0; // @[executor.scala 518:26]
  assign pipe5_io_vliw_in_1 = pipe4_io_vliw_out_1; // @[executor.scala 518:26]
  assign pipe5_io_vliw_in_2 = pipe4_io_vliw_out_2; // @[executor.scala 518:26]
  assign pipe5_io_vliw_in_3 = pipe4_io_vliw_out_3; // @[executor.scala 518:26]
  assign pipe5_io_field_in_0 = pipe4_io_field_out_0; // @[executor.scala 519:26]
  assign pipe5_io_field_in_1 = pipe4_io_field_out_1; // @[executor.scala 519:26]
  assign pipe5_io_field_in_2 = pipe4_io_field_out_2; // @[executor.scala 519:26]
  assign pipe5_io_field_in_3 = pipe4_io_field_out_3; // @[executor.scala 519:26]
  assign pipe5_io_mask_in_0 = pipe4_io_mask_out_0; // @[executor.scala 520:26]
  assign pipe5_io_mask_in_1 = pipe4_io_mask_out_1; // @[executor.scala 520:26]
  assign pipe5_io_mask_in_2 = pipe4_io_mask_out_2; // @[executor.scala 520:26]
  assign pipe5_io_mask_in_3 = pipe4_io_mask_out_3; // @[executor.scala 520:26]
  assign pipe5_io_bias_in_0 = pipe4_io_bias_out_0; // @[executor.scala 521:26]
  assign pipe5_io_bias_in_1 = pipe4_io_bias_out_1; // @[executor.scala 521:26]
  assign pipe5_io_bias_in_2 = pipe4_io_bias_out_2; // @[executor.scala 521:26]
  assign pipe5_io_bias_in_3 = pipe4_io_bias_out_3; // @[executor.scala 521:26]
  assign pipe5_io_dst_offset_in_0 = pipe4_io_dst_offset_out_0; // @[executor.scala 522:28]
  assign pipe5_io_dst_offset_in_1 = pipe4_io_dst_offset_out_1; // @[executor.scala 522:28]
  assign pipe5_io_dst_offset_in_2 = pipe4_io_dst_offset_out_2; // @[executor.scala 522:28]
  assign pipe5_io_dst_offset_in_3 = pipe4_io_dst_offset_out_3; // @[executor.scala 522:28]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_96 = pipe5_io_pipe_phv_out_data_96; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_97 = pipe5_io_pipe_phv_out_data_97; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_98 = pipe5_io_pipe_phv_out_data_98; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_99 = pipe5_io_pipe_phv_out_data_99; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_100 = pipe5_io_pipe_phv_out_data_100; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_101 = pipe5_io_pipe_phv_out_data_101; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_102 = pipe5_io_pipe_phv_out_data_102; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_103 = pipe5_io_pipe_phv_out_data_103; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_104 = pipe5_io_pipe_phv_out_data_104; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_105 = pipe5_io_pipe_phv_out_data_105; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_106 = pipe5_io_pipe_phv_out_data_106; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_107 = pipe5_io_pipe_phv_out_data_107; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_108 = pipe5_io_pipe_phv_out_data_108; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_109 = pipe5_io_pipe_phv_out_data_109; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_110 = pipe5_io_pipe_phv_out_data_110; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_111 = pipe5_io_pipe_phv_out_data_111; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_112 = pipe5_io_pipe_phv_out_data_112; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_113 = pipe5_io_pipe_phv_out_data_113; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_114 = pipe5_io_pipe_phv_out_data_114; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_115 = pipe5_io_pipe_phv_out_data_115; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_116 = pipe5_io_pipe_phv_out_data_116; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_117 = pipe5_io_pipe_phv_out_data_117; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_118 = pipe5_io_pipe_phv_out_data_118; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_119 = pipe5_io_pipe_phv_out_data_119; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_120 = pipe5_io_pipe_phv_out_data_120; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_121 = pipe5_io_pipe_phv_out_data_121; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_122 = pipe5_io_pipe_phv_out_data_122; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_123 = pipe5_io_pipe_phv_out_data_123; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_124 = pipe5_io_pipe_phv_out_data_124; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_125 = pipe5_io_pipe_phv_out_data_125; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_126 = pipe5_io_pipe_phv_out_data_126; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_127 = pipe5_io_pipe_phv_out_data_127; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_128 = pipe5_io_pipe_phv_out_data_128; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_129 = pipe5_io_pipe_phv_out_data_129; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_130 = pipe5_io_pipe_phv_out_data_130; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_131 = pipe5_io_pipe_phv_out_data_131; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_132 = pipe5_io_pipe_phv_out_data_132; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_133 = pipe5_io_pipe_phv_out_data_133; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_134 = pipe5_io_pipe_phv_out_data_134; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_135 = pipe5_io_pipe_phv_out_data_135; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_136 = pipe5_io_pipe_phv_out_data_136; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_137 = pipe5_io_pipe_phv_out_data_137; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_138 = pipe5_io_pipe_phv_out_data_138; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_139 = pipe5_io_pipe_phv_out_data_139; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_140 = pipe5_io_pipe_phv_out_data_140; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_141 = pipe5_io_pipe_phv_out_data_141; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_142 = pipe5_io_pipe_phv_out_data_142; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_143 = pipe5_io_pipe_phv_out_data_143; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_144 = pipe5_io_pipe_phv_out_data_144; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_145 = pipe5_io_pipe_phv_out_data_145; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_146 = pipe5_io_pipe_phv_out_data_146; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_147 = pipe5_io_pipe_phv_out_data_147; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_148 = pipe5_io_pipe_phv_out_data_148; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_149 = pipe5_io_pipe_phv_out_data_149; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_150 = pipe5_io_pipe_phv_out_data_150; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_151 = pipe5_io_pipe_phv_out_data_151; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_152 = pipe5_io_pipe_phv_out_data_152; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_153 = pipe5_io_pipe_phv_out_data_153; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_154 = pipe5_io_pipe_phv_out_data_154; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_155 = pipe5_io_pipe_phv_out_data_155; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_156 = pipe5_io_pipe_phv_out_data_156; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_157 = pipe5_io_pipe_phv_out_data_157; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_158 = pipe5_io_pipe_phv_out_data_158; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_159 = pipe5_io_pipe_phv_out_data_159; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_160 = pipe5_io_pipe_phv_out_data_160; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_161 = pipe5_io_pipe_phv_out_data_161; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_162 = pipe5_io_pipe_phv_out_data_162; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_163 = pipe5_io_pipe_phv_out_data_163; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_164 = pipe5_io_pipe_phv_out_data_164; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_165 = pipe5_io_pipe_phv_out_data_165; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_166 = pipe5_io_pipe_phv_out_data_166; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_167 = pipe5_io_pipe_phv_out_data_167; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_168 = pipe5_io_pipe_phv_out_data_168; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_169 = pipe5_io_pipe_phv_out_data_169; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_170 = pipe5_io_pipe_phv_out_data_170; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_171 = pipe5_io_pipe_phv_out_data_171; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_172 = pipe5_io_pipe_phv_out_data_172; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_173 = pipe5_io_pipe_phv_out_data_173; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_174 = pipe5_io_pipe_phv_out_data_174; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_175 = pipe5_io_pipe_phv_out_data_175; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_176 = pipe5_io_pipe_phv_out_data_176; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_177 = pipe5_io_pipe_phv_out_data_177; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_178 = pipe5_io_pipe_phv_out_data_178; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_179 = pipe5_io_pipe_phv_out_data_179; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_180 = pipe5_io_pipe_phv_out_data_180; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_181 = pipe5_io_pipe_phv_out_data_181; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_182 = pipe5_io_pipe_phv_out_data_182; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_183 = pipe5_io_pipe_phv_out_data_183; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_184 = pipe5_io_pipe_phv_out_data_184; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_185 = pipe5_io_pipe_phv_out_data_185; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_186 = pipe5_io_pipe_phv_out_data_186; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_187 = pipe5_io_pipe_phv_out_data_187; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_188 = pipe5_io_pipe_phv_out_data_188; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_189 = pipe5_io_pipe_phv_out_data_189; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_190 = pipe5_io_pipe_phv_out_data_190; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_191 = pipe5_io_pipe_phv_out_data_191; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_192 = pipe5_io_pipe_phv_out_data_192; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_193 = pipe5_io_pipe_phv_out_data_193; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_194 = pipe5_io_pipe_phv_out_data_194; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_195 = pipe5_io_pipe_phv_out_data_195; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_196 = pipe5_io_pipe_phv_out_data_196; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_197 = pipe5_io_pipe_phv_out_data_197; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_198 = pipe5_io_pipe_phv_out_data_198; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_199 = pipe5_io_pipe_phv_out_data_199; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_200 = pipe5_io_pipe_phv_out_data_200; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_201 = pipe5_io_pipe_phv_out_data_201; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_202 = pipe5_io_pipe_phv_out_data_202; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_203 = pipe5_io_pipe_phv_out_data_203; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_204 = pipe5_io_pipe_phv_out_data_204; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_205 = pipe5_io_pipe_phv_out_data_205; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_206 = pipe5_io_pipe_phv_out_data_206; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_207 = pipe5_io_pipe_phv_out_data_207; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_208 = pipe5_io_pipe_phv_out_data_208; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_209 = pipe5_io_pipe_phv_out_data_209; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_210 = pipe5_io_pipe_phv_out_data_210; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_211 = pipe5_io_pipe_phv_out_data_211; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_212 = pipe5_io_pipe_phv_out_data_212; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_213 = pipe5_io_pipe_phv_out_data_213; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_214 = pipe5_io_pipe_phv_out_data_214; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_215 = pipe5_io_pipe_phv_out_data_215; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_216 = pipe5_io_pipe_phv_out_data_216; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_217 = pipe5_io_pipe_phv_out_data_217; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_218 = pipe5_io_pipe_phv_out_data_218; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_219 = pipe5_io_pipe_phv_out_data_219; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_220 = pipe5_io_pipe_phv_out_data_220; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_221 = pipe5_io_pipe_phv_out_data_221; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_222 = pipe5_io_pipe_phv_out_data_222; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_223 = pipe5_io_pipe_phv_out_data_223; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_224 = pipe5_io_pipe_phv_out_data_224; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_225 = pipe5_io_pipe_phv_out_data_225; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_226 = pipe5_io_pipe_phv_out_data_226; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_227 = pipe5_io_pipe_phv_out_data_227; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_228 = pipe5_io_pipe_phv_out_data_228; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_229 = pipe5_io_pipe_phv_out_data_229; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_230 = pipe5_io_pipe_phv_out_data_230; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_231 = pipe5_io_pipe_phv_out_data_231; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_232 = pipe5_io_pipe_phv_out_data_232; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_233 = pipe5_io_pipe_phv_out_data_233; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_234 = pipe5_io_pipe_phv_out_data_234; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_235 = pipe5_io_pipe_phv_out_data_235; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_236 = pipe5_io_pipe_phv_out_data_236; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_237 = pipe5_io_pipe_phv_out_data_237; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_238 = pipe5_io_pipe_phv_out_data_238; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_239 = pipe5_io_pipe_phv_out_data_239; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_240 = pipe5_io_pipe_phv_out_data_240; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_241 = pipe5_io_pipe_phv_out_data_241; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_242 = pipe5_io_pipe_phv_out_data_242; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_243 = pipe5_io_pipe_phv_out_data_243; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_244 = pipe5_io_pipe_phv_out_data_244; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_245 = pipe5_io_pipe_phv_out_data_245; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_246 = pipe5_io_pipe_phv_out_data_246; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_247 = pipe5_io_pipe_phv_out_data_247; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_248 = pipe5_io_pipe_phv_out_data_248; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_249 = pipe5_io_pipe_phv_out_data_249; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_250 = pipe5_io_pipe_phv_out_data_250; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_251 = pipe5_io_pipe_phv_out_data_251; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_252 = pipe5_io_pipe_phv_out_data_252; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_253 = pipe5_io_pipe_phv_out_data_253; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_254 = pipe5_io_pipe_phv_out_data_254; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_255 = pipe5_io_pipe_phv_out_data_255; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[executor.scala 524:26]
  assign pipe6_io_vliw_in_0 = pipe5_io_vliw_out_0; // @[executor.scala 525:26]
  assign pipe6_io_vliw_in_1 = pipe5_io_vliw_out_1; // @[executor.scala 525:26]
  assign pipe6_io_vliw_in_2 = pipe5_io_vliw_out_2; // @[executor.scala 525:26]
  assign pipe6_io_vliw_in_3 = pipe5_io_vliw_out_3; // @[executor.scala 525:26]
  assign pipe6_io_field_in_0 = pipe5_io_field_out_0; // @[executor.scala 526:26]
  assign pipe6_io_field_in_1 = pipe5_io_field_out_1; // @[executor.scala 526:26]
  assign pipe6_io_field_in_2 = pipe5_io_field_out_2; // @[executor.scala 526:26]
  assign pipe6_io_field_in_3 = pipe5_io_field_out_3; // @[executor.scala 526:26]
  assign pipe6_io_mask_in_0 = pipe5_io_mask_out_0; // @[executor.scala 527:26]
  assign pipe6_io_mask_in_1 = pipe5_io_mask_out_1; // @[executor.scala 527:26]
  assign pipe6_io_mask_in_2 = pipe5_io_mask_out_2; // @[executor.scala 527:26]
  assign pipe6_io_mask_in_3 = pipe5_io_mask_out_3; // @[executor.scala 527:26]
  assign pipe6_io_dst_offset_in_0 = pipe5_io_dst_offset_out_0; // @[executor.scala 528:28]
  assign pipe6_io_dst_offset_in_1 = pipe5_io_dst_offset_out_1; // @[executor.scala 528:28]
  assign pipe6_io_dst_offset_in_2 = pipe5_io_dst_offset_out_2; // @[executor.scala 528:28]
  assign pipe6_io_dst_offset_in_3 = pipe5_io_dst_offset_out_3; // @[executor.scala 528:28]
endmodule
