module PrimitiveWriteBackPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [14:0] io_nid_in,
  input  [1:0]  io_tag_in_0,
  input  [1:0]  io_tag_in_1,
  input  [1:0]  io_tag_in_2,
  input  [1:0]  io_tag_in_3,
  input  [1:0]  io_tag_in_4,
  input  [1:0]  io_tag_in_5,
  input  [1:0]  io_tag_in_6,
  input  [1:0]  io_tag_in_7,
  input  [1:0]  io_tag_in_8,
  input  [1:0]  io_tag_in_9,
  input  [1:0]  io_tag_in_10,
  input  [1:0]  io_tag_in_11,
  input  [1:0]  io_tag_in_12,
  input  [1:0]  io_tag_in_13,
  input  [1:0]  io_tag_in_14,
  input  [1:0]  io_tag_in_15,
  input  [1:0]  io_tag_in_16,
  input  [1:0]  io_tag_in_17,
  input  [1:0]  io_tag_in_18,
  input  [1:0]  io_tag_in_19,
  input  [1:0]  io_tag_in_20,
  input  [1:0]  io_tag_in_21,
  input  [1:0]  io_tag_in_22,
  input  [1:0]  io_tag_in_23,
  input  [1:0]  io_tag_in_24,
  input  [1:0]  io_tag_in_25,
  input  [1:0]  io_tag_in_26,
  input  [1:0]  io_tag_in_27,
  input  [1:0]  io_tag_in_28,
  input  [1:0]  io_tag_in_29,
  input  [1:0]  io_tag_in_30,
  input  [1:0]  io_tag_in_31,
  input  [1:0]  io_tag_in_32,
  input  [1:0]  io_tag_in_33,
  input  [1:0]  io_tag_in_34,
  input  [1:0]  io_tag_in_35,
  input  [1:0]  io_tag_in_36,
  input  [1:0]  io_tag_in_37,
  input  [1:0]  io_tag_in_38,
  input  [1:0]  io_tag_in_39,
  input  [1:0]  io_tag_in_40,
  input  [1:0]  io_tag_in_41,
  input  [1:0]  io_tag_in_42,
  input  [1:0]  io_tag_in_43,
  input  [1:0]  io_tag_in_44,
  input  [1:0]  io_tag_in_45,
  input  [1:0]  io_tag_in_46,
  input  [1:0]  io_tag_in_47,
  input  [1:0]  io_tag_in_48,
  input  [1:0]  io_tag_in_49,
  input  [1:0]  io_tag_in_50,
  input  [1:0]  io_tag_in_51,
  input  [1:0]  io_tag_in_52,
  input  [1:0]  io_tag_in_53,
  input  [1:0]  io_tag_in_54,
  input  [1:0]  io_tag_in_55,
  input  [1:0]  io_tag_in_56,
  input  [1:0]  io_tag_in_57,
  input  [1:0]  io_tag_in_58,
  input  [1:0]  io_tag_in_59,
  input  [1:0]  io_tag_in_60,
  input  [1:0]  io_tag_in_61,
  input  [1:0]  io_tag_in_62,
  input  [1:0]  io_tag_in_63,
  input  [1:0]  io_tag_in_64,
  input  [1:0]  io_tag_in_65,
  input  [1:0]  io_tag_in_66,
  input  [1:0]  io_tag_in_67,
  input  [1:0]  io_tag_in_68,
  input  [1:0]  io_tag_in_69,
  input  [7:0]  io_field_set_field8_0,
  input  [7:0]  io_field_set_field8_1,
  input  [7:0]  io_field_set_field8_2,
  input  [7:0]  io_field_set_field8_3,
  input  [7:0]  io_field_set_field8_4,
  input  [7:0]  io_field_set_field8_5,
  input  [7:0]  io_field_set_field8_6,
  input  [7:0]  io_field_set_field8_7,
  input  [7:0]  io_field_set_field8_8,
  input  [7:0]  io_field_set_field8_9,
  input  [7:0]  io_field_set_field8_10,
  input  [7:0]  io_field_set_field8_11,
  input  [7:0]  io_field_set_field8_12,
  input  [7:0]  io_field_set_field8_13,
  input  [7:0]  io_field_set_field8_14,
  input  [7:0]  io_field_set_field8_15,
  input  [7:0]  io_field_set_field8_16,
  input  [7:0]  io_field_set_field8_17,
  input  [7:0]  io_field_set_field8_18,
  input  [7:0]  io_field_set_field8_19,
  input  [7:0]  io_field_set_field8_20,
  input  [7:0]  io_field_set_field8_21,
  input  [7:0]  io_field_set_field8_22,
  input  [7:0]  io_field_set_field8_23,
  input  [7:0]  io_field_set_field8_24,
  input  [7:0]  io_field_set_field8_25,
  input  [7:0]  io_field_set_field8_26,
  input  [7:0]  io_field_set_field8_27,
  input  [7:0]  io_field_set_field8_28,
  input  [7:0]  io_field_set_field8_29,
  input  [7:0]  io_field_set_field8_30,
  input  [7:0]  io_field_set_field8_31,
  input  [15:0] io_field_set_field16_0,
  input  [15:0] io_field_set_field16_1,
  input  [15:0] io_field_set_field16_2,
  input  [15:0] io_field_set_field16_3,
  input  [15:0] io_field_set_field16_4,
  input  [15:0] io_field_set_field16_5,
  input  [15:0] io_field_set_field16_6,
  input  [15:0] io_field_set_field16_7,
  input  [15:0] io_field_set_field16_8,
  input  [15:0] io_field_set_field16_9,
  input  [15:0] io_field_set_field16_10,
  input  [15:0] io_field_set_field16_11,
  input  [15:0] io_field_set_field16_12,
  input  [15:0] io_field_set_field16_13,
  input  [15:0] io_field_set_field16_14,
  input  [15:0] io_field_set_field16_15,
  input  [15:0] io_field_set_field16_16,
  input  [15:0] io_field_set_field16_17,
  input  [15:0] io_field_set_field16_18,
  input  [15:0] io_field_set_field16_19,
  input  [15:0] io_field_set_field16_20,
  input  [15:0] io_field_set_field16_21,
  input  [15:0] io_field_set_field16_22,
  input  [15:0] io_field_set_field16_23,
  input  [15:0] io_field_set_field16_24,
  input  [15:0] io_field_set_field16_25,
  input  [15:0] io_field_set_field16_26,
  input  [15:0] io_field_set_field16_27,
  input  [15:0] io_field_set_field16_28,
  input  [15:0] io_field_set_field16_29,
  input  [15:0] io_field_set_field16_30,
  input  [15:0] io_field_set_field16_31,
  input  [15:0] io_field_set_field16_32,
  input  [15:0] io_field_set_field16_33,
  input  [15:0] io_field_set_field16_34,
  input  [15:0] io_field_set_field16_35,
  input  [15:0] io_field_set_field16_36,
  input  [15:0] io_field_set_field16_37
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_1; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_2; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_3; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_4; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_5; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_6; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_7; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_8; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_9; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_10; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_11; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_12; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_13; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_14; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_15; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_16; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_17; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_18; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_19; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_20; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_21; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_22; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_23; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_24; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_25; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_26; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_27; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_28; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_29; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_30; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_31; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_32; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_33; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_34; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_35; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_36; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_37; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_38; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_39; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_40; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_41; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_42; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_43; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_44; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_45; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_46; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_47; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_48; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_49; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_50; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_51; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_52; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_53; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_54; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_55; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_56; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_57; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_58; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_59; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_60; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_61; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_62; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_63; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_64; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_65; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_66; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_67; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_68; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_69; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_70; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_71; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_72; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_73; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_74; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_75; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_76; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_77; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_78; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_79; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_80; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_81; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_82; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_83; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_84; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_85; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_86; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_87; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_88; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_89; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_90; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_91; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_92; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_93; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_94; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_95; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_96; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_97; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_98; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_99; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_100; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_101; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_102; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_103; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_104; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_105; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_106; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_107; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_108; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_109; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_110; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_111; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_112; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_113; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_114; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_115; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_116; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_117; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_118; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_119; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_120; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_121; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_122; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_123; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_124; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_125; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_126; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_127; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_128; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_129; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_130; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_131; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_132; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_133; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_134; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_135; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_136; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_137; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_138; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_139; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_140; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_141; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_142; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_143; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_144; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_145; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_146; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_147; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_148; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_149; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_150; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_151; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_152; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_153; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_154; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_155; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_156; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_157; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_158; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_159; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_160; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_161; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_162; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_163; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_164; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_165; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_166; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_167; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_168; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_169; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_170; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_171; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_172; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_173; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_174; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_175; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_176; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_177; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_178; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_179; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_180; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_181; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_182; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_183; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_184; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_185; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_186; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_187; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_188; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_189; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_190; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_191; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_192; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_193; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_194; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_195; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_196; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_197; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_198; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_199; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_200; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_201; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_202; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_203; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_204; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_205; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_206; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_207; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_208; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_209; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_210; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_211; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_212; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_213; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_214; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_215; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_216; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_217; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_218; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_219; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_220; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_221; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_222; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_223; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_224; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_225; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_226; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_227; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_228; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_229; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_230; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_231; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_232; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_233; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_234; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_235; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_236; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_237; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_238; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_239; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_240; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_241; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_242; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_243; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_244; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_245; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_246; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_247; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_248; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_249; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_250; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_251; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_252; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_253; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_254; // @[executor_pisa.scala 244:22]
  reg [7:0] phv_data_255; // @[executor_pisa.scala 244:22]
  reg [3:0] phv_next_processor_id; // @[executor_pisa.scala 244:22]
  reg  phv_next_config_id; // @[executor_pisa.scala 244:22]
  reg [7:0] fs_field8_0; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_1; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_2; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_3; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_4; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_5; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_6; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_7; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_8; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_9; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_10; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_11; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_12; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_13; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_14; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_15; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_16; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_17; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_18; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_19; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_20; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_21; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_22; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_23; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_24; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_25; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_26; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_27; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_28; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_29; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_30; // @[executor_pisa.scala 248:21]
  reg [7:0] fs_field8_31; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_0; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_1; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_2; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_3; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_4; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_5; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_6; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_7; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_8; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_9; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_10; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_11; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_12; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_13; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_14; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_15; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_16; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_17; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_18; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_19; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_20; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_21; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_22; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_23; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_24; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_25; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_26; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_27; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_28; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_29; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_30; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_31; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_32; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_33; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_34; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_35; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_36; // @[executor_pisa.scala 248:21]
  reg [15:0] fs_field16_37; // @[executor_pisa.scala 248:21]
  reg [1:0] tag_0; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_1; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_2; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_3; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_4; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_5; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_6; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_7; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_8; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_9; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_10; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_11; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_12; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_13; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_14; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_15; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_16; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_17; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_18; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_19; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_20; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_21; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_22; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_23; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_24; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_25; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_26; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_27; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_28; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_29; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_30; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_31; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_32; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_33; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_34; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_35; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_36; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_37; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_38; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_39; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_40; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_41; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_42; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_43; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_44; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_45; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_46; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_47; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_48; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_49; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_50; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_51; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_52; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_53; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_54; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_55; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_56; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_57; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_58; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_59; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_60; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_61; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_62; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_63; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_64; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_65; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_66; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_67; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_68; // @[executor_pisa.scala 251:22]
  reg [1:0] tag_69; // @[executor_pisa.scala 251:22]
  reg [14:0] nid; // @[executor_pisa.scala 254:22]
  wire  _add1_T_2 = tag_0[0] ^ tag_0[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1 = _add1_T_2 ? fs_field8_0 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T = tag_0 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2 = _add2_T ? 8'h0 : phv_data_0; // @[executor_pisa.scala 268:24]
  wire  _add1_T_6 = tag_1[0] ^ tag_1[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_1 = _add1_T_6 ? fs_field8_1 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_2 = tag_1 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_1 = _add2_T_2 ? 8'h0 : phv_data_1; // @[executor_pisa.scala 268:24]
  wire  _add1_T_10 = tag_2[0] ^ tag_2[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_2 = _add1_T_10 ? fs_field8_2 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_4 = tag_2 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_2 = _add2_T_4 ? 8'h0 : phv_data_2; // @[executor_pisa.scala 268:24]
  wire  _add1_T_14 = tag_3[0] ^ tag_3[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_3 = _add1_T_14 ? fs_field8_3 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_6 = tag_3 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_3 = _add2_T_6 ? 8'h0 : phv_data_3; // @[executor_pisa.scala 268:24]
  wire  _add1_T_18 = tag_4[0] ^ tag_4[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_4 = _add1_T_18 ? fs_field8_4 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_8 = tag_4 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_4 = _add2_T_8 ? 8'h0 : phv_data_4; // @[executor_pisa.scala 268:24]
  wire  _add1_T_22 = tag_5[0] ^ tag_5[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_5 = _add1_T_22 ? fs_field8_5 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_10 = tag_5 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_5 = _add2_T_10 ? 8'h0 : phv_data_5; // @[executor_pisa.scala 268:24]
  wire  _add1_T_26 = tag_6[0] ^ tag_6[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_6 = _add1_T_26 ? fs_field8_6 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_12 = tag_6 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_6 = _add2_T_12 ? 8'h0 : phv_data_6; // @[executor_pisa.scala 268:24]
  wire  _add1_T_30 = tag_7[0] ^ tag_7[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_7 = _add1_T_30 ? fs_field8_7 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_14 = tag_7 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_7 = _add2_T_14 ? 8'h0 : phv_data_7; // @[executor_pisa.scala 268:24]
  wire  _add1_T_34 = tag_8[0] ^ tag_8[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_8 = _add1_T_34 ? fs_field8_8 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_16 = tag_8 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_8 = _add2_T_16 ? 8'h0 : phv_data_8; // @[executor_pisa.scala 268:24]
  wire  _add1_T_38 = tag_9[0] ^ tag_9[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_9 = _add1_T_38 ? fs_field8_9 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_18 = tag_9 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_9 = _add2_T_18 ? 8'h0 : phv_data_9; // @[executor_pisa.scala 268:24]
  wire  _add1_T_42 = tag_10[0] ^ tag_10[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_10 = _add1_T_42 ? fs_field8_10 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_20 = tag_10 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_10 = _add2_T_20 ? 8'h0 : phv_data_10; // @[executor_pisa.scala 268:24]
  wire  _add1_T_46 = tag_11[0] ^ tag_11[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_11 = _add1_T_46 ? fs_field8_11 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_22 = tag_11 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_11 = _add2_T_22 ? 8'h0 : phv_data_11; // @[executor_pisa.scala 268:24]
  wire  _add1_T_50 = tag_12[0] ^ tag_12[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_12 = _add1_T_50 ? fs_field8_12 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_24 = tag_12 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_12 = _add2_T_24 ? 8'h0 : phv_data_12; // @[executor_pisa.scala 268:24]
  wire  _add1_T_54 = tag_13[0] ^ tag_13[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_13 = _add1_T_54 ? fs_field8_13 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_26 = tag_13 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_13 = _add2_T_26 ? 8'h0 : phv_data_13; // @[executor_pisa.scala 268:24]
  wire  _add1_T_58 = tag_14[0] ^ tag_14[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_14 = _add1_T_58 ? fs_field8_14 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_28 = tag_14 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_14 = _add2_T_28 ? 8'h0 : phv_data_14; // @[executor_pisa.scala 268:24]
  wire  _add1_T_62 = tag_15[0] ^ tag_15[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_15 = _add1_T_62 ? fs_field8_15 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_30 = tag_15 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_15 = _add2_T_30 ? 8'h0 : phv_data_15; // @[executor_pisa.scala 268:24]
  wire  _add1_T_66 = tag_16[0] ^ tag_16[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_16 = _add1_T_66 ? fs_field8_16 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_32 = tag_16 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_16 = _add2_T_32 ? 8'h0 : phv_data_16; // @[executor_pisa.scala 268:24]
  wire  _add1_T_70 = tag_17[0] ^ tag_17[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_17 = _add1_T_70 ? fs_field8_17 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_34 = tag_17 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_17 = _add2_T_34 ? 8'h0 : phv_data_17; // @[executor_pisa.scala 268:24]
  wire  _add1_T_74 = tag_18[0] ^ tag_18[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_18 = _add1_T_74 ? fs_field8_18 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_36 = tag_18 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_18 = _add2_T_36 ? 8'h0 : phv_data_18; // @[executor_pisa.scala 268:24]
  wire  _add1_T_78 = tag_19[0] ^ tag_19[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_19 = _add1_T_78 ? fs_field8_19 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_38 = tag_19 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_19 = _add2_T_38 ? 8'h0 : phv_data_19; // @[executor_pisa.scala 268:24]
  wire  _add1_T_82 = tag_20[0] ^ tag_20[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_20 = _add1_T_82 ? fs_field8_20 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_40 = tag_20 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_20 = _add2_T_40 ? 8'h0 : phv_data_20; // @[executor_pisa.scala 268:24]
  wire  _add1_T_86 = tag_21[0] ^ tag_21[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_21 = _add1_T_86 ? fs_field8_21 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_42 = tag_21 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_21 = _add2_T_42 ? 8'h0 : phv_data_21; // @[executor_pisa.scala 268:24]
  wire  _add1_T_90 = tag_22[0] ^ tag_22[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_22 = _add1_T_90 ? fs_field8_22 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_44 = tag_22 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_22 = _add2_T_44 ? 8'h0 : phv_data_22; // @[executor_pisa.scala 268:24]
  wire  _add1_T_94 = tag_23[0] ^ tag_23[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_23 = _add1_T_94 ? fs_field8_23 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_46 = tag_23 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_23 = _add2_T_46 ? 8'h0 : phv_data_23; // @[executor_pisa.scala 268:24]
  wire  _add1_T_98 = tag_24[0] ^ tag_24[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_24 = _add1_T_98 ? fs_field8_24 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_48 = tag_24 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_24 = _add2_T_48 ? 8'h0 : phv_data_24; // @[executor_pisa.scala 268:24]
  wire  _add1_T_102 = tag_25[0] ^ tag_25[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_25 = _add1_T_102 ? fs_field8_25 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_50 = tag_25 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_25 = _add2_T_50 ? 8'h0 : phv_data_25; // @[executor_pisa.scala 268:24]
  wire  _add1_T_106 = tag_26[0] ^ tag_26[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_26 = _add1_T_106 ? fs_field8_26 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_52 = tag_26 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_26 = _add2_T_52 ? 8'h0 : phv_data_26; // @[executor_pisa.scala 268:24]
  wire  _add1_T_110 = tag_27[0] ^ tag_27[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_27 = _add1_T_110 ? fs_field8_27 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_54 = tag_27 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_27 = _add2_T_54 ? 8'h0 : phv_data_27; // @[executor_pisa.scala 268:24]
  wire  _add1_T_114 = tag_28[0] ^ tag_28[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_28 = _add1_T_114 ? fs_field8_28 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_56 = tag_28 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_28 = _add2_T_56 ? 8'h0 : phv_data_28; // @[executor_pisa.scala 268:24]
  wire  _add1_T_118 = tag_29[0] ^ tag_29[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_29 = _add1_T_118 ? fs_field8_29 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_58 = tag_29 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_29 = _add2_T_58 ? 8'h0 : phv_data_29; // @[executor_pisa.scala 268:24]
  wire  _add1_T_122 = tag_30[0] ^ tag_30[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_30 = _add1_T_122 ? fs_field8_30 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_60 = tag_30 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_30 = _add2_T_60 ? 8'h0 : phv_data_30; // @[executor_pisa.scala 268:24]
  wire  _add1_T_126 = tag_31[0] ^ tag_31[1]; // @[executor_pisa.scala 264:30]
  wire [7:0] add1_31 = _add1_T_126 ? fs_field8_31 : 8'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_62 = tag_31 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [7:0] add2_31 = _add2_T_62 ? 8'h0 : phv_data_31; // @[executor_pisa.scala 268:24]
  wire  _add1_T_130 = tag_32[0] ^ tag_32[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_32 = _add1_T_130 ? fs_field16_0 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_64 = tag_32 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_65 = {phv_data_32,phv_data_33}; // @[Cat.scala 30:58]
  wire [15:0] add2_32 = _add2_T_64 ? 16'h0 : _add2_T_65; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_65 = add1_32 + add2_32; // @[executor_pisa.scala 273:51]
  wire  _add1_T_134 = tag_33[0] ^ tag_33[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_33 = _add1_T_134 ? fs_field16_1 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_67 = tag_33 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_68 = {phv_data_34,phv_data_35}; // @[Cat.scala 30:58]
  wire [15:0] add2_33 = _add2_T_67 ? 16'h0 : _add2_T_68; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_67 = add1_33 + add2_33; // @[executor_pisa.scala 273:51]
  wire  _add1_T_138 = tag_34[0] ^ tag_34[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_34 = _add1_T_138 ? fs_field16_2 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_70 = tag_34 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_71 = {phv_data_36,phv_data_37}; // @[Cat.scala 30:58]
  wire [15:0] add2_34 = _add2_T_70 ? 16'h0 : _add2_T_71; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_69 = add1_34 + add2_34; // @[executor_pisa.scala 273:51]
  wire  _add1_T_142 = tag_35[0] ^ tag_35[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_35 = _add1_T_142 ? fs_field16_3 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_73 = tag_35 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_74 = {phv_data_38,phv_data_39}; // @[Cat.scala 30:58]
  wire [15:0] add2_35 = _add2_T_73 ? 16'h0 : _add2_T_74; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_71 = add1_35 + add2_35; // @[executor_pisa.scala 273:51]
  wire  _add1_T_146 = tag_36[0] ^ tag_36[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_36 = _add1_T_146 ? fs_field16_4 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_76 = tag_36 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_77 = {phv_data_40,phv_data_41}; // @[Cat.scala 30:58]
  wire [15:0] add2_36 = _add2_T_76 ? 16'h0 : _add2_T_77; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_73 = add1_36 + add2_36; // @[executor_pisa.scala 273:51]
  wire  _add1_T_150 = tag_37[0] ^ tag_37[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_37 = _add1_T_150 ? fs_field16_5 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_79 = tag_37 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_80 = {phv_data_42,phv_data_43}; // @[Cat.scala 30:58]
  wire [15:0] add2_37 = _add2_T_79 ? 16'h0 : _add2_T_80; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_75 = add1_37 + add2_37; // @[executor_pisa.scala 273:51]
  wire  _add1_T_154 = tag_38[0] ^ tag_38[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_38 = _add1_T_154 ? fs_field16_6 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_82 = tag_38 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_83 = {phv_data_44,phv_data_45}; // @[Cat.scala 30:58]
  wire [15:0] add2_38 = _add2_T_82 ? 16'h0 : _add2_T_83; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_77 = add1_38 + add2_38; // @[executor_pisa.scala 273:51]
  wire  _add1_T_158 = tag_39[0] ^ tag_39[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_39 = _add1_T_158 ? fs_field16_7 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_85 = tag_39 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_86 = {phv_data_46,phv_data_47}; // @[Cat.scala 30:58]
  wire [15:0] add2_39 = _add2_T_85 ? 16'h0 : _add2_T_86; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_79 = add1_39 + add2_39; // @[executor_pisa.scala 273:51]
  wire  _add1_T_162 = tag_40[0] ^ tag_40[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_40 = _add1_T_162 ? fs_field16_8 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_88 = tag_40 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_89 = {phv_data_48,phv_data_49}; // @[Cat.scala 30:58]
  wire [15:0] add2_40 = _add2_T_88 ? 16'h0 : _add2_T_89; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_81 = add1_40 + add2_40; // @[executor_pisa.scala 273:51]
  wire  _add1_T_166 = tag_41[0] ^ tag_41[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_41 = _add1_T_166 ? fs_field16_9 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_91 = tag_41 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_92 = {phv_data_50,phv_data_51}; // @[Cat.scala 30:58]
  wire [15:0] add2_41 = _add2_T_91 ? 16'h0 : _add2_T_92; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_83 = add1_41 + add2_41; // @[executor_pisa.scala 273:51]
  wire  _add1_T_170 = tag_42[0] ^ tag_42[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_42 = _add1_T_170 ? fs_field16_10 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_94 = tag_42 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_95 = {phv_data_52,phv_data_53}; // @[Cat.scala 30:58]
  wire [15:0] add2_42 = _add2_T_94 ? 16'h0 : _add2_T_95; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_85 = add1_42 + add2_42; // @[executor_pisa.scala 273:51]
  wire  _add1_T_174 = tag_43[0] ^ tag_43[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_43 = _add1_T_174 ? fs_field16_11 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_97 = tag_43 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_98 = {phv_data_54,phv_data_55}; // @[Cat.scala 30:58]
  wire [15:0] add2_43 = _add2_T_97 ? 16'h0 : _add2_T_98; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_87 = add1_43 + add2_43; // @[executor_pisa.scala 273:51]
  wire  _add1_T_178 = tag_44[0] ^ tag_44[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_44 = _add1_T_178 ? fs_field16_12 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_100 = tag_44 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_101 = {phv_data_56,phv_data_57}; // @[Cat.scala 30:58]
  wire [15:0] add2_44 = _add2_T_100 ? 16'h0 : _add2_T_101; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_89 = add1_44 + add2_44; // @[executor_pisa.scala 273:51]
  wire  _add1_T_182 = tag_45[0] ^ tag_45[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_45 = _add1_T_182 ? fs_field16_13 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_103 = tag_45 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_104 = {phv_data_58,phv_data_59}; // @[Cat.scala 30:58]
  wire [15:0] add2_45 = _add2_T_103 ? 16'h0 : _add2_T_104; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_91 = add1_45 + add2_45; // @[executor_pisa.scala 273:51]
  wire  _add1_T_186 = tag_46[0] ^ tag_46[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_46 = _add1_T_186 ? fs_field16_14 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_106 = tag_46 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_107 = {phv_data_60,phv_data_61}; // @[Cat.scala 30:58]
  wire [15:0] add2_46 = _add2_T_106 ? 16'h0 : _add2_T_107; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_93 = add1_46 + add2_46; // @[executor_pisa.scala 273:51]
  wire  _add1_T_190 = tag_47[0] ^ tag_47[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_47 = _add1_T_190 ? fs_field16_15 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_109 = tag_47 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_110 = {phv_data_62,phv_data_63}; // @[Cat.scala 30:58]
  wire [15:0] add2_47 = _add2_T_109 ? 16'h0 : _add2_T_110; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_95 = add1_47 + add2_47; // @[executor_pisa.scala 273:51]
  wire  _add1_T_194 = tag_48[0] ^ tag_48[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_48 = _add1_T_194 ? fs_field16_16 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_112 = tag_48 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_113 = {phv_data_64,phv_data_65}; // @[Cat.scala 30:58]
  wire [15:0] add2_48 = _add2_T_112 ? 16'h0 : _add2_T_113; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_97 = add1_48 + add2_48; // @[executor_pisa.scala 273:51]
  wire  _add1_T_198 = tag_49[0] ^ tag_49[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_49 = _add1_T_198 ? fs_field16_17 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_115 = tag_49 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_116 = {phv_data_66,phv_data_67}; // @[Cat.scala 30:58]
  wire [15:0] add2_49 = _add2_T_115 ? 16'h0 : _add2_T_116; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_99 = add1_49 + add2_49; // @[executor_pisa.scala 273:51]
  wire  _add1_T_202 = tag_50[0] ^ tag_50[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_50 = _add1_T_202 ? fs_field16_18 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_118 = tag_50 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_119 = {phv_data_68,phv_data_69}; // @[Cat.scala 30:58]
  wire [15:0] add2_50 = _add2_T_118 ? 16'h0 : _add2_T_119; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_101 = add1_50 + add2_50; // @[executor_pisa.scala 273:51]
  wire  _add1_T_206 = tag_51[0] ^ tag_51[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_51 = _add1_T_206 ? fs_field16_19 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_121 = tag_51 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_122 = {phv_data_70,phv_data_71}; // @[Cat.scala 30:58]
  wire [15:0] add2_51 = _add2_T_121 ? 16'h0 : _add2_T_122; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_103 = add1_51 + add2_51; // @[executor_pisa.scala 273:51]
  wire  _add1_T_210 = tag_52[0] ^ tag_52[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_52 = _add1_T_210 ? fs_field16_20 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_124 = tag_52 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_125 = {phv_data_72,phv_data_73}; // @[Cat.scala 30:58]
  wire [15:0] add2_52 = _add2_T_124 ? 16'h0 : _add2_T_125; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_105 = add1_52 + add2_52; // @[executor_pisa.scala 273:51]
  wire  _add1_T_214 = tag_53[0] ^ tag_53[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_53 = _add1_T_214 ? fs_field16_21 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_127 = tag_53 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_128 = {phv_data_74,phv_data_75}; // @[Cat.scala 30:58]
  wire [15:0] add2_53 = _add2_T_127 ? 16'h0 : _add2_T_128; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_107 = add1_53 + add2_53; // @[executor_pisa.scala 273:51]
  wire  _add1_T_218 = tag_54[0] ^ tag_54[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_54 = _add1_T_218 ? fs_field16_22 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_130 = tag_54 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_131 = {phv_data_76,phv_data_77}; // @[Cat.scala 30:58]
  wire [15:0] add2_54 = _add2_T_130 ? 16'h0 : _add2_T_131; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_109 = add1_54 + add2_54; // @[executor_pisa.scala 273:51]
  wire  _add1_T_222 = tag_55[0] ^ tag_55[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_55 = _add1_T_222 ? fs_field16_23 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_133 = tag_55 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_134 = {phv_data_78,phv_data_79}; // @[Cat.scala 30:58]
  wire [15:0] add2_55 = _add2_T_133 ? 16'h0 : _add2_T_134; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_111 = add1_55 + add2_55; // @[executor_pisa.scala 273:51]
  wire  _add1_T_226 = tag_56[0] ^ tag_56[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_56 = _add1_T_226 ? fs_field16_24 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_136 = tag_56 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_137 = {phv_data_80,phv_data_81}; // @[Cat.scala 30:58]
  wire [15:0] add2_56 = _add2_T_136 ? 16'h0 : _add2_T_137; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_113 = add1_56 + add2_56; // @[executor_pisa.scala 273:51]
  wire  _add1_T_230 = tag_57[0] ^ tag_57[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_57 = _add1_T_230 ? fs_field16_25 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_139 = tag_57 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_140 = {phv_data_82,phv_data_83}; // @[Cat.scala 30:58]
  wire [15:0] add2_57 = _add2_T_139 ? 16'h0 : _add2_T_140; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_115 = add1_57 + add2_57; // @[executor_pisa.scala 273:51]
  wire  _add1_T_234 = tag_58[0] ^ tag_58[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_58 = _add1_T_234 ? fs_field16_26 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_142 = tag_58 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_143 = {phv_data_84,phv_data_85}; // @[Cat.scala 30:58]
  wire [15:0] add2_58 = _add2_T_142 ? 16'h0 : _add2_T_143; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_117 = add1_58 + add2_58; // @[executor_pisa.scala 273:51]
  wire  _add1_T_238 = tag_59[0] ^ tag_59[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_59 = _add1_T_238 ? fs_field16_27 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_145 = tag_59 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_146 = {phv_data_86,phv_data_87}; // @[Cat.scala 30:58]
  wire [15:0] add2_59 = _add2_T_145 ? 16'h0 : _add2_T_146; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_119 = add1_59 + add2_59; // @[executor_pisa.scala 273:51]
  wire  _add1_T_242 = tag_60[0] ^ tag_60[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_60 = _add1_T_242 ? fs_field16_28 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_148 = tag_60 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_149 = {phv_data_88,phv_data_89}; // @[Cat.scala 30:58]
  wire [15:0] add2_60 = _add2_T_148 ? 16'h0 : _add2_T_149; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_121 = add1_60 + add2_60; // @[executor_pisa.scala 273:51]
  wire  _add1_T_246 = tag_61[0] ^ tag_61[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_61 = _add1_T_246 ? fs_field16_29 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_151 = tag_61 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_152 = {phv_data_90,phv_data_91}; // @[Cat.scala 30:58]
  wire [15:0] add2_61 = _add2_T_151 ? 16'h0 : _add2_T_152; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_123 = add1_61 + add2_61; // @[executor_pisa.scala 273:51]
  wire  _add1_T_250 = tag_62[0] ^ tag_62[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_62 = _add1_T_250 ? fs_field16_30 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_154 = tag_62 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_155 = {phv_data_92,phv_data_93}; // @[Cat.scala 30:58]
  wire [15:0] add2_62 = _add2_T_154 ? 16'h0 : _add2_T_155; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_125 = add1_62 + add2_62; // @[executor_pisa.scala 273:51]
  wire  _add1_T_254 = tag_63[0] ^ tag_63[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_63 = _add1_T_254 ? fs_field16_31 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_157 = tag_63 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_158 = {phv_data_94,phv_data_95}; // @[Cat.scala 30:58]
  wire [15:0] add2_63 = _add2_T_157 ? 16'h0 : _add2_T_158; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_127 = add1_63 + add2_63; // @[executor_pisa.scala 273:51]
  wire  _add1_T_258 = tag_64[0] ^ tag_64[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_64 = _add1_T_258 ? fs_field16_32 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_160 = tag_64 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_161 = {phv_data_96,phv_data_97}; // @[Cat.scala 30:58]
  wire [15:0] add2_64 = _add2_T_160 ? 16'h0 : _add2_T_161; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_129 = add1_64 + add2_64; // @[executor_pisa.scala 273:51]
  wire  _add1_T_262 = tag_65[0] ^ tag_65[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_65 = _add1_T_262 ? fs_field16_33 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_163 = tag_65 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_164 = {phv_data_98,phv_data_99}; // @[Cat.scala 30:58]
  wire [15:0] add2_65 = _add2_T_163 ? 16'h0 : _add2_T_164; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_131 = add1_65 + add2_65; // @[executor_pisa.scala 273:51]
  wire  _add1_T_266 = tag_66[0] ^ tag_66[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_66 = _add1_T_266 ? fs_field16_34 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_166 = tag_66 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_167 = {phv_data_100,phv_data_101}; // @[Cat.scala 30:58]
  wire [15:0] add2_66 = _add2_T_166 ? 16'h0 : _add2_T_167; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_133 = add1_66 + add2_66; // @[executor_pisa.scala 273:51]
  wire  _add1_T_270 = tag_67[0] ^ tag_67[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_67 = _add1_T_270 ? fs_field16_35 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_169 = tag_67 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_170 = {phv_data_102,phv_data_103}; // @[Cat.scala 30:58]
  wire [15:0] add2_67 = _add2_T_169 ? 16'h0 : _add2_T_170; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_135 = add1_67 + add2_67; // @[executor_pisa.scala 273:51]
  wire  _add1_T_274 = tag_68[0] ^ tag_68[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_68 = _add1_T_274 ? fs_field16_36 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_172 = tag_68 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_173 = {phv_data_104,phv_data_105}; // @[Cat.scala 30:58]
  wire [15:0] add2_68 = _add2_T_172 ? 16'h0 : _add2_T_173; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_137 = add1_68 + add2_68; // @[executor_pisa.scala 273:51]
  wire  _add1_T_278 = tag_69[0] ^ tag_69[1]; // @[executor_pisa.scala 264:30]
  wire [15:0] add1_69 = _add1_T_278 ? fs_field16_37 : 16'h0; // @[executor_pisa.scala 263:24]
  wire  _add2_T_175 = tag_69 == 2'h2; // @[executor_pisa.scala 269:27]
  wire [15:0] _add2_T_176 = {phv_data_106,phv_data_107}; // @[Cat.scala 30:58]
  wire [15:0] add2_69 = _add2_T_175 ? 16'h0 : _add2_T_176; // @[executor_pisa.scala 268:24]
  wire [15:0] _T_139 = add1_69 + add2_69; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_0 = add1 + add2; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_1 = add1_1 + add2_1; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_2 = add1_2 + add2_2; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_3 = add1_3 + add2_3; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_4 = add1_4 + add2_4; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_5 = add1_5 + add2_5; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_6 = add1_6 + add2_6; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_7 = add1_7 + add2_7; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_8 = add1_8 + add2_8; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_9 = add1_9 + add2_9; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_10 = add1_10 + add2_10; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_11 = add1_11 + add2_11; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_12 = add1_12 + add2_12; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_13 = add1_13 + add2_13; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_14 = add1_14 + add2_14; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_15 = add1_15 + add2_15; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_16 = add1_16 + add2_16; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_17 = add1_17 + add2_17; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_18 = add1_18 + add2_18; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_19 = add1_19 + add2_19; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_20 = add1_20 + add2_20; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_21 = add1_21 + add2_21; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_22 = add1_22 + add2_22; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_23 = add1_23 + add2_23; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_24 = add1_24 + add2_24; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_25 = add1_25 + add2_25; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_26 = add1_26 + add2_26; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_27 = add1_27 + add2_27; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_28 = add1_28 + add2_28; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_29 = add1_29 + add2_29; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_30 = add1_30 + add2_30; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_31 = add1_31 + add2_31; // @[executor_pisa.scala 273:51]
  assign io_pipe_phv_out_data_32 = _T_65[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_33 = _T_65[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_34 = _T_67[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_35 = _T_67[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_36 = _T_69[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_37 = _T_69[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_38 = _T_71[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_39 = _T_71[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_40 = _T_73[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_41 = _T_73[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_42 = _T_75[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_43 = _T_75[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_44 = _T_77[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_45 = _T_77[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_46 = _T_79[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_47 = _T_79[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_48 = _T_81[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_49 = _T_81[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_50 = _T_83[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_51 = _T_83[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_52 = _T_85[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_53 = _T_85[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_54 = _T_87[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_55 = _T_87[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_56 = _T_89[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_57 = _T_89[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_58 = _T_91[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_59 = _T_91[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_60 = _T_93[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_61 = _T_93[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_62 = _T_95[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_63 = _T_95[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_64 = _T_97[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_65 = _T_97[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_66 = _T_99[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_67 = _T_99[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_68 = _T_101[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_69 = _T_101[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_70 = _T_103[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_71 = _T_103[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_72 = _T_105[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_73 = _T_105[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_74 = _T_107[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_75 = _T_107[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_76 = _T_109[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_77 = _T_109[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_78 = _T_111[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_79 = _T_111[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_80 = _T_113[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_81 = _T_113[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_82 = _T_115[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_83 = _T_115[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_84 = _T_117[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_85 = _T_117[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_86 = _T_119[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_87 = _T_119[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_88 = _T_121[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_89 = _T_121[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_90 = _T_123[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_91 = _T_123[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_92 = _T_125[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_93 = _T_125[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_94 = _T_127[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_95 = _T_127[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_96 = _T_129[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_97 = _T_129[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_98 = _T_131[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_99 = _T_131[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_100 = _T_133[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_101 = _T_133[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_102 = _T_135[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_103 = _T_135[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_104 = _T_137[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_105 = _T_137[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_106 = _T_139[15:8]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_107 = _T_139[7:0]; // @[executor_pisa.scala 232:46]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[executor_pisa.scala 246:25]
  assign io_pipe_phv_out_next_processor_id = nid[14] ? nid[13:10] : phv_next_processor_id; // @[executor_pisa.scala 276:24 executor_pisa.scala 277:47 executor_pisa.scala 246:25]
  assign io_pipe_phv_out_next_config_id = nid[14] ? nid[0] : phv_next_config_id; // @[executor_pisa.scala 276:24 executor_pisa.scala 278:47 executor_pisa.scala 246:25]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor_pisa.scala 245:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor_pisa.scala 245:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor_pisa.scala 245:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor_pisa.scala 245:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor_pisa.scala 245:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor_pisa.scala 245:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor_pisa.scala 245:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor_pisa.scala 245:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor_pisa.scala 245:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor_pisa.scala 245:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor_pisa.scala 245:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor_pisa.scala 245:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor_pisa.scala 245:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor_pisa.scala 245:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor_pisa.scala 245:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor_pisa.scala 245:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor_pisa.scala 245:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor_pisa.scala 245:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor_pisa.scala 245:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor_pisa.scala 245:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor_pisa.scala 245:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor_pisa.scala 245:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor_pisa.scala 245:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor_pisa.scala 245:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor_pisa.scala 245:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor_pisa.scala 245:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor_pisa.scala 245:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor_pisa.scala 245:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor_pisa.scala 245:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor_pisa.scala 245:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor_pisa.scala 245:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor_pisa.scala 245:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor_pisa.scala 245:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor_pisa.scala 245:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor_pisa.scala 245:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor_pisa.scala 245:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor_pisa.scala 245:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor_pisa.scala 245:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor_pisa.scala 245:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor_pisa.scala 245:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor_pisa.scala 245:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor_pisa.scala 245:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor_pisa.scala 245:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor_pisa.scala 245:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor_pisa.scala 245:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor_pisa.scala 245:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor_pisa.scala 245:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor_pisa.scala 245:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor_pisa.scala 245:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor_pisa.scala 245:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor_pisa.scala 245:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor_pisa.scala 245:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor_pisa.scala 245:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor_pisa.scala 245:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor_pisa.scala 245:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor_pisa.scala 245:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor_pisa.scala 245:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor_pisa.scala 245:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor_pisa.scala 245:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor_pisa.scala 245:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor_pisa.scala 245:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor_pisa.scala 245:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor_pisa.scala 245:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor_pisa.scala 245:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor_pisa.scala 245:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor_pisa.scala 245:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor_pisa.scala 245:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor_pisa.scala 245:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor_pisa.scala 245:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor_pisa.scala 245:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor_pisa.scala 245:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor_pisa.scala 245:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor_pisa.scala 245:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor_pisa.scala 245:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor_pisa.scala 245:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor_pisa.scala 245:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor_pisa.scala 245:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor_pisa.scala 245:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor_pisa.scala 245:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor_pisa.scala 245:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor_pisa.scala 245:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor_pisa.scala 245:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor_pisa.scala 245:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor_pisa.scala 245:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor_pisa.scala 245:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor_pisa.scala 245:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor_pisa.scala 245:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor_pisa.scala 245:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor_pisa.scala 245:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor_pisa.scala 245:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor_pisa.scala 245:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor_pisa.scala 245:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor_pisa.scala 245:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor_pisa.scala 245:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor_pisa.scala 245:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor_pisa.scala 245:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor_pisa.scala 245:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor_pisa.scala 245:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor_pisa.scala 245:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor_pisa.scala 245:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor_pisa.scala 245:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor_pisa.scala 245:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor_pisa.scala 245:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor_pisa.scala 245:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor_pisa.scala 245:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor_pisa.scala 245:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor_pisa.scala 245:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor_pisa.scala 245:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor_pisa.scala 245:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor_pisa.scala 245:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor_pisa.scala 245:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor_pisa.scala 245:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor_pisa.scala 245:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor_pisa.scala 245:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor_pisa.scala 245:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor_pisa.scala 245:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor_pisa.scala 245:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor_pisa.scala 245:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor_pisa.scala 245:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor_pisa.scala 245:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor_pisa.scala 245:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor_pisa.scala 245:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor_pisa.scala 245:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor_pisa.scala 245:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor_pisa.scala 245:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor_pisa.scala 245:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor_pisa.scala 245:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor_pisa.scala 245:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor_pisa.scala 245:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor_pisa.scala 245:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor_pisa.scala 245:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor_pisa.scala 245:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor_pisa.scala 245:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor_pisa.scala 245:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor_pisa.scala 245:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor_pisa.scala 245:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor_pisa.scala 245:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor_pisa.scala 245:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor_pisa.scala 245:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor_pisa.scala 245:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor_pisa.scala 245:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor_pisa.scala 245:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor_pisa.scala 245:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor_pisa.scala 245:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor_pisa.scala 245:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor_pisa.scala 245:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor_pisa.scala 245:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor_pisa.scala 245:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor_pisa.scala 245:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor_pisa.scala 245:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor_pisa.scala 245:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor_pisa.scala 245:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor_pisa.scala 245:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor_pisa.scala 245:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor_pisa.scala 245:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor_pisa.scala 245:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor_pisa.scala 245:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor_pisa.scala 245:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor_pisa.scala 245:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor_pisa.scala 245:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor_pisa.scala 245:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor_pisa.scala 245:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor_pisa.scala 245:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor_pisa.scala 245:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor_pisa.scala 245:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor_pisa.scala 245:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor_pisa.scala 245:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor_pisa.scala 245:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor_pisa.scala 245:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor_pisa.scala 245:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor_pisa.scala 245:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor_pisa.scala 245:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor_pisa.scala 245:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor_pisa.scala 245:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor_pisa.scala 245:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor_pisa.scala 245:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor_pisa.scala 245:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor_pisa.scala 245:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor_pisa.scala 245:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor_pisa.scala 245:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor_pisa.scala 245:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor_pisa.scala 245:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor_pisa.scala 245:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor_pisa.scala 245:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor_pisa.scala 245:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor_pisa.scala 245:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor_pisa.scala 245:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor_pisa.scala 245:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor_pisa.scala 245:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor_pisa.scala 245:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor_pisa.scala 245:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor_pisa.scala 245:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor_pisa.scala 245:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor_pisa.scala 245:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor_pisa.scala 245:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor_pisa.scala 245:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor_pisa.scala 245:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor_pisa.scala 245:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor_pisa.scala 245:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor_pisa.scala 245:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor_pisa.scala 245:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor_pisa.scala 245:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor_pisa.scala 245:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor_pisa.scala 245:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor_pisa.scala 245:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor_pisa.scala 245:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor_pisa.scala 245:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor_pisa.scala 245:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor_pisa.scala 245:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor_pisa.scala 245:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor_pisa.scala 245:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor_pisa.scala 245:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor_pisa.scala 245:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor_pisa.scala 245:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor_pisa.scala 245:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor_pisa.scala 245:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor_pisa.scala 245:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor_pisa.scala 245:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor_pisa.scala 245:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor_pisa.scala 245:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor_pisa.scala 245:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor_pisa.scala 245:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor_pisa.scala 245:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor_pisa.scala 245:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor_pisa.scala 245:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor_pisa.scala 245:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor_pisa.scala 245:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor_pisa.scala 245:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor_pisa.scala 245:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor_pisa.scala 245:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor_pisa.scala 245:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor_pisa.scala 245:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor_pisa.scala 245:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor_pisa.scala 245:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor_pisa.scala 245:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor_pisa.scala 245:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor_pisa.scala 245:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor_pisa.scala 245:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor_pisa.scala 245:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor_pisa.scala 245:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor_pisa.scala 245:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor_pisa.scala 245:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor_pisa.scala 245:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor_pisa.scala 245:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor_pisa.scala 245:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor_pisa.scala 245:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor_pisa.scala 245:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor_pisa.scala 245:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor_pisa.scala 245:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor_pisa.scala 245:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor_pisa.scala 245:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor_pisa.scala 245:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor_pisa.scala 245:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor_pisa.scala 245:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor_pisa.scala 245:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor_pisa.scala 245:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor_pisa.scala 245:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 245:13]
    fs_field8_0 <= io_field_set_field8_0; // @[executor_pisa.scala 249:12]
    fs_field8_1 <= io_field_set_field8_1; // @[executor_pisa.scala 249:12]
    fs_field8_2 <= io_field_set_field8_2; // @[executor_pisa.scala 249:12]
    fs_field8_3 <= io_field_set_field8_3; // @[executor_pisa.scala 249:12]
    fs_field8_4 <= io_field_set_field8_4; // @[executor_pisa.scala 249:12]
    fs_field8_5 <= io_field_set_field8_5; // @[executor_pisa.scala 249:12]
    fs_field8_6 <= io_field_set_field8_6; // @[executor_pisa.scala 249:12]
    fs_field8_7 <= io_field_set_field8_7; // @[executor_pisa.scala 249:12]
    fs_field8_8 <= io_field_set_field8_8; // @[executor_pisa.scala 249:12]
    fs_field8_9 <= io_field_set_field8_9; // @[executor_pisa.scala 249:12]
    fs_field8_10 <= io_field_set_field8_10; // @[executor_pisa.scala 249:12]
    fs_field8_11 <= io_field_set_field8_11; // @[executor_pisa.scala 249:12]
    fs_field8_12 <= io_field_set_field8_12; // @[executor_pisa.scala 249:12]
    fs_field8_13 <= io_field_set_field8_13; // @[executor_pisa.scala 249:12]
    fs_field8_14 <= io_field_set_field8_14; // @[executor_pisa.scala 249:12]
    fs_field8_15 <= io_field_set_field8_15; // @[executor_pisa.scala 249:12]
    fs_field8_16 <= io_field_set_field8_16; // @[executor_pisa.scala 249:12]
    fs_field8_17 <= io_field_set_field8_17; // @[executor_pisa.scala 249:12]
    fs_field8_18 <= io_field_set_field8_18; // @[executor_pisa.scala 249:12]
    fs_field8_19 <= io_field_set_field8_19; // @[executor_pisa.scala 249:12]
    fs_field8_20 <= io_field_set_field8_20; // @[executor_pisa.scala 249:12]
    fs_field8_21 <= io_field_set_field8_21; // @[executor_pisa.scala 249:12]
    fs_field8_22 <= io_field_set_field8_22; // @[executor_pisa.scala 249:12]
    fs_field8_23 <= io_field_set_field8_23; // @[executor_pisa.scala 249:12]
    fs_field8_24 <= io_field_set_field8_24; // @[executor_pisa.scala 249:12]
    fs_field8_25 <= io_field_set_field8_25; // @[executor_pisa.scala 249:12]
    fs_field8_26 <= io_field_set_field8_26; // @[executor_pisa.scala 249:12]
    fs_field8_27 <= io_field_set_field8_27; // @[executor_pisa.scala 249:12]
    fs_field8_28 <= io_field_set_field8_28; // @[executor_pisa.scala 249:12]
    fs_field8_29 <= io_field_set_field8_29; // @[executor_pisa.scala 249:12]
    fs_field8_30 <= io_field_set_field8_30; // @[executor_pisa.scala 249:12]
    fs_field8_31 <= io_field_set_field8_31; // @[executor_pisa.scala 249:12]
    fs_field16_0 <= io_field_set_field16_0; // @[executor_pisa.scala 249:12]
    fs_field16_1 <= io_field_set_field16_1; // @[executor_pisa.scala 249:12]
    fs_field16_2 <= io_field_set_field16_2; // @[executor_pisa.scala 249:12]
    fs_field16_3 <= io_field_set_field16_3; // @[executor_pisa.scala 249:12]
    fs_field16_4 <= io_field_set_field16_4; // @[executor_pisa.scala 249:12]
    fs_field16_5 <= io_field_set_field16_5; // @[executor_pisa.scala 249:12]
    fs_field16_6 <= io_field_set_field16_6; // @[executor_pisa.scala 249:12]
    fs_field16_7 <= io_field_set_field16_7; // @[executor_pisa.scala 249:12]
    fs_field16_8 <= io_field_set_field16_8; // @[executor_pisa.scala 249:12]
    fs_field16_9 <= io_field_set_field16_9; // @[executor_pisa.scala 249:12]
    fs_field16_10 <= io_field_set_field16_10; // @[executor_pisa.scala 249:12]
    fs_field16_11 <= io_field_set_field16_11; // @[executor_pisa.scala 249:12]
    fs_field16_12 <= io_field_set_field16_12; // @[executor_pisa.scala 249:12]
    fs_field16_13 <= io_field_set_field16_13; // @[executor_pisa.scala 249:12]
    fs_field16_14 <= io_field_set_field16_14; // @[executor_pisa.scala 249:12]
    fs_field16_15 <= io_field_set_field16_15; // @[executor_pisa.scala 249:12]
    fs_field16_16 <= io_field_set_field16_16; // @[executor_pisa.scala 249:12]
    fs_field16_17 <= io_field_set_field16_17; // @[executor_pisa.scala 249:12]
    fs_field16_18 <= io_field_set_field16_18; // @[executor_pisa.scala 249:12]
    fs_field16_19 <= io_field_set_field16_19; // @[executor_pisa.scala 249:12]
    fs_field16_20 <= io_field_set_field16_20; // @[executor_pisa.scala 249:12]
    fs_field16_21 <= io_field_set_field16_21; // @[executor_pisa.scala 249:12]
    fs_field16_22 <= io_field_set_field16_22; // @[executor_pisa.scala 249:12]
    fs_field16_23 <= io_field_set_field16_23; // @[executor_pisa.scala 249:12]
    fs_field16_24 <= io_field_set_field16_24; // @[executor_pisa.scala 249:12]
    fs_field16_25 <= io_field_set_field16_25; // @[executor_pisa.scala 249:12]
    fs_field16_26 <= io_field_set_field16_26; // @[executor_pisa.scala 249:12]
    fs_field16_27 <= io_field_set_field16_27; // @[executor_pisa.scala 249:12]
    fs_field16_28 <= io_field_set_field16_28; // @[executor_pisa.scala 249:12]
    fs_field16_29 <= io_field_set_field16_29; // @[executor_pisa.scala 249:12]
    fs_field16_30 <= io_field_set_field16_30; // @[executor_pisa.scala 249:12]
    fs_field16_31 <= io_field_set_field16_31; // @[executor_pisa.scala 249:12]
    fs_field16_32 <= io_field_set_field16_32; // @[executor_pisa.scala 249:12]
    fs_field16_33 <= io_field_set_field16_33; // @[executor_pisa.scala 249:12]
    fs_field16_34 <= io_field_set_field16_34; // @[executor_pisa.scala 249:12]
    fs_field16_35 <= io_field_set_field16_35; // @[executor_pisa.scala 249:12]
    fs_field16_36 <= io_field_set_field16_36; // @[executor_pisa.scala 249:12]
    fs_field16_37 <= io_field_set_field16_37; // @[executor_pisa.scala 249:12]
    tag_0 <= io_tag_in_0; // @[executor_pisa.scala 252:13]
    tag_1 <= io_tag_in_1; // @[executor_pisa.scala 252:13]
    tag_2 <= io_tag_in_2; // @[executor_pisa.scala 252:13]
    tag_3 <= io_tag_in_3; // @[executor_pisa.scala 252:13]
    tag_4 <= io_tag_in_4; // @[executor_pisa.scala 252:13]
    tag_5 <= io_tag_in_5; // @[executor_pisa.scala 252:13]
    tag_6 <= io_tag_in_6; // @[executor_pisa.scala 252:13]
    tag_7 <= io_tag_in_7; // @[executor_pisa.scala 252:13]
    tag_8 <= io_tag_in_8; // @[executor_pisa.scala 252:13]
    tag_9 <= io_tag_in_9; // @[executor_pisa.scala 252:13]
    tag_10 <= io_tag_in_10; // @[executor_pisa.scala 252:13]
    tag_11 <= io_tag_in_11; // @[executor_pisa.scala 252:13]
    tag_12 <= io_tag_in_12; // @[executor_pisa.scala 252:13]
    tag_13 <= io_tag_in_13; // @[executor_pisa.scala 252:13]
    tag_14 <= io_tag_in_14; // @[executor_pisa.scala 252:13]
    tag_15 <= io_tag_in_15; // @[executor_pisa.scala 252:13]
    tag_16 <= io_tag_in_16; // @[executor_pisa.scala 252:13]
    tag_17 <= io_tag_in_17; // @[executor_pisa.scala 252:13]
    tag_18 <= io_tag_in_18; // @[executor_pisa.scala 252:13]
    tag_19 <= io_tag_in_19; // @[executor_pisa.scala 252:13]
    tag_20 <= io_tag_in_20; // @[executor_pisa.scala 252:13]
    tag_21 <= io_tag_in_21; // @[executor_pisa.scala 252:13]
    tag_22 <= io_tag_in_22; // @[executor_pisa.scala 252:13]
    tag_23 <= io_tag_in_23; // @[executor_pisa.scala 252:13]
    tag_24 <= io_tag_in_24; // @[executor_pisa.scala 252:13]
    tag_25 <= io_tag_in_25; // @[executor_pisa.scala 252:13]
    tag_26 <= io_tag_in_26; // @[executor_pisa.scala 252:13]
    tag_27 <= io_tag_in_27; // @[executor_pisa.scala 252:13]
    tag_28 <= io_tag_in_28; // @[executor_pisa.scala 252:13]
    tag_29 <= io_tag_in_29; // @[executor_pisa.scala 252:13]
    tag_30 <= io_tag_in_30; // @[executor_pisa.scala 252:13]
    tag_31 <= io_tag_in_31; // @[executor_pisa.scala 252:13]
    tag_32 <= io_tag_in_32; // @[executor_pisa.scala 252:13]
    tag_33 <= io_tag_in_33; // @[executor_pisa.scala 252:13]
    tag_34 <= io_tag_in_34; // @[executor_pisa.scala 252:13]
    tag_35 <= io_tag_in_35; // @[executor_pisa.scala 252:13]
    tag_36 <= io_tag_in_36; // @[executor_pisa.scala 252:13]
    tag_37 <= io_tag_in_37; // @[executor_pisa.scala 252:13]
    tag_38 <= io_tag_in_38; // @[executor_pisa.scala 252:13]
    tag_39 <= io_tag_in_39; // @[executor_pisa.scala 252:13]
    tag_40 <= io_tag_in_40; // @[executor_pisa.scala 252:13]
    tag_41 <= io_tag_in_41; // @[executor_pisa.scala 252:13]
    tag_42 <= io_tag_in_42; // @[executor_pisa.scala 252:13]
    tag_43 <= io_tag_in_43; // @[executor_pisa.scala 252:13]
    tag_44 <= io_tag_in_44; // @[executor_pisa.scala 252:13]
    tag_45 <= io_tag_in_45; // @[executor_pisa.scala 252:13]
    tag_46 <= io_tag_in_46; // @[executor_pisa.scala 252:13]
    tag_47 <= io_tag_in_47; // @[executor_pisa.scala 252:13]
    tag_48 <= io_tag_in_48; // @[executor_pisa.scala 252:13]
    tag_49 <= io_tag_in_49; // @[executor_pisa.scala 252:13]
    tag_50 <= io_tag_in_50; // @[executor_pisa.scala 252:13]
    tag_51 <= io_tag_in_51; // @[executor_pisa.scala 252:13]
    tag_52 <= io_tag_in_52; // @[executor_pisa.scala 252:13]
    tag_53 <= io_tag_in_53; // @[executor_pisa.scala 252:13]
    tag_54 <= io_tag_in_54; // @[executor_pisa.scala 252:13]
    tag_55 <= io_tag_in_55; // @[executor_pisa.scala 252:13]
    tag_56 <= io_tag_in_56; // @[executor_pisa.scala 252:13]
    tag_57 <= io_tag_in_57; // @[executor_pisa.scala 252:13]
    tag_58 <= io_tag_in_58; // @[executor_pisa.scala 252:13]
    tag_59 <= io_tag_in_59; // @[executor_pisa.scala 252:13]
    tag_60 <= io_tag_in_60; // @[executor_pisa.scala 252:13]
    tag_61 <= io_tag_in_61; // @[executor_pisa.scala 252:13]
    tag_62 <= io_tag_in_62; // @[executor_pisa.scala 252:13]
    tag_63 <= io_tag_in_63; // @[executor_pisa.scala 252:13]
    tag_64 <= io_tag_in_64; // @[executor_pisa.scala 252:13]
    tag_65 <= io_tag_in_65; // @[executor_pisa.scala 252:13]
    tag_66 <= io_tag_in_66; // @[executor_pisa.scala 252:13]
    tag_67 <= io_tag_in_67; // @[executor_pisa.scala 252:13]
    tag_68 <= io_tag_in_68; // @[executor_pisa.scala 252:13]
    tag_69 <= io_tag_in_69; // @[executor_pisa.scala 252:13]
    nid <= io_nid_in; // @[executor_pisa.scala 255:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  phv_next_config_id = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  fs_field8_0 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  fs_field8_1 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  fs_field8_2 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  fs_field8_3 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  fs_field8_4 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  fs_field8_5 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  fs_field8_6 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  fs_field8_7 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  fs_field8_8 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  fs_field8_9 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  fs_field8_10 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  fs_field8_11 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  fs_field8_12 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  fs_field8_13 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  fs_field8_14 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  fs_field8_15 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  fs_field8_16 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  fs_field8_17 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  fs_field8_18 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  fs_field8_19 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  fs_field8_20 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  fs_field8_21 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  fs_field8_22 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  fs_field8_23 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  fs_field8_24 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  fs_field8_25 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  fs_field8_26 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  fs_field8_27 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  fs_field8_28 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  fs_field8_29 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  fs_field8_30 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  fs_field8_31 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  fs_field16_0 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  fs_field16_1 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  fs_field16_2 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  fs_field16_3 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  fs_field16_4 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  fs_field16_5 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  fs_field16_6 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  fs_field16_7 = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  fs_field16_8 = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  fs_field16_9 = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  fs_field16_10 = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  fs_field16_11 = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  fs_field16_12 = _RAND_302[15:0];
  _RAND_303 = {1{`RANDOM}};
  fs_field16_13 = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  fs_field16_14 = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  fs_field16_15 = _RAND_305[15:0];
  _RAND_306 = {1{`RANDOM}};
  fs_field16_16 = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  fs_field16_17 = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  fs_field16_18 = _RAND_308[15:0];
  _RAND_309 = {1{`RANDOM}};
  fs_field16_19 = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  fs_field16_20 = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  fs_field16_21 = _RAND_311[15:0];
  _RAND_312 = {1{`RANDOM}};
  fs_field16_22 = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  fs_field16_23 = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  fs_field16_24 = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  fs_field16_25 = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  fs_field16_26 = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  fs_field16_27 = _RAND_317[15:0];
  _RAND_318 = {1{`RANDOM}};
  fs_field16_28 = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  fs_field16_29 = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  fs_field16_30 = _RAND_320[15:0];
  _RAND_321 = {1{`RANDOM}};
  fs_field16_31 = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  fs_field16_32 = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  fs_field16_33 = _RAND_323[15:0];
  _RAND_324 = {1{`RANDOM}};
  fs_field16_34 = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  fs_field16_35 = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  fs_field16_36 = _RAND_326[15:0];
  _RAND_327 = {1{`RANDOM}};
  fs_field16_37 = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  tag_0 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  tag_1 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  tag_2 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  tag_3 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  tag_4 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  tag_5 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  tag_6 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  tag_7 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  tag_8 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  tag_9 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  tag_10 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  tag_11 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  tag_12 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  tag_13 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  tag_14 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  tag_15 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  tag_16 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  tag_17 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  tag_18 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  tag_19 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  tag_20 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  tag_21 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  tag_22 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  tag_23 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  tag_24 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  tag_25 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  tag_26 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  tag_27 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  tag_28 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  tag_29 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  tag_30 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  tag_31 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  tag_32 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  tag_33 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  tag_34 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  tag_35 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  tag_36 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  tag_37 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  tag_38 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  tag_39 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  tag_40 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  tag_41 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  tag_42 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  tag_43 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  tag_44 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  tag_45 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  tag_46 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  tag_47 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  tag_48 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  tag_49 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  tag_50 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  tag_51 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  tag_52 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  tag_53 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  tag_54 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  tag_55 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  tag_56 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  tag_57 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  tag_58 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  tag_59 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  tag_60 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  tag_61 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  tag_62 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  tag_63 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  tag_64 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  tag_65 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  tag_66 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  tag_67 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  tag_68 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  tag_69 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  nid = _RAND_398[14:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
